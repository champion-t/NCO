module counter (clk,
    csb00,
    csb01,
    rst,
    addr00,
    addr01,
    denum,
    din00,
    din01,
    num,
    sine_out,
    vccd1,
    vssd1);
 input clk;
 input csb00;
 input csb01;
 input rst;
 input [7:0] addr00;
 input [7:0] addr01;
 input [3:0] denum;
 input [15:0] din00;
 input [15:0] din01;
 input [3:0] num;
 output [15:0] sine_out;
 inout vccd1;
 inout vssd1;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire \sine_out_reg0[0] ;
 wire \sine_out_reg0[10] ;
 wire \sine_out_reg0[11] ;
 wire \sine_out_reg0[12] ;
 wire \sine_out_reg0[13] ;
 wire \sine_out_reg0[14] ;
 wire \sine_out_reg0[15] ;
 wire \sine_out_reg0[1] ;
 wire \sine_out_reg0[2] ;
 wire \sine_out_reg0[3] ;
 wire \sine_out_reg0[4] ;
 wire \sine_out_reg0[5] ;
 wire \sine_out_reg0[6] ;
 wire \sine_out_reg0[7] ;
 wire \sine_out_reg0[8] ;
 wire \sine_out_reg0[9] ;
 wire \sine_out_reg1[0] ;
 wire \sine_out_reg1[10] ;
 wire \sine_out_reg1[11] ;
 wire \sine_out_reg1[12] ;
 wire \sine_out_reg1[13] ;
 wire \sine_out_reg1[14] ;
 wire \sine_out_reg1[15] ;
 wire \sine_out_reg1[1] ;
 wire \sine_out_reg1[2] ;
 wire \sine_out_reg1[3] ;
 wire \sine_out_reg1[4] ;
 wire \sine_out_reg1[5] ;
 wire \sine_out_reg1[6] ;
 wire \sine_out_reg1[7] ;
 wire \sine_out_reg1[8] ;
 wire \sine_out_reg1[9] ;
 wire \sine_out_temp0[0] ;
 wire \sine_out_temp0[10] ;
 wire \sine_out_temp0[11] ;
 wire \sine_out_temp0[12] ;
 wire \sine_out_temp0[13] ;
 wire \sine_out_temp0[14] ;
 wire \sine_out_temp0[15] ;
 wire \sine_out_temp0[1] ;
 wire \sine_out_temp0[2] ;
 wire \sine_out_temp0[3] ;
 wire \sine_out_temp0[4] ;
 wire \sine_out_temp0[5] ;
 wire \sine_out_temp0[6] ;
 wire \sine_out_temp0[7] ;
 wire \sine_out_temp0[8] ;
 wire \sine_out_temp0[9] ;
 wire \sine_out_temp1[0] ;
 wire \sine_out_temp1[10] ;
 wire \sine_out_temp1[11] ;
 wire \sine_out_temp1[12] ;
 wire \sine_out_temp1[13] ;
 wire \sine_out_temp1[14] ;
 wire \sine_out_temp1[15] ;
 wire \sine_out_temp1[1] ;
 wire \sine_out_temp1[2] ;
 wire \sine_out_temp1[3] ;
 wire \sine_out_temp1[4] ;
 wire \sine_out_temp1[5] ;
 wire \sine_out_temp1[6] ;
 wire \sine_out_temp1[7] ;
 wire \sine_out_temp1[8] ;
 wire \sine_out_temp1[9] ;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;
 wire \tcout[8] ;
 wire \tcout_delay[0] ;
 wire \tcout_delay[1] ;

 sky130_fd_sc_hd__inv_2 _297_ (.A(denum[3]),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _298_ (.A(denum[2]),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _299_ (.A(denum[0]),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _300_ (.A(num[0]),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _301_ (.A(num[3]),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _302_ (.A(num[1]),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _303_ (.A(num[2]),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _304_ (.A(rst),
    .Y(_025_));
 sky130_fd_sc_hd__or2_2 _305_ (.A(num[3]),
    .B(num[2]),
    .X(_057_));
 sky130_fd_sc_hd__or4b_2 _306_ (.A(num[3]),
    .B(num[1]),
    .C(num[2]),
    .D_N(num[0]),
    .X(_058_));
 sky130_fd_sc_hd__or3b_2 _307_ (.A(_050_),
    .B(num[1]),
    .C_N(_058_),
    .X(_059_));
 sky130_fd_sc_hd__nand2_2 _308_ (.A(_050_),
    .B(num[1]),
    .Y(_060_));
 sky130_fd_sc_hd__nand2_2 _309_ (.A(_051_),
    .B(num[0]),
    .Y(_061_));
 sky130_fd_sc_hd__and3_2 _310_ (.A(_059_),
    .B(_060_),
    .C(_061_),
    .X(_062_));
 sky130_fd_sc_hd__a221o_2 _311_ (.A1(_051_),
    .A2(num[0]),
    .B1(num[1]),
    .B2(_050_),
    .C1(_057_),
    .X(_063_));
 sky130_fd_sc_hd__a21boi_2 _312_ (.A1(denum[3]),
    .A2(_058_),
    .B1_N(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__a21oi_2 _313_ (.A1(_059_),
    .A2(_060_),
    .B1(_061_),
    .Y(_065_));
 sky130_fd_sc_hd__o21ba_2 _314_ (.A1(_062_),
    .A2(_065_),
    .B1_N(_063_),
    .X(_066_));
 sky130_fd_sc_hd__nand2_2 _315_ (.A(_050_),
    .B(num[3]),
    .Y(_067_));
 sky130_fd_sc_hd__a2111o_2 _316_ (.A1(_050_),
    .A2(num[1]),
    .B1(_057_),
    .C1(_051_),
    .D1(_053_),
    .X(_068_));
 sky130_fd_sc_hd__nand2_2 _317_ (.A(denum[2]),
    .B(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__and3_2 _318_ (.A(denum[2]),
    .B(_055_),
    .C(_068_),
    .X(_070_));
 sky130_fd_sc_hd__a21o_2 _319_ (.A1(denum[2]),
    .A2(_068_),
    .B1(_055_),
    .X(_071_));
 sky130_fd_sc_hd__and2b_2 _320_ (.A_N(_070_),
    .B(_071_),
    .X(_072_));
 sky130_fd_sc_hd__or2_2 _321_ (.A(denum[1]),
    .B(_053_),
    .X(_073_));
 sky130_fd_sc_hd__a21oi_2 _322_ (.A1(_071_),
    .A2(_073_),
    .B1(_070_),
    .Y(_074_));
 sky130_fd_sc_hd__nand2_2 _323_ (.A(num[2]),
    .B(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__or2_2 _324_ (.A(num[2]),
    .B(_074_),
    .X(_076_));
 sky130_fd_sc_hd__a311o_2 _325_ (.A1(_054_),
    .A2(_075_),
    .A3(_076_),
    .B1(_064_),
    .C1(_066_),
    .X(_077_));
 sky130_fd_sc_hd__nor2_2 _326_ (.A(num[3]),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__o31a_2 _327_ (.A1(num[2]),
    .A2(_064_),
    .A3(_066_),
    .B1(_074_),
    .X(_079_));
 sky130_fd_sc_hd__a21o_2 _328_ (.A1(_050_),
    .A2(num[2]),
    .B1(num[3]),
    .X(_080_));
 sky130_fd_sc_hd__nor2_2 _329_ (.A(_079_),
    .B(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__xnor2_2 _330_ (.A(_072_),
    .B(_073_),
    .Y(_082_));
 sky130_fd_sc_hd__mux2_1 _331_ (.A0(_069_),
    .A1(_082_),
    .S(_081_),
    .X(_083_));
 sky130_fd_sc_hd__nor2_2 _332_ (.A(num[2]),
    .B(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__xnor2_2 _333_ (.A(_056_),
    .B(_083_),
    .Y(_085_));
 sky130_fd_sc_hd__o31ai_2 _334_ (.A1(_053_),
    .A2(_079_),
    .A3(_080_),
    .B1(denum[1]),
    .Y(_086_));
 sky130_fd_sc_hd__or4_2 _335_ (.A(denum[1]),
    .B(_053_),
    .C(_079_),
    .D(_080_),
    .X(_087_));
 sky130_fd_sc_hd__and2_2 _336_ (.A(_086_),
    .B(_087_),
    .X(_088_));
 sky130_fd_sc_hd__a21o_2 _337_ (.A1(_086_),
    .A2(_087_),
    .B1(num[1]),
    .X(_089_));
 sky130_fd_sc_hd__nand3_2 _338_ (.A(num[1]),
    .B(_086_),
    .C(_087_),
    .Y(_090_));
 sky130_fd_sc_hd__nand2_2 _339_ (.A(_052_),
    .B(num[0]),
    .Y(_091_));
 sky130_fd_sc_hd__and3_2 _340_ (.A(_089_),
    .B(_090_),
    .C(_091_),
    .X(_092_));
 sky130_fd_sc_hd__a21bo_2 _341_ (.A1(_090_),
    .A2(_091_),
    .B1_N(_089_),
    .X(_093_));
 sky130_fd_sc_hd__a211o_2 _342_ (.A1(_085_),
    .A2(_093_),
    .B1(_078_),
    .C1(_084_),
    .X(_094_));
 sky130_fd_sc_hd__and2_2 _343_ (.A(_067_),
    .B(_094_),
    .X(_095_));
 sky130_fd_sc_hd__inv_2 _344_ (.A(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__xnor2_2 _345_ (.A(_085_),
    .B(_093_),
    .Y(_097_));
 sky130_fd_sc_hd__mux2_1 _346_ (.A0(_083_),
    .A1(_097_),
    .S(_095_),
    .X(_098_));
 sky130_fd_sc_hd__xnor2_2 _347_ (.A(num[3]),
    .B(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_2 _348_ (.A1(_089_),
    .A2(_090_),
    .B1(_091_),
    .Y(_100_));
 sky130_fd_sc_hd__or2_2 _349_ (.A(_092_),
    .B(_100_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _350_ (.A0(_088_),
    .A1(_101_),
    .S(_095_),
    .X(_102_));
 sky130_fd_sc_hd__or2_2 _351_ (.A(num[2]),
    .B(_102_),
    .X(_103_));
 sky130_fd_sc_hd__and2_2 _352_ (.A(num[2]),
    .B(_102_),
    .X(_104_));
 sky130_fd_sc_hd__a31o_2 _353_ (.A1(num[0]),
    .A2(_067_),
    .A3(_094_),
    .B1(_052_),
    .X(_105_));
 sky130_fd_sc_hd__nand3b_2 _354_ (.A_N(_091_),
    .B(_094_),
    .C(_067_),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_2 _355_ (.A(_105_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__a21oi_2 _356_ (.A1(_105_),
    .A2(_106_),
    .B1(num[1]),
    .Y(_108_));
 sky130_fd_sc_hd__and3_2 _357_ (.A(num[1]),
    .B(_105_),
    .C(_106_),
    .X(_109_));
 sky130_fd_sc_hd__or2_2 _358_ (.A(_108_),
    .B(_109_),
    .X(_110_));
 sky130_fd_sc_hd__o21ba_2 _359_ (.A1(num[0]),
    .A2(_109_),
    .B1_N(_108_),
    .X(_111_));
 sky130_fd_sc_hd__a21o_2 _360_ (.A1(_103_),
    .A2(_111_),
    .B1(_104_),
    .X(_112_));
 sky130_fd_sc_hd__a211o_2 _361_ (.A1(_103_),
    .A2(_111_),
    .B1(_104_),
    .C1(_099_),
    .X(_113_));
 sky130_fd_sc_hd__or3_2 _362_ (.A(_062_),
    .B(_063_),
    .C(_065_),
    .X(_114_));
 sky130_fd_sc_hd__o221a_2 _363_ (.A1(_077_),
    .A2(_095_),
    .B1(_098_),
    .B2(num[3]),
    .C1(_114_),
    .X(_115_));
 sky130_fd_sc_hd__and2_2 _364_ (.A(_113_),
    .B(_115_),
    .X(_116_));
 sky130_fd_sc_hd__nand2_2 _365_ (.A(_113_),
    .B(_115_),
    .Y(_117_));
 sky130_fd_sc_hd__a21bo_2 _366_ (.A1(_098_),
    .A2(_115_),
    .B1_N(_113_),
    .X(_118_));
 sky130_fd_sc_hd__a21oi_2 _367_ (.A1(_099_),
    .A2(_112_),
    .B1(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__xnor2_2 _368_ (.A(_056_),
    .B(_102_),
    .Y(_120_));
 sky130_fd_sc_hd__nand2_2 _369_ (.A(_111_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__or2_2 _370_ (.A(_111_),
    .B(_120_),
    .X(_122_));
 sky130_fd_sc_hd__nand3b_2 _371_ (.A_N(_102_),
    .B(_113_),
    .C(_115_),
    .Y(_123_));
 sky130_fd_sc_hd__a22o_2 _372_ (.A1(_113_),
    .A2(_115_),
    .B1(_121_),
    .B2(_122_),
    .X(_124_));
 sky130_fd_sc_hd__and2_2 _373_ (.A(_123_),
    .B(_124_),
    .X(_125_));
 sky130_fd_sc_hd__a21oi_2 _374_ (.A1(_123_),
    .A2(_124_),
    .B1(num[3]),
    .Y(_126_));
 sky130_fd_sc_hd__nand2_2 _375_ (.A(num[3]),
    .B(_125_),
    .Y(_127_));
 sky130_fd_sc_hd__and3_2 _376_ (.A(_107_),
    .B(_113_),
    .C(_115_),
    .X(_128_));
 sky130_fd_sc_hd__xnor2_2 _377_ (.A(_053_),
    .B(_110_),
    .Y(_129_));
 sky130_fd_sc_hd__a21o_2 _378_ (.A1(_113_),
    .A2(_115_),
    .B1(_129_),
    .X(_130_));
 sky130_fd_sc_hd__o21a_2 _379_ (.A1(_107_),
    .A2(_117_),
    .B1(_130_),
    .X(_131_));
 sky130_fd_sc_hd__inv_2 _380_ (.A(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__o211a_2 _381_ (.A1(_107_),
    .A2(_117_),
    .B1(_130_),
    .C1(_056_),
    .X(_133_));
 sky130_fd_sc_hd__a211o_2 _382_ (.A1(_117_),
    .A2(_129_),
    .B1(_128_),
    .C1(_056_),
    .X(_134_));
 sky130_fd_sc_hd__and2b_2 _383_ (.A_N(_133_),
    .B(_134_),
    .X(_135_));
 sky130_fd_sc_hd__a21oi_2 _384_ (.A1(num[0]),
    .A2(_116_),
    .B1(num[1]),
    .Y(_136_));
 sky130_fd_sc_hd__a21oi_2 _385_ (.A1(_134_),
    .A2(_136_),
    .B1(_133_),
    .Y(_137_));
 sky130_fd_sc_hd__a211o_2 _386_ (.A1(_134_),
    .A2(_136_),
    .B1(_126_),
    .C1(_133_),
    .X(_138_));
 sky130_fd_sc_hd__a21oi_2 _387_ (.A1(_127_),
    .A2(_138_),
    .B1(_119_),
    .Y(_139_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__xnor2_2 _389_ (.A(_135_),
    .B(_136_),
    .Y(_141_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(_141_),
    .A1(_132_),
    .S(_139_),
    .X(_142_));
 sky130_fd_sc_hd__nand2_2 _391_ (.A(num[3]),
    .B(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__a211oi_2 _392_ (.A1(_127_),
    .A2(_138_),
    .B1(_053_),
    .C1(_119_),
    .Y(_144_));
 sky130_fd_sc_hd__and3_2 _393_ (.A(num[0]),
    .B(num[1]),
    .C(_116_),
    .X(_145_));
 sky130_fd_sc_hd__or2_2 _394_ (.A(_136_),
    .B(_145_),
    .X(_146_));
 sky130_fd_sc_hd__o2bb2a_2 _395_ (.A1_N(_117_),
    .A2_N(_144_),
    .B1(_146_),
    .B2(_139_),
    .X(_147_));
 sky130_fd_sc_hd__nand2_2 _396_ (.A(num[2]),
    .B(_147_),
    .Y(_148_));
 sky130_fd_sc_hd__nor2_2 _397_ (.A(num[1]),
    .B(_144_),
    .Y(_149_));
 sky130_fd_sc_hd__o21bai_2 _398_ (.A1(num[2]),
    .A2(_147_),
    .B1_N(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__and2_2 _399_ (.A(_148_),
    .B(_150_),
    .X(_151_));
 sky130_fd_sc_hd__nand2_2 _400_ (.A(_143_),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__or2_2 _401_ (.A(num[3]),
    .B(_142_),
    .X(_153_));
 sky130_fd_sc_hd__xnor2_2 _402_ (.A(_054_),
    .B(_137_),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_2 _403_ (.A(_119_),
    .B(_125_),
    .Y(_155_));
 sky130_fd_sc_hd__mux2_1 _404_ (.A0(_125_),
    .A1(_155_),
    .S(_154_),
    .X(_156_));
 sky130_fd_sc_hd__o21ai_2 _405_ (.A1(num[3]),
    .A2(_142_),
    .B1(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__a31oi_2 _406_ (.A1(_143_),
    .A2(_148_),
    .A3(_150_),
    .B1(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__nand2_2 _407_ (.A(_143_),
    .B(_153_),
    .Y(_159_));
 sky130_fd_sc_hd__xor2_2 _408_ (.A(_151_),
    .B(_159_),
    .X(_160_));
 sky130_fd_sc_hd__mux2_1 _409_ (.A0(_160_),
    .A1(_142_),
    .S(_158_),
    .X(_161_));
 sky130_fd_sc_hd__a21o_2 _410_ (.A1(_152_),
    .A2(_153_),
    .B1(_156_),
    .X(_162_));
 sky130_fd_sc_hd__nand3_2 _411_ (.A(_119_),
    .B(_127_),
    .C(_138_),
    .Y(_163_));
 sky130_fd_sc_hd__nand4_2 _412_ (.A(_114_),
    .B(_161_),
    .C(_162_),
    .D(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__xnor2_2 _413_ (.A(_056_),
    .B(_147_),
    .Y(_165_));
 sky130_fd_sc_hd__xnor2_2 _414_ (.A(_149_),
    .B(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__mux2_1 _415_ (.A0(_166_),
    .A1(_147_),
    .S(_158_),
    .X(_167_));
 sky130_fd_sc_hd__nor2_2 _416_ (.A(num[3]),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__nand2_2 _417_ (.A(num[3]),
    .B(_167_),
    .Y(_169_));
 sky130_fd_sc_hd__a311oi_2 _418_ (.A1(_143_),
    .A2(_148_),
    .A3(_150_),
    .B1(_157_),
    .C1(_053_),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_2 _419_ (.A(num[1]),
    .B(_144_),
    .Y(_171_));
 sky130_fd_sc_hd__nand2b_2 _420_ (.A_N(_149_),
    .B(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__o2bb2a_2 _421_ (.A1_N(_140_),
    .A2_N(_170_),
    .B1(_172_),
    .B2(_158_),
    .X(_173_));
 sky130_fd_sc_hd__nor2_2 _422_ (.A(num[2]),
    .B(_173_),
    .Y(_174_));
 sky130_fd_sc_hd__xnor2_2 _423_ (.A(_056_),
    .B(_173_),
    .Y(_175_));
 sky130_fd_sc_hd__nor2_2 _424_ (.A(num[1]),
    .B(_170_),
    .Y(_176_));
 sky130_fd_sc_hd__a21o_2 _425_ (.A1(_175_),
    .A2(_176_),
    .B1(_174_),
    .X(_177_));
 sky130_fd_sc_hd__a211o_2 _426_ (.A1(_175_),
    .A2(_176_),
    .B1(_168_),
    .C1(_174_),
    .X(_178_));
 sky130_fd_sc_hd__a21o_2 _427_ (.A1(_169_),
    .A2(_178_),
    .B1(_164_),
    .X(_179_));
 sky130_fd_sc_hd__xnor2_2 _428_ (.A(_175_),
    .B(_176_),
    .Y(_180_));
 sky130_fd_sc_hd__mux2_1 _429_ (.A0(_173_),
    .A1(_180_),
    .S(_179_),
    .X(_181_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__or2_2 _431_ (.A(num[3]),
    .B(_181_),
    .X(_183_));
 sky130_fd_sc_hd__xnor2_2 _432_ (.A(num[3]),
    .B(_181_),
    .Y(_184_));
 sky130_fd_sc_hd__a211o_2 _433_ (.A1(_169_),
    .A2(_178_),
    .B1(_053_),
    .C1(_164_),
    .X(_185_));
 sky130_fd_sc_hd__and2_2 _434_ (.A(num[1]),
    .B(_170_),
    .X(_186_));
 sky130_fd_sc_hd__nor2_2 _435_ (.A(_176_),
    .B(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__o2bb2a_2 _436_ (.A1_N(_187_),
    .A2_N(_179_),
    .B1(_158_),
    .B2(_185_),
    .X(_188_));
 sky130_fd_sc_hd__and2_2 _437_ (.A(num[2]),
    .B(_188_),
    .X(_189_));
 sky130_fd_sc_hd__and2_2 _438_ (.A(_055_),
    .B(_185_),
    .X(_190_));
 sky130_fd_sc_hd__o21ba_2 _439_ (.A1(num[2]),
    .A2(_188_),
    .B1_N(_190_),
    .X(_191_));
 sky130_fd_sc_hd__or2_2 _440_ (.A(_189_),
    .B(_191_),
    .X(_192_));
 sky130_fd_sc_hd__nand2b_2 _441_ (.A_N(_168_),
    .B(_169_),
    .Y(_193_));
 sky130_fd_sc_hd__xor2_2 _442_ (.A(_177_),
    .B(_193_),
    .X(_194_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(_167_),
    .A1(_194_),
    .S(_179_),
    .X(_195_));
 sky130_fd_sc_hd__o311a_2 _444_ (.A1(_184_),
    .A2(_189_),
    .A3(_191_),
    .B1(_195_),
    .C1(_183_),
    .X(_196_));
 sky130_fd_sc_hd__xnor2_2 _445_ (.A(_056_),
    .B(_188_),
    .Y(_197_));
 sky130_fd_sc_hd__xnor2_2 _446_ (.A(_190_),
    .B(_197_),
    .Y(_198_));
 sky130_fd_sc_hd__mux2_1 _447_ (.A0(_198_),
    .A1(_188_),
    .S(_196_),
    .X(_199_));
 sky130_fd_sc_hd__and2_2 _448_ (.A(num[3]),
    .B(_199_),
    .X(_200_));
 sky130_fd_sc_hd__nand2_2 _449_ (.A(num[3]),
    .B(_199_),
    .Y(_201_));
 sky130_fd_sc_hd__nand2_2 _450_ (.A(num[0]),
    .B(_179_),
    .Y(_202_));
 sky130_fd_sc_hd__nor2_2 _451_ (.A(_055_),
    .B(_185_),
    .Y(_203_));
 sky130_fd_sc_hd__or2_2 _452_ (.A(_190_),
    .B(_203_),
    .X(_204_));
 sky130_fd_sc_hd__mux2_1 _453_ (.A0(_204_),
    .A1(_202_),
    .S(_196_),
    .X(_205_));
 sky130_fd_sc_hd__nor2_2 _454_ (.A(num[2]),
    .B(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__xnor2_2 _455_ (.A(_056_),
    .B(_205_),
    .Y(_207_));
 sky130_fd_sc_hd__a21oi_2 _456_ (.A1(num[0]),
    .A2(_196_),
    .B1(num[1]),
    .Y(_208_));
 sky130_fd_sc_hd__a21o_2 _457_ (.A1(_207_),
    .A2(_208_),
    .B1(_206_),
    .X(_209_));
 sky130_fd_sc_hd__nor2_2 _458_ (.A(num[3]),
    .B(_199_),
    .Y(_210_));
 sky130_fd_sc_hd__nor2_2 _459_ (.A(_200_),
    .B(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__a21oi_2 _460_ (.A1(_184_),
    .A2(_192_),
    .B1(_196_),
    .Y(_212_));
 sky130_fd_sc_hd__o21a_2 _461_ (.A1(_184_),
    .A2(_192_),
    .B1(_212_),
    .X(_213_));
 sky130_fd_sc_hd__and3_2 _462_ (.A(_164_),
    .B(_169_),
    .C(_178_),
    .X(_214_));
 sky130_fd_sc_hd__a2111o_2 _463_ (.A1(_182_),
    .A2(_196_),
    .B1(_210_),
    .C1(_213_),
    .D1(_214_),
    .X(_215_));
 sky130_fd_sc_hd__a21oi_2 _464_ (.A1(_201_),
    .A2(_209_),
    .B1(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__xnor2_2 _465_ (.A(_207_),
    .B(_208_),
    .Y(_217_));
 sky130_fd_sc_hd__mux2_1 _466_ (.A0(_217_),
    .A1(_205_),
    .S(_216_),
    .X(_218_));
 sky130_fd_sc_hd__nand2_2 _467_ (.A(num[3]),
    .B(_218_),
    .Y(_219_));
 sky130_fd_sc_hd__a211o_2 _468_ (.A1(_201_),
    .A2(_209_),
    .B1(_215_),
    .C1(_053_),
    .X(_220_));
 sky130_fd_sc_hd__and3_2 _469_ (.A(num[0]),
    .B(num[1]),
    .C(_196_),
    .X(_221_));
 sky130_fd_sc_hd__o32a_2 _470_ (.A1(_208_),
    .A2(_216_),
    .A3(_221_),
    .B1(_220_),
    .B2(_196_),
    .X(_222_));
 sky130_fd_sc_hd__nand2_2 _471_ (.A(num[2]),
    .B(_222_),
    .Y(_223_));
 sky130_fd_sc_hd__and2_2 _472_ (.A(_055_),
    .B(_220_),
    .X(_224_));
 sky130_fd_sc_hd__o21bai_2 _473_ (.A1(num[2]),
    .A2(_222_),
    .B1_N(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__xnor2_2 _474_ (.A(_209_),
    .B(_211_),
    .Y(_226_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(_226_),
    .A1(_199_),
    .S(_216_),
    .X(_227_));
 sky130_fd_sc_hd__inv_2 _476_ (.A(_227_),
    .Y(_228_));
 sky130_fd_sc_hd__o21ai_2 _477_ (.A1(num[3]),
    .A2(_218_),
    .B1(_227_),
    .Y(_229_));
 sky130_fd_sc_hd__a31oi_2 _478_ (.A1(_219_),
    .A2(_223_),
    .A3(_225_),
    .B1(_229_),
    .Y(_230_));
 sky130_fd_sc_hd__a311o_2 _479_ (.A1(_219_),
    .A2(_223_),
    .A3(_225_),
    .B1(_229_),
    .C1(_053_),
    .X(_231_));
 sky130_fd_sc_hd__or3b_2 _480_ (.A(num[1]),
    .B(num[2]),
    .C_N(_231_),
    .X(_232_));
 sky130_fd_sc_hd__nor2_2 _481_ (.A(_055_),
    .B(_220_),
    .Y(_233_));
 sky130_fd_sc_hd__o32a_2 _482_ (.A1(_224_),
    .A2(_230_),
    .A3(_233_),
    .B1(_231_),
    .B2(_216_),
    .X(_234_));
 sky130_fd_sc_hd__xnor2_2 _483_ (.A(_056_),
    .B(_222_),
    .Y(_235_));
 sky130_fd_sc_hd__xnor2_2 _484_ (.A(_224_),
    .B(_235_),
    .Y(_236_));
 sky130_fd_sc_hd__mux2_1 _485_ (.A0(_236_),
    .A1(_222_),
    .S(_230_),
    .X(_237_));
 sky130_fd_sc_hd__a21oi_2 _486_ (.A1(_055_),
    .A2(_231_),
    .B1(_056_),
    .Y(_238_));
 sky130_fd_sc_hd__a221o_2 _487_ (.A1(_232_),
    .A2(_234_),
    .B1(_237_),
    .B2(num[3]),
    .C1(_238_),
    .X(_239_));
 sky130_fd_sc_hd__a21bo_2 _488_ (.A1(_218_),
    .A2(_227_),
    .B1_N(_230_),
    .X(_240_));
 sky130_fd_sc_hd__a22o_2 _489_ (.A1(_223_),
    .A2(_225_),
    .B1(_228_),
    .B2(_219_),
    .X(_241_));
 sky130_fd_sc_hd__a21oi_2 _490_ (.A1(_229_),
    .A2(_241_),
    .B1(_214_),
    .Y(_242_));
 sky130_fd_sc_hd__o211a_2 _491_ (.A1(num[3]),
    .A2(_237_),
    .B1(_240_),
    .C1(_242_),
    .X(_243_));
 sky130_fd_sc_hd__and2_2 _492_ (.A(_239_),
    .B(_243_),
    .X(_244_));
 sky130_fd_sc_hd__and4_2 _493_ (.A(_216_),
    .B(_230_),
    .C(_239_),
    .D(_243_),
    .X(_245_));
 sky130_fd_sc_hd__nand2_2 _494_ (.A(_196_),
    .B(_245_),
    .Y(_246_));
 sky130_fd_sc_hd__and4_2 _495_ (.A(_139_),
    .B(_158_),
    .C(_196_),
    .D(_245_),
    .X(_247_));
 sky130_fd_sc_hd__nand4_2 _496_ (.A(_139_),
    .B(_158_),
    .C(_196_),
    .D(_245_),
    .Y(_248_));
 sky130_fd_sc_hd__xnor2_2 _497_ (.A(_117_),
    .B(_247_),
    .Y(_249_));
 sky130_fd_sc_hd__xnor2_2 _498_ (.A(\tcout[7] ),
    .B(_249_),
    .Y(_250_));
 sky130_fd_sc_hd__a31o_2 _499_ (.A1(_158_),
    .A2(_196_),
    .A3(_245_),
    .B1(_139_),
    .X(_251_));
 sky130_fd_sc_hd__and3_2 _500_ (.A(\tcout[6] ),
    .B(_248_),
    .C(_251_),
    .X(_252_));
 sky130_fd_sc_hd__xnor2_2 _501_ (.A(_158_),
    .B(_246_),
    .Y(_253_));
 sky130_fd_sc_hd__xnor2_2 _502_ (.A(\tcout[5] ),
    .B(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__a21oi_2 _503_ (.A1(_248_),
    .A2(_251_),
    .B1(\tcout[6] ),
    .Y(_255_));
 sky130_fd_sc_hd__xor2_2 _504_ (.A(_196_),
    .B(_245_),
    .X(_256_));
 sky130_fd_sc_hd__xnor2_2 _505_ (.A(\tcout[3] ),
    .B(_256_),
    .Y(_257_));
 sky130_fd_sc_hd__a21oi_2 _506_ (.A1(_196_),
    .A2(_245_),
    .B1(_179_),
    .Y(_258_));
 sky130_fd_sc_hd__xnor2_2 _507_ (.A(\tcout[4] ),
    .B(_258_),
    .Y(_259_));
 sky130_fd_sc_hd__a31o_2 _508_ (.A1(_230_),
    .A2(_239_),
    .A3(_243_),
    .B1(_216_),
    .X(_260_));
 sky130_fd_sc_hd__and2b_2 _509_ (.A_N(_245_),
    .B(_260_),
    .X(_261_));
 sky130_fd_sc_hd__xnor2_2 _510_ (.A(\tcout[1] ),
    .B(_230_),
    .Y(_262_));
 sky130_fd_sc_hd__nand2_2 _511_ (.A(\tcout[0] ),
    .B(_262_),
    .Y(_263_));
 sky130_fd_sc_hd__o21ba_2 _512_ (.A1(\tcout[0] ),
    .A2(_262_),
    .B1_N(_244_),
    .X(_264_));
 sky130_fd_sc_hd__a221o_2 _513_ (.A1(\tcout[8] ),
    .A2(_096_),
    .B1(_244_),
    .B2(_263_),
    .C1(_264_),
    .X(_265_));
 sky130_fd_sc_hd__xnor2_2 _514_ (.A(\tcout[2] ),
    .B(_261_),
    .Y(_266_));
 sky130_fd_sc_hd__or4_2 _515_ (.A(_257_),
    .B(_259_),
    .C(_265_),
    .D(_266_),
    .X(_267_));
 sky130_fd_sc_hd__or2_2 _516_ (.A(\tcout[8] ),
    .B(_096_),
    .X(_268_));
 sky130_fd_sc_hd__and3_2 _517_ (.A(_116_),
    .B(_247_),
    .C(_268_),
    .X(_269_));
 sky130_fd_sc_hd__a21oi_2 _518_ (.A1(_116_),
    .A2(_247_),
    .B1(_268_),
    .Y(_270_));
 sky130_fd_sc_hd__or4_2 _519_ (.A(_252_),
    .B(_255_),
    .C(_269_),
    .D(_270_),
    .X(_271_));
 sky130_fd_sc_hd__or4_2 _520_ (.A(_250_),
    .B(_254_),
    .C(_267_),
    .D(_271_),
    .X(_272_));
 sky130_fd_sc_hd__and2b_2 _521_ (.A_N(\tcout[0] ),
    .B(_272_),
    .X(_016_));
 sky130_fd_sc_hd__or2_2 _522_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .X(_273_));
 sky130_fd_sc_hd__nand2_2 _523_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .Y(_274_));
 sky130_fd_sc_hd__and3_2 _524_ (.A(_272_),
    .B(_273_),
    .C(_274_),
    .X(_017_));
 sky130_fd_sc_hd__nand3_2 _525_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .Y(_275_));
 sky130_fd_sc_hd__a21o_2 _526_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1(\tcout[2] ),
    .X(_276_));
 sky130_fd_sc_hd__and3_2 _527_ (.A(_272_),
    .B(_275_),
    .C(_276_),
    .X(_018_));
 sky130_fd_sc_hd__and4_2 _528_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .D(\tcout[3] ),
    .X(_277_));
 sky130_fd_sc_hd__inv_2 _529_ (.A(_277_),
    .Y(_278_));
 sky130_fd_sc_hd__a31o_2 _530_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .A3(\tcout[2] ),
    .B1(\tcout[3] ),
    .X(_279_));
 sky130_fd_sc_hd__and3_2 _531_ (.A(_272_),
    .B(_278_),
    .C(_279_),
    .X(_019_));
 sky130_fd_sc_hd__nand2_2 _532_ (.A(\tcout[4] ),
    .B(_277_),
    .Y(_280_));
 sky130_fd_sc_hd__or2_2 _533_ (.A(\tcout[4] ),
    .B(_277_),
    .X(_281_));
 sky130_fd_sc_hd__and3_2 _534_ (.A(_272_),
    .B(_280_),
    .C(_281_),
    .X(_020_));
 sky130_fd_sc_hd__and3_2 _535_ (.A(\tcout[4] ),
    .B(\tcout[5] ),
    .C(_277_),
    .X(_282_));
 sky130_fd_sc_hd__inv_2 _536_ (.A(_282_),
    .Y(_283_));
 sky130_fd_sc_hd__a21o_2 _537_ (.A1(\tcout[4] ),
    .A2(_277_),
    .B1(\tcout[5] ),
    .X(_284_));
 sky130_fd_sc_hd__and3_2 _538_ (.A(_272_),
    .B(_283_),
    .C(_284_),
    .X(_021_));
 sky130_fd_sc_hd__and2_2 _539_ (.A(\tcout[6] ),
    .B(_282_),
    .X(_285_));
 sky130_fd_sc_hd__nand2_2 _540_ (.A(\tcout[6] ),
    .B(_282_),
    .Y(_286_));
 sky130_fd_sc_hd__or2_2 _541_ (.A(\tcout[6] ),
    .B(_282_),
    .X(_287_));
 sky130_fd_sc_hd__and3_2 _542_ (.A(_272_),
    .B(_286_),
    .C(_287_),
    .X(_022_));
 sky130_fd_sc_hd__nand2_2 _543_ (.A(\tcout[7] ),
    .B(_285_),
    .Y(_288_));
 sky130_fd_sc_hd__or2_2 _544_ (.A(\tcout[7] ),
    .B(_285_),
    .X(_289_));
 sky130_fd_sc_hd__and3_2 _545_ (.A(_272_),
    .B(_288_),
    .C(_289_),
    .X(_023_));
 sky130_fd_sc_hd__xnor2_2 _546_ (.A(\tcout[8] ),
    .B(_288_),
    .Y(_290_));
 sky130_fd_sc_hd__and2_2 _547_ (.A(_272_),
    .B(_290_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _548_ (.A0(\sine_out_reg0[0] ),
    .A1(\sine_out_reg1[0] ),
    .S(\tcout_delay[0] ),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _549_ (.A0(\sine_out_reg0[1] ),
    .A1(\sine_out_reg1[1] ),
    .S(\tcout_delay[0] ),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _550_ (.A0(\sine_out_reg0[2] ),
    .A1(\sine_out_reg1[2] ),
    .S(\tcout_delay[0] ),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _551_ (.A0(\sine_out_reg0[3] ),
    .A1(\sine_out_reg1[3] ),
    .S(\tcout_delay[0] ),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _552_ (.A0(\sine_out_reg0[4] ),
    .A1(\sine_out_reg1[4] ),
    .S(\tcout_delay[0] ),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _553_ (.A0(\sine_out_reg0[5] ),
    .A1(\sine_out_reg1[5] ),
    .S(\tcout_delay[0] ),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _554_ (.A0(\sine_out_reg0[6] ),
    .A1(\sine_out_reg1[6] ),
    .S(\tcout_delay[0] ),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _555_ (.A0(\sine_out_reg0[7] ),
    .A1(\sine_out_reg1[7] ),
    .S(\tcout_delay[0] ),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _556_ (.A0(\sine_out_reg0[8] ),
    .A1(\sine_out_reg1[8] ),
    .S(\tcout_delay[0] ),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _557_ (.A0(\sine_out_reg0[9] ),
    .A1(\sine_out_reg1[9] ),
    .S(\tcout_delay[0] ),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _558_ (.A0(\sine_out_reg0[10] ),
    .A1(\sine_out_reg1[10] ),
    .S(\tcout_delay[0] ),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _559_ (.A0(\sine_out_reg0[11] ),
    .A1(\sine_out_reg1[11] ),
    .S(\tcout_delay[0] ),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _560_ (.A0(\sine_out_reg0[12] ),
    .A1(\sine_out_reg1[12] ),
    .S(\tcout_delay[0] ),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _561_ (.A0(\sine_out_reg0[13] ),
    .A1(\sine_out_reg1[13] ),
    .S(\tcout_delay[0] ),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _562_ (.A0(\sine_out_reg0[14] ),
    .A1(\sine_out_reg1[14] ),
    .S(\tcout_delay[0] ),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _563_ (.A0(\sine_out_reg0[15] ),
    .A1(\sine_out_reg1[15] ),
    .S(\tcout_delay[0] ),
    .X(_006_));
 sky130_fd_sc_hd__inv_2 _564_ (.A(rst),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _565_ (.A(rst),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _566_ (.A(rst),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _567_ (.A(rst),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _568_ (.A(rst),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _569_ (.A(rst),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _570_ (.A(rst),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _571_ (.A(rst),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _572_ (.A(rst),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _573_ (.A(rst),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _574_ (.A(rst),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _575_ (.A(rst),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _576_ (.A(rst),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _577_ (.A(rst),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _578_ (.A(rst),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _579_ (.A(rst),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _580_ (.A(rst),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _581_ (.A(rst),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _582_ (.A(rst),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _583_ (.A(rst),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _584_ (.A(rst),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _585_ (.A(rst),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _586_ (.A(rst),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _587_ (.A(rst),
    .Y(_049_));
 sky130_fd_sc_hd__dfrtp_2 _588_ (.CLK(clk),
    .D(_000_),
    .RESET_B(_025_),
    .Q(sine_out[0]));
 sky130_fd_sc_hd__dfrtp_2 _589_ (.CLK(clk),
    .D(_007_),
    .RESET_B(_026_),
    .Q(sine_out[1]));
 sky130_fd_sc_hd__dfrtp_2 _590_ (.CLK(clk),
    .D(_008_),
    .RESET_B(_027_),
    .Q(sine_out[2]));
 sky130_fd_sc_hd__dfrtp_2 _591_ (.CLK(clk),
    .D(_009_),
    .RESET_B(_028_),
    .Q(sine_out[3]));
 sky130_fd_sc_hd__dfrtp_2 _592_ (.CLK(clk),
    .D(_010_),
    .RESET_B(_029_),
    .Q(sine_out[4]));
 sky130_fd_sc_hd__dfrtp_2 _593_ (.CLK(clk),
    .D(_011_),
    .RESET_B(_030_),
    .Q(sine_out[5]));
 sky130_fd_sc_hd__dfrtp_2 _594_ (.CLK(clk),
    .D(_012_),
    .RESET_B(_031_),
    .Q(sine_out[6]));
 sky130_fd_sc_hd__dfrtp_2 _595_ (.CLK(clk),
    .D(_013_),
    .RESET_B(_032_),
    .Q(sine_out[7]));
 sky130_fd_sc_hd__dfrtp_2 _596_ (.CLK(clk),
    .D(_014_),
    .RESET_B(_033_),
    .Q(sine_out[8]));
 sky130_fd_sc_hd__dfrtp_2 _597_ (.CLK(clk),
    .D(_015_),
    .RESET_B(_034_),
    .Q(sine_out[9]));
 sky130_fd_sc_hd__dfrtp_2 _598_ (.CLK(clk),
    .D(_001_),
    .RESET_B(_035_),
    .Q(sine_out[10]));
 sky130_fd_sc_hd__dfrtp_2 _599_ (.CLK(clk),
    .D(_002_),
    .RESET_B(_036_),
    .Q(sine_out[11]));
 sky130_fd_sc_hd__dfrtp_2 _600_ (.CLK(clk),
    .D(_003_),
    .RESET_B(_037_),
    .Q(sine_out[12]));
 sky130_fd_sc_hd__dfrtp_2 _601_ (.CLK(clk),
    .D(_004_),
    .RESET_B(_038_),
    .Q(sine_out[13]));
 sky130_fd_sc_hd__dfrtp_2 _602_ (.CLK(clk),
    .D(_005_),
    .RESET_B(_039_),
    .Q(sine_out[14]));
 sky130_fd_sc_hd__dfrtp_2 _603_ (.CLK(clk),
    .D(_006_),
    .RESET_B(_040_),
    .Q(sine_out[15]));
 sky130_fd_sc_hd__dfrtp_2 _604_ (.CLK(clk),
    .D(_016_),
    .RESET_B(_041_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_2 _605_ (.CLK(clk),
    .D(_017_),
    .RESET_B(_042_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_2 _606_ (.CLK(clk),
    .D(_018_),
    .RESET_B(_043_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_2 _607_ (.CLK(clk),
    .D(_019_),
    .RESET_B(_044_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_2 _608_ (.CLK(clk),
    .D(_020_),
    .RESET_B(_045_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_2 _609_ (.CLK(clk),
    .D(_021_),
    .RESET_B(_046_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_2 _610_ (.CLK(clk),
    .D(_022_),
    .RESET_B(_047_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_2 _611_ (.CLK(clk),
    .D(_023_),
    .RESET_B(_048_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__dfrtp_2 _612_ (.CLK(clk),
    .D(_024_),
    .RESET_B(_049_),
    .Q(\tcout[8] ));
 sky130_fd_sc_hd__dfxtp_2 _613_ (.CLK(clk),
    .D(\sine_out_temp0[0] ),
    .Q(\sine_out_reg0[0] ));
 sky130_fd_sc_hd__dfxtp_2 _614_ (.CLK(clk),
    .D(\sine_out_temp0[1] ),
    .Q(\sine_out_reg0[1] ));
 sky130_fd_sc_hd__dfxtp_2 _615_ (.CLK(clk),
    .D(\sine_out_temp0[2] ),
    .Q(\sine_out_reg0[2] ));
 sky130_fd_sc_hd__dfxtp_2 _616_ (.CLK(clk),
    .D(\sine_out_temp0[3] ),
    .Q(\sine_out_reg0[3] ));
 sky130_fd_sc_hd__dfxtp_2 _617_ (.CLK(clk),
    .D(\sine_out_temp0[4] ),
    .Q(\sine_out_reg0[4] ));
 sky130_fd_sc_hd__dfxtp_2 _618_ (.CLK(clk),
    .D(\sine_out_temp0[5] ),
    .Q(\sine_out_reg0[5] ));
 sky130_fd_sc_hd__dfxtp_2 _619_ (.CLK(clk),
    .D(\sine_out_temp0[6] ),
    .Q(\sine_out_reg0[6] ));
 sky130_fd_sc_hd__dfxtp_2 _620_ (.CLK(clk),
    .D(\sine_out_temp0[7] ),
    .Q(\sine_out_reg0[7] ));
 sky130_fd_sc_hd__dfxtp_2 _621_ (.CLK(clk),
    .D(\sine_out_temp0[8] ),
    .Q(\sine_out_reg0[8] ));
 sky130_fd_sc_hd__dfxtp_2 _622_ (.CLK(clk),
    .D(\sine_out_temp0[9] ),
    .Q(\sine_out_reg0[9] ));
 sky130_fd_sc_hd__dfxtp_2 _623_ (.CLK(clk),
    .D(\sine_out_temp0[10] ),
    .Q(\sine_out_reg0[10] ));
 sky130_fd_sc_hd__dfxtp_2 _624_ (.CLK(clk),
    .D(\sine_out_temp0[11] ),
    .Q(\sine_out_reg0[11] ));
 sky130_fd_sc_hd__dfxtp_2 _625_ (.CLK(clk),
    .D(\sine_out_temp0[12] ),
    .Q(\sine_out_reg0[12] ));
 sky130_fd_sc_hd__dfxtp_2 _626_ (.CLK(clk),
    .D(\sine_out_temp0[13] ),
    .Q(\sine_out_reg0[13] ));
 sky130_fd_sc_hd__dfxtp_2 _627_ (.CLK(clk),
    .D(\sine_out_temp0[14] ),
    .Q(\sine_out_reg0[14] ));
 sky130_fd_sc_hd__dfxtp_2 _628_ (.CLK(clk),
    .D(\sine_out_temp0[15] ),
    .Q(\sine_out_reg0[15] ));
 sky130_fd_sc_hd__dfxtp_2 _629_ (.CLK(clk),
    .D(\sine_out_temp1[0] ),
    .Q(\sine_out_reg1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _630_ (.CLK(clk),
    .D(\sine_out_temp1[1] ),
    .Q(\sine_out_reg1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _631_ (.CLK(clk),
    .D(\sine_out_temp1[2] ),
    .Q(\sine_out_reg1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _632_ (.CLK(clk),
    .D(\sine_out_temp1[3] ),
    .Q(\sine_out_reg1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _633_ (.CLK(clk),
    .D(\sine_out_temp1[4] ),
    .Q(\sine_out_reg1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _634_ (.CLK(clk),
    .D(\sine_out_temp1[5] ),
    .Q(\sine_out_reg1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _635_ (.CLK(clk),
    .D(\sine_out_temp1[6] ),
    .Q(\sine_out_reg1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _636_ (.CLK(clk),
    .D(\sine_out_temp1[7] ),
    .Q(\sine_out_reg1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _637_ (.CLK(clk),
    .D(\sine_out_temp1[8] ),
    .Q(\sine_out_reg1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _638_ (.CLK(clk),
    .D(\sine_out_temp1[9] ),
    .Q(\sine_out_reg1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _639_ (.CLK(clk),
    .D(\sine_out_temp1[10] ),
    .Q(\sine_out_reg1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _640_ (.CLK(clk),
    .D(\sine_out_temp1[11] ),
    .Q(\sine_out_reg1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _641_ (.CLK(clk),
    .D(\sine_out_temp1[12] ),
    .Q(\sine_out_reg1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _642_ (.CLK(clk),
    .D(\sine_out_temp1[13] ),
    .Q(\sine_out_reg1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _643_ (.CLK(clk),
    .D(\sine_out_temp1[14] ),
    .Q(\sine_out_reg1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _644_ (.CLK(clk),
    .D(\sine_out_temp1[15] ),
    .Q(\sine_out_reg1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _645_ (.CLK(clk),
    .D(\tcout_delay[1] ),
    .Q(\tcout_delay[0] ));
 sky130_fd_sc_hd__dfxtp_2 _646_ (.CLK(clk),
    .D(\tcout[8] ),
    .Q(\tcout_delay[1] ));
 sky130_fd_sc_hd__conb_1 _647_ (.HI(_291_));
 sky130_fd_sc_hd__conb_1 _648_ (.HI(_292_));
 sky130_fd_sc_hd__conb_1 _649_ (.HI(_293_));
 sky130_fd_sc_hd__conb_1 _650_ (.HI(_294_));
 sky130_fd_sc_hd__conb_1 _651_ (.LO(_295_));
 sky130_fd_sc_hd__conb_1 _652_ (.LO(_296_));
 sky130_sram_1kbyte_1rw1r_32x256_8 mem_i (.csb0(csb00),
    .csb1(_295_),
    .web0(_296_),
    .clk0(clk),
    .clk1(clk),
    .addr0({addr00[7],
    addr00[6],
    addr00[5],
    addr00[4],
    addr00[3],
    addr00[2],
    addr00[1],
    addr00[0]}),
    .addr1({\tcout[7] ,
    \tcout[6] ,
    \tcout[5] ,
    \tcout[4] ,
    \tcout[3] ,
    \tcout[2] ,
    \tcout[1] ,
    \tcout[0] }),
    .din0({din01[15],
    din01[14],
    din01[13],
    din01[12],
    din01[11],
    din01[10],
    din01[9],
    din01[8],
    din01[7],
    din01[6],
    din01[5],
    din01[4],
    din01[3],
    din01[2],
    din01[1],
    din01[0],
    din00[15],
    din00[14],
    din00[13],
    din00[12],
    din00[11],
    din00[10],
    din00[9],
    din00[8],
    din00[7],
    din00[6],
    din00[5],
    din00[4],
    din00[3],
    din00[2],
    din00[1],
    din00[0]}),
    .dout0({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .dout1({\sine_out_temp1[15] ,
    \sine_out_temp1[14] ,
    \sine_out_temp1[13] ,
    \sine_out_temp1[12] ,
    \sine_out_temp1[11] ,
    \sine_out_temp1[10] ,
    \sine_out_temp1[9] ,
    \sine_out_temp1[8] ,
    \sine_out_temp1[7] ,
    \sine_out_temp1[6] ,
    \sine_out_temp1[5] ,
    \sine_out_temp1[4] ,
    \sine_out_temp1[3] ,
    \sine_out_temp1[2] ,
    \sine_out_temp1[1] ,
    \sine_out_temp1[0] ,
    \sine_out_temp0[15] ,
    \sine_out_temp0[14] ,
    \sine_out_temp0[13] ,
    \sine_out_temp0[12] ,
    \sine_out_temp0[11] ,
    \sine_out_temp0[10] ,
    \sine_out_temp0[9] ,
    \sine_out_temp0[8] ,
    \sine_out_temp0[7] ,
    \sine_out_temp0[6] ,
    \sine_out_temp0[5] ,
    \sine_out_temp0[4] ,
    \sine_out_temp0[3] ,
    \sine_out_temp0[2] ,
    \sine_out_temp0[1] ,
    \sine_out_temp0[0] }),
    .wmask0({_294_,
    _293_,
    _292_,
    _291_}));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_2_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_2_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_2_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_2_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_2_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_2_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_2_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_2_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_2_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_2_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_2_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_2_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_2_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_2_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_2_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_2_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_2_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_2_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_2_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_2_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_2_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_2_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_2_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_2_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_2_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_2_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_2_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_2_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_2_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_2_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_2_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_1_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_1_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_1_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_1_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_1_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_1_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_1_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_1_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_1_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_1_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_1_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_1_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_1_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_1_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_1_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_1_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_1_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_1_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_1_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_1_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_1_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_1_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_1_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_1_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_1_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_1_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_1_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_1_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_1_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_1_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_1_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_1_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_1_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_1_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_1_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_1_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_1_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_1_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_1_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_1_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_1_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_1_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_1_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_1_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_1_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_1_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_1_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_1_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Left_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Left_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Left_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Left_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_2_Left_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_2_Left_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_2_Left_459 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_2_Left_460 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_2_Left_461 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_2_Left_462 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_2_Left_463 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_2_Left_464 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_2_Left_465 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_2_Left_466 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_2_Left_467 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_2_Left_468 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_2_Left_469 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_2_Left_470 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_2_Left_471 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_2_Left_472 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_2_Left_473 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_2_Left_474 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_2_Left_475 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_2_Left_476 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_2_Left_477 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_2_Left_478 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Left_479 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Left_480 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Left_481 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Left_482 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Left_483 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Left_484 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Left_485 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Left_486 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Left_487 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Left_488 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Left_489 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Left_490 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Left_491 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Left_492 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Left_493 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Left_494 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Left_495 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_2_Left_496 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_2_Left_497 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_2_Left_498 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_2_Left_499 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_2_Left_500 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_2_Left_501 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_2_Left_502 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_2_Left_503 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_2_Left_504 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_505 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_506 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_507 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_508 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_509 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_510 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_511 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_512 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_513 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_514 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_515 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_516 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_517 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_518 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_519 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_520 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_521 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_522 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_523 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_524 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_525 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_526 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_527 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_528 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_529 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_530 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_531 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_532 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_533 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_534 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_535 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_536 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_537 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_538 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_539 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_540 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_541 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_542 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_543 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_544 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_545 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_546 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_547 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_548 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_549 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_550 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_551 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_552 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_553 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_554 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_555 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_556 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_557 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_558 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_559 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_560 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_561 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_562 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_563 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Right_564 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Right_565 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Right_566 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Right_567 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Right_568 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Right_569 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Right_570 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Right_571 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Right_572 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Right_573 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Right_574 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Right_575 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Right_576 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Right_577 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Right_578 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Right_579 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Right_580 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Right_581 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Right_582 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Right_583 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Right_584 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Right_585 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Right_586 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Right_587 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Right_588 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Right_589 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Right_590 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Right_591 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Right_592 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Right_593 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Right_594 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Right_595 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Right_596 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Right_597 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Right_598 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Right_599 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Right_600 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Right_601 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Right_602 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Right_603 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Right_604 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Right_605 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Right_606 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Right_607 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Right_608 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Right_609 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Right_610 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_1_Right_611 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_1_Right_612 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_1_Right_613 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_1_Right_614 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_1_Right_615 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_1_Right_616 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_1_Right_617 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_1_Right_618 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_1_Right_619 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_1_Right_620 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_1_Right_621 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_1_Right_622 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_1_Right_623 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_1_Right_624 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_1_Right_625 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_1_Right_626 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_1_Right_627 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_1_Right_628 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_1_Right_629 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_1_Right_630 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_1_Right_631 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_1_Right_632 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_1_Right_633 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_1_Right_634 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_1_Right_635 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_1_Right_636 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_1_Right_637 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_1_Right_638 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_1_Right_639 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_1_Right_640 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_1_Right_641 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_1_Right_642 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_1_Right_643 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_1_Right_644 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_1_Right_645 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_1_Right_646 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_1_Right_647 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_1_Right_648 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_1_Right_649 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_1_Right_650 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_1_Right_651 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_1_Right_652 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_1_Right_653 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_1_Right_654 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_1_Right_655 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_1_Right_656 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_1_Right_657 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_1_Right_658 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_2_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_2_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_2_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2_1664 ();
endmodule
