magic
tech sky130A
magscale 1 2
timestamp 1740921364
<< checkpaint >>
rect -3932 -3932 23544 25688
<< viali >>
rect 8493 18921 8527 18955
rect 10149 18921 10183 18955
rect 11897 18921 11931 18955
rect 8309 18717 8343 18751
rect 9965 18717 9999 18751
rect 11713 18717 11747 18751
rect 14657 18717 14691 18751
rect 7757 18649 7791 18683
rect 8125 18649 8159 18683
rect 9597 18649 9631 18683
rect 9781 18649 9815 18683
rect 14749 18581 14783 18615
rect 7849 18377 7883 18411
rect 8033 18377 8067 18411
rect 9413 18377 9447 18411
rect 13277 18377 13311 18411
rect 11897 18309 11931 18343
rect 2329 18241 2363 18275
rect 3801 18241 3835 18275
rect 7113 18241 7147 18275
rect 7297 18241 7331 18275
rect 7852 18241 7886 18275
rect 8493 18241 8527 18275
rect 8769 18241 8803 18275
rect 8953 18241 8987 18275
rect 9587 18241 9621 18275
rect 9873 18241 9907 18275
rect 10425 18241 10459 18275
rect 10701 18241 10735 18275
rect 10885 18241 10919 18275
rect 12541 18241 12575 18275
rect 13001 18241 13035 18275
rect 13185 18241 13219 18275
rect 15301 18241 15335 18275
rect 15761 18241 15795 18275
rect 15945 18241 15979 18275
rect 16313 18241 16347 18275
rect 16405 18241 16439 18275
rect 16681 18241 16715 18275
rect 7205 18173 7239 18207
rect 7389 18173 7423 18207
rect 8309 18173 8343 18207
rect 8401 18173 8435 18207
rect 8585 18173 8619 18207
rect 10057 18173 10091 18207
rect 10241 18173 10275 18207
rect 10333 18173 10367 18207
rect 10517 18173 10551 18207
rect 12633 18173 12667 18207
rect 14749 18173 14783 18207
rect 15025 18173 15059 18207
rect 15209 18173 15243 18207
rect 7481 18105 7515 18139
rect 8125 18105 8159 18139
rect 9689 18105 9723 18139
rect 9781 18105 9815 18139
rect 12909 18105 12943 18139
rect 13185 18105 13219 18139
rect 15669 18105 15703 18139
rect 2237 18037 2271 18071
rect 3617 18037 3651 18071
rect 10793 18037 10827 18071
rect 11989 18037 12023 18071
rect 16773 18037 16807 18071
rect 7113 17833 7147 17867
rect 7665 17833 7699 17867
rect 10057 17833 10091 17867
rect 10793 17833 10827 17867
rect 11345 17833 11379 17867
rect 12817 17833 12851 17867
rect 13001 17833 13035 17867
rect 13093 17833 13127 17867
rect 13829 17833 13863 17867
rect 8401 17765 8435 17799
rect 12357 17765 12391 17799
rect 10701 17697 10735 17731
rect 11161 17697 11195 17731
rect 11989 17697 12023 17731
rect 14381 17697 14415 17731
rect 15945 17697 15979 17731
rect 16221 17697 16255 17731
rect 1685 17629 1719 17663
rect 3893 17629 3927 17663
rect 4077 17629 4111 17663
rect 5181 17629 5215 17663
rect 7297 17629 7331 17663
rect 7573 17629 7607 17663
rect 7849 17629 7883 17663
rect 7941 17629 7975 17663
rect 8217 17629 8251 17663
rect 8309 17629 8343 17663
rect 8677 17629 8711 17663
rect 9229 17629 9263 17663
rect 9505 17629 9539 17663
rect 10241 17629 10275 17663
rect 10425 17629 10459 17663
rect 10517 17629 10551 17663
rect 10885 17629 10919 17663
rect 10977 17629 11011 17663
rect 11069 17629 11103 17663
rect 11253 17629 11287 17663
rect 11529 17629 11563 17663
rect 12081 17629 12115 17663
rect 12357 17629 12391 17663
rect 13369 17629 13403 17663
rect 13921 17629 13955 17663
rect 14105 17629 14139 17663
rect 12863 17595 12897 17629
rect 3433 17561 3467 17595
rect 3617 17561 3651 17595
rect 8033 17561 8067 17595
rect 8401 17561 8435 17595
rect 9689 17561 9723 17595
rect 11621 17561 11655 17595
rect 11713 17561 11747 17595
rect 11831 17561 11865 17595
rect 12633 17561 12667 17595
rect 13093 17561 13127 17595
rect 1501 17493 1535 17527
rect 3249 17493 3283 17527
rect 4077 17493 4111 17527
rect 4997 17493 5031 17527
rect 7481 17493 7515 17527
rect 8585 17493 8619 17527
rect 9321 17493 9355 17527
rect 12173 17493 12207 17527
rect 13277 17493 13311 17527
rect 15853 17493 15887 17527
rect 17693 17493 17727 17527
rect 7665 17289 7699 17323
rect 8309 17289 8343 17323
rect 9689 17289 9723 17323
rect 12265 17289 12299 17323
rect 17785 17289 17819 17323
rect 2605 17221 2639 17255
rect 7849 17221 7883 17255
rect 8585 17221 8619 17255
rect 14749 17221 14783 17255
rect 1869 17153 1903 17187
rect 3341 17153 3375 17187
rect 3433 17153 3467 17187
rect 3525 17153 3559 17187
rect 3709 17153 3743 17187
rect 4629 17153 4663 17187
rect 4813 17153 4847 17187
rect 5733 17153 5767 17187
rect 6929 17153 6963 17187
rect 7113 17153 7147 17187
rect 7205 17153 7239 17187
rect 7757 17153 7791 17187
rect 7941 17153 7975 17187
rect 8493 17153 8527 17187
rect 8677 17153 8711 17187
rect 8861 17153 8895 17187
rect 8953 17153 8987 17187
rect 9045 17153 9079 17187
rect 9193 17153 9227 17187
rect 9321 17153 9355 17187
rect 9413 17153 9447 17187
rect 9551 17153 9585 17187
rect 10149 17153 10183 17187
rect 10241 17153 10275 17187
rect 10425 17153 10459 17187
rect 11713 17153 11747 17187
rect 11805 17153 11839 17187
rect 11989 17153 12023 17187
rect 12081 17153 12115 17187
rect 14105 17153 14139 17187
rect 14565 17153 14599 17187
rect 16497 17153 16531 17187
rect 16681 17153 16715 17187
rect 17693 17153 17727 17187
rect 2145 17085 2179 17119
rect 7481 17085 7515 17119
rect 7573 17085 7607 17119
rect 9965 17085 9999 17119
rect 10057 17085 10091 17119
rect 16957 17085 16991 17119
rect 2421 17017 2455 17051
rect 9781 17017 9815 17051
rect 1685 16949 1719 16983
rect 2053 16949 2087 16983
rect 3065 16949 3099 16983
rect 4997 16949 5031 16983
rect 5641 16949 5675 16983
rect 6929 16949 6963 16983
rect 7297 16949 7331 16983
rect 10609 16949 10643 16983
rect 13921 16949 13955 16983
rect 14473 16949 14507 16983
rect 1501 16745 1535 16779
rect 3433 16745 3467 16779
rect 4445 16745 4479 16779
rect 7389 16745 7423 16779
rect 9229 16745 9263 16779
rect 9597 16745 9631 16779
rect 10425 16745 10459 16779
rect 11621 16745 11655 16779
rect 11989 16745 12023 16779
rect 12817 16745 12851 16779
rect 14841 16745 14875 16779
rect 15742 16745 15776 16779
rect 17233 16745 17267 16779
rect 2789 16677 2823 16711
rect 2881 16677 2915 16711
rect 7021 16677 7055 16711
rect 14749 16677 14783 16711
rect 14933 16677 14967 16711
rect 2145 16609 2179 16643
rect 3801 16609 3835 16643
rect 6285 16609 6319 16643
rect 11805 16609 11839 16643
rect 11897 16609 11931 16643
rect 14381 16609 14415 16643
rect 15485 16609 15519 16643
rect 1869 16541 1903 16575
rect 1961 16541 1995 16575
rect 2697 16541 2731 16575
rect 2973 16541 3007 16575
rect 3157 16541 3191 16575
rect 3524 16541 3558 16575
rect 3617 16541 3651 16575
rect 3985 16541 4019 16575
rect 4261 16541 4295 16575
rect 4353 16541 4387 16575
rect 4808 16541 4842 16575
rect 5125 16541 5159 16575
rect 5273 16541 5307 16575
rect 5917 16541 5951 16575
rect 6193 16541 6227 16575
rect 6653 16541 6687 16575
rect 6745 16541 6779 16575
rect 6929 16541 6963 16575
rect 7113 16541 7147 16575
rect 7205 16541 7239 16575
rect 9321 16541 9355 16575
rect 9505 16541 9539 16575
rect 9689 16541 9723 16575
rect 10057 16541 10091 16575
rect 10149 16541 10183 16575
rect 10425 16541 10459 16575
rect 11529 16541 11563 16575
rect 12081 16541 12115 16575
rect 12173 16541 12207 16575
rect 13093 16541 13127 16575
rect 13185 16541 13219 16575
rect 13277 16541 13311 16575
rect 13461 16541 13495 16575
rect 15117 16541 15151 16575
rect 15393 16541 15427 16575
rect 17509 16541 17543 16575
rect 4169 16473 4203 16507
rect 4905 16473 4939 16507
rect 4997 16473 5031 16507
rect 6469 16473 6503 16507
rect 7481 16473 7515 16507
rect 7849 16473 7883 16507
rect 8033 16473 8067 16507
rect 8217 16473 8251 16507
rect 9781 16473 9815 16507
rect 17417 16473 17451 16507
rect 2513 16405 2547 16439
rect 4629 16405 4663 16439
rect 9879 16405 9913 16439
rect 9965 16405 9999 16439
rect 10241 16405 10275 16439
rect 11805 16405 11839 16439
rect 15301 16405 15335 16439
rect 1961 16201 1995 16235
rect 2513 16201 2547 16235
rect 10793 16201 10827 16235
rect 11345 16201 11379 16235
rect 11529 16201 11563 16235
rect 13093 16201 13127 16235
rect 14105 16201 14139 16235
rect 7205 16133 7239 16167
rect 10885 16133 10919 16167
rect 13645 16133 13679 16167
rect 13829 16133 13863 16167
rect 14473 16133 14507 16167
rect 16865 16133 16899 16167
rect 17693 16133 17727 16167
rect 14243 16099 14277 16133
rect 1869 16065 1903 16099
rect 2697 16065 2731 16099
rect 2973 16065 3007 16099
rect 4169 16065 4203 16099
rect 4261 16065 4295 16099
rect 4445 16065 4479 16099
rect 4537 16065 4571 16099
rect 5181 16065 5215 16099
rect 5733 16065 5767 16099
rect 5917 16065 5951 16099
rect 6377 16065 6411 16099
rect 6929 16065 6963 16099
rect 7021 16065 7055 16099
rect 7389 16065 7423 16099
rect 9137 16065 9171 16099
rect 9505 16065 9539 16099
rect 9781 16065 9815 16099
rect 10149 16065 10183 16099
rect 10242 16065 10276 16099
rect 10425 16065 10459 16099
rect 10517 16065 10551 16099
rect 10614 16065 10648 16099
rect 11161 16065 11195 16099
rect 11805 16065 11839 16099
rect 11897 16065 11931 16099
rect 11989 16065 12023 16099
rect 12449 16065 12483 16099
rect 13277 16065 13311 16099
rect 13461 16065 13495 16099
rect 13553 16065 13587 16099
rect 14657 16065 14691 16099
rect 15669 16065 15703 16099
rect 15945 16065 15979 16099
rect 16037 16065 16071 16099
rect 17509 16065 17543 16099
rect 2145 15997 2179 16031
rect 2789 15997 2823 16031
rect 2881 15997 2915 16031
rect 11069 15997 11103 16031
rect 11713 15997 11747 16031
rect 12173 15997 12207 16031
rect 17325 15997 17359 16031
rect 5733 15929 5767 15963
rect 6837 15929 6871 15963
rect 7573 15929 7607 15963
rect 12633 15929 12667 15963
rect 17233 15929 17267 15963
rect 1501 15861 1535 15895
rect 3985 15861 4019 15895
rect 9321 15861 9355 15895
rect 9873 15861 9907 15895
rect 10057 15861 10091 15895
rect 11161 15861 11195 15895
rect 12265 15861 12299 15895
rect 14013 15861 14047 15895
rect 14289 15861 14323 15895
rect 14933 15861 14967 15895
rect 16221 15861 16255 15895
rect 16681 15861 16715 15895
rect 16865 15861 16899 15895
rect 1501 15657 1535 15691
rect 3525 15657 3559 15691
rect 4261 15657 4295 15691
rect 5457 15657 5491 15691
rect 8033 15657 8067 15691
rect 9781 15657 9815 15691
rect 10241 15657 10275 15691
rect 10425 15657 10459 15691
rect 12173 15657 12207 15691
rect 15853 15657 15887 15691
rect 6561 15589 6595 15623
rect 3617 15521 3651 15555
rect 5089 15521 5123 15555
rect 6193 15521 6227 15555
rect 6285 15521 6319 15555
rect 9321 15521 9355 15555
rect 9505 15521 9539 15555
rect 12265 15521 12299 15555
rect 1685 15453 1719 15487
rect 2237 15453 2271 15487
rect 2789 15453 2823 15487
rect 2973 15453 3007 15487
rect 3065 15453 3099 15487
rect 3341 15453 3375 15487
rect 3433 15453 3467 15487
rect 4169 15453 4203 15487
rect 4353 15453 4387 15487
rect 5181 15453 5215 15487
rect 5549 15453 5583 15487
rect 5641 15453 5675 15487
rect 5825 15453 5859 15487
rect 6837 15453 6871 15487
rect 7021 15453 7055 15487
rect 7481 15453 7515 15487
rect 7573 15453 7607 15487
rect 7757 15453 7791 15487
rect 7849 15453 7883 15487
rect 8493 15453 8527 15487
rect 9413 15453 9447 15487
rect 9597 15453 9631 15487
rect 11529 15453 11563 15487
rect 11713 15453 11747 15487
rect 11805 15453 11839 15487
rect 11897 15453 11931 15487
rect 12449 15453 12483 15487
rect 12725 15453 12759 15487
rect 13921 15453 13955 15487
rect 14105 15453 14139 15487
rect 15945 15453 15979 15487
rect 6101 15385 6135 15419
rect 10057 15385 10091 15419
rect 14381 15385 14415 15419
rect 16221 15385 16255 15419
rect 2053 15317 2087 15351
rect 6745 15317 6779 15351
rect 7021 15317 7055 15351
rect 8401 15317 8435 15351
rect 10257 15317 10291 15351
rect 12633 15317 12667 15351
rect 13829 15317 13863 15351
rect 17693 15317 17727 15351
rect 5181 15113 5215 15147
rect 5365 15113 5399 15147
rect 7849 15113 7883 15147
rect 9505 15113 9539 15147
rect 9689 15113 9723 15147
rect 10057 15113 10091 15147
rect 14105 15113 14139 15147
rect 14657 15113 14691 15147
rect 4721 15045 4755 15079
rect 8861 15045 8895 15079
rect 13277 15045 13311 15079
rect 1685 14977 1719 15011
rect 2697 14977 2731 15011
rect 2881 14977 2915 15011
rect 3525 14977 3559 15011
rect 3709 14977 3743 15011
rect 4537 14977 4571 15011
rect 5549 14977 5583 15011
rect 6561 14977 6595 15011
rect 7021 14977 7055 15011
rect 7205 14977 7239 15011
rect 8125 14977 8159 15011
rect 8401 14977 8435 15011
rect 8769 14977 8803 15011
rect 8953 14977 8987 15011
rect 9321 14977 9355 15011
rect 9505 14977 9539 15011
rect 9597 14977 9631 15011
rect 9781 14977 9815 15011
rect 10241 14977 10275 15011
rect 10333 14977 10367 15011
rect 10517 14977 10551 15011
rect 10609 14977 10643 15011
rect 13093 14977 13127 15011
rect 13553 14977 13587 15011
rect 14289 14977 14323 15011
rect 14565 14977 14599 15011
rect 15025 14977 15059 15011
rect 15853 14977 15887 15011
rect 16923 14977 16957 15011
rect 17325 14977 17359 15011
rect 6653 14909 6687 14943
rect 7849 14909 7883 14943
rect 8677 14909 8711 14943
rect 12909 14909 12943 14943
rect 13001 14909 13035 14943
rect 14473 14909 14507 14943
rect 15669 14909 15703 14943
rect 17233 14909 17267 14943
rect 5089 14841 5123 14875
rect 16681 14841 16715 14875
rect 1501 14773 1535 14807
rect 2881 14773 2915 14807
rect 3525 14773 3559 14807
rect 4261 14773 4295 14807
rect 6653 14773 6687 14807
rect 6929 14773 6963 14807
rect 7205 14773 7239 14807
rect 8033 14773 8067 14807
rect 8217 14773 8251 14807
rect 8585 14773 8619 14807
rect 13369 14773 13403 14807
rect 1593 14569 1627 14603
rect 3433 14569 3467 14603
rect 4721 14569 4755 14603
rect 6377 14569 6411 14603
rect 7389 14569 7423 14603
rect 7665 14569 7699 14603
rect 10057 14569 10091 14603
rect 10977 14569 11011 14603
rect 12081 14569 12115 14603
rect 14657 14569 14691 14603
rect 15761 14569 15795 14603
rect 17877 14569 17911 14603
rect 2145 14501 2179 14535
rect 5089 14501 5123 14535
rect 7573 14501 7607 14535
rect 8493 14501 8527 14535
rect 8585 14501 8619 14535
rect 12449 14501 12483 14535
rect 12633 14501 12667 14535
rect 14841 14501 14875 14535
rect 2053 14433 2087 14467
rect 3617 14433 3651 14467
rect 4169 14433 4203 14467
rect 6469 14433 6503 14467
rect 7205 14433 7239 14467
rect 8401 14433 8435 14467
rect 12909 14433 12943 14467
rect 1777 14365 1811 14399
rect 1961 14365 1995 14399
rect 2421 14365 2455 14399
rect 2789 14365 2823 14399
rect 2973 14365 3007 14399
rect 3157 14365 3191 14399
rect 3249 14365 3283 14399
rect 3341 14365 3375 14399
rect 3985 14365 4019 14399
rect 4077 14365 4111 14399
rect 4261 14365 4295 14399
rect 4445 14365 4479 14399
rect 6009 14365 6043 14399
rect 7389 14365 7423 14399
rect 7941 14365 7975 14399
rect 8033 14365 8067 14399
rect 8125 14365 8159 14399
rect 8309 14365 8343 14399
rect 8677 14365 8711 14399
rect 10241 14365 10275 14399
rect 10333 14365 10367 14399
rect 10425 14365 10459 14399
rect 10517 14365 10551 14399
rect 10701 14365 10735 14399
rect 10793 14365 10827 14399
rect 12265 14365 12299 14399
rect 12541 14365 12575 14399
rect 12633 14365 12667 14399
rect 12725 14365 12759 14399
rect 14565 14365 14599 14399
rect 17785 14365 17819 14399
rect 2145 14297 2179 14331
rect 2881 14297 2915 14331
rect 3801 14297 3835 14331
rect 4721 14297 4755 14331
rect 6929 14297 6963 14331
rect 9045 14297 9079 14331
rect 10977 14297 11011 14331
rect 15025 14297 15059 14331
rect 15209 14297 15243 14331
rect 17049 14297 17083 14331
rect 2329 14229 2363 14263
rect 2605 14229 2639 14263
rect 3617 14229 3651 14263
rect 4537 14229 4571 14263
rect 5733 14229 5767 14263
rect 6101 14229 6135 14263
rect 6193 14229 6227 14263
rect 9137 14229 9171 14263
rect 1961 14025 1995 14059
rect 2789 14025 2823 14059
rect 6101 14025 6135 14059
rect 6377 14025 6411 14059
rect 7481 14025 7515 14059
rect 8585 14025 8619 14059
rect 9965 14025 9999 14059
rect 11345 14025 11379 14059
rect 11621 14025 11655 14059
rect 11989 14025 12023 14059
rect 12909 14025 12943 14059
rect 14105 14025 14139 14059
rect 14289 14025 14323 14059
rect 15761 14025 15795 14059
rect 17785 14025 17819 14059
rect 1869 13957 1903 13991
rect 2421 13957 2455 13991
rect 2637 13957 2671 13991
rect 3709 13957 3743 13991
rect 6653 13957 6687 13991
rect 6745 13957 6779 13991
rect 8953 13957 8987 13991
rect 15393 13957 15427 13991
rect 18061 13957 18095 13991
rect 3065 13889 3099 13923
rect 3157 13889 3191 13923
rect 3341 13889 3375 13923
rect 3433 13889 3467 13923
rect 3893 13889 3927 13923
rect 4077 13889 4111 13923
rect 4261 13889 4295 13923
rect 4445 13889 4479 13923
rect 4905 13889 4939 13923
rect 5089 13889 5123 13923
rect 5917 13889 5951 13923
rect 6193 13889 6227 13923
rect 6556 13889 6590 13923
rect 6928 13889 6962 13923
rect 7021 13889 7055 13923
rect 7113 13889 7147 13923
rect 8769 13889 8803 13923
rect 9045 13889 9079 13923
rect 9597 13889 9631 13923
rect 9873 13889 9907 13923
rect 10057 13889 10091 13923
rect 10149 13889 10183 13923
rect 11069 13889 11103 13923
rect 11529 13889 11563 13923
rect 11713 13889 11747 13923
rect 12173 13889 12207 13923
rect 12449 13889 12483 13923
rect 12541 13889 12575 13923
rect 12725 13889 12759 13923
rect 12817 13889 12851 13923
rect 13001 13889 13035 13923
rect 14013 13889 14047 13923
rect 14381 13889 14415 13923
rect 15301 13889 15335 13923
rect 15485 13889 15519 13923
rect 15669 13889 15703 13923
rect 16773 13889 16807 13923
rect 17601 13889 17635 13923
rect 2145 13821 2179 13855
rect 4629 13821 4663 13855
rect 4997 13821 5031 13855
rect 5733 13821 5767 13855
rect 7205 13821 7239 13855
rect 10425 13821 10459 13855
rect 11345 13821 11379 13855
rect 12357 13821 12391 13855
rect 14197 13821 14231 13855
rect 2881 13753 2915 13787
rect 1501 13685 1535 13719
rect 2605 13685 2639 13719
rect 7297 13685 7331 13719
rect 9321 13685 9355 13719
rect 11161 13685 11195 13719
rect 17141 13685 17175 13719
rect 1501 13481 1535 13515
rect 2421 13481 2455 13515
rect 3801 13481 3835 13515
rect 6009 13481 6043 13515
rect 6377 13481 6411 13515
rect 8769 13481 8803 13515
rect 9505 13481 9539 13515
rect 13737 13481 13771 13515
rect 14105 13481 14139 13515
rect 6561 13413 6595 13447
rect 4445 13345 4479 13379
rect 8401 13345 8435 13379
rect 9321 13345 9355 13379
rect 10149 13345 10183 13379
rect 11069 13345 11103 13379
rect 13645 13345 13679 13379
rect 1685 13277 1719 13311
rect 2605 13277 2639 13311
rect 2881 13277 2915 13311
rect 4169 13277 4203 13311
rect 5917 13277 5951 13311
rect 6193 13277 6227 13311
rect 6745 13277 6779 13311
rect 8309 13277 8343 13311
rect 8493 13277 8527 13311
rect 8585 13277 8619 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9689 13277 9723 13311
rect 9873 13277 9907 13311
rect 10011 13277 10045 13311
rect 10793 13277 10827 13311
rect 12081 13277 12115 13311
rect 12357 13277 12391 13311
rect 12633 13277 12667 13311
rect 12817 13277 12851 13311
rect 13369 13277 13403 13311
rect 14381 13277 14415 13311
rect 14473 13277 14507 13311
rect 14565 13277 14599 13311
rect 14749 13277 14783 13311
rect 16405 13277 16439 13311
rect 2789 13209 2823 13243
rect 4261 13209 4295 13243
rect 9781 13209 9815 13243
rect 12449 13209 12483 13243
rect 11897 13141 11931 13175
rect 12265 13141 12299 13175
rect 13921 13141 13955 13175
rect 17693 13141 17727 13175
rect 6929 12937 6963 12971
rect 8585 12937 8619 12971
rect 13921 12937 13955 12971
rect 17141 12937 17175 12971
rect 3249 12869 3283 12903
rect 12817 12869 12851 12903
rect 15761 12869 15795 12903
rect 17509 12869 17543 12903
rect 3065 12801 3099 12835
rect 3341 12801 3375 12835
rect 4629 12801 4663 12835
rect 4905 12801 4939 12835
rect 4997 12801 5031 12835
rect 5181 12801 5215 12835
rect 6561 12801 6595 12835
rect 7113 12801 7147 12835
rect 8217 12801 8251 12835
rect 8401 12801 8435 12835
rect 8861 12801 8895 12835
rect 8953 12801 8987 12835
rect 9045 12801 9079 12835
rect 9229 12801 9263 12835
rect 10609 12801 10643 12835
rect 10793 12801 10827 12835
rect 10885 12801 10919 12835
rect 12725 12801 12759 12835
rect 12909 12801 12943 12835
rect 13185 12801 13219 12835
rect 13277 12801 13311 12835
rect 13369 12801 13403 12835
rect 13737 12801 13771 12835
rect 14013 12801 14047 12835
rect 14197 12801 14231 12835
rect 14381 12801 14415 12835
rect 14473 12801 14507 12835
rect 14657 12801 14691 12835
rect 14749 12801 14783 12835
rect 15209 12801 15243 12835
rect 16681 12801 16715 12835
rect 16957 12801 16991 12835
rect 17325 12801 17359 12835
rect 17877 12801 17911 12835
rect 4537 12733 4571 12767
rect 6653 12733 6687 12767
rect 13093 12733 13127 12767
rect 15301 12733 15335 12767
rect 15393 12733 15427 12767
rect 3065 12665 3099 12699
rect 8309 12665 8343 12699
rect 10425 12665 10459 12699
rect 13553 12665 13587 12699
rect 5181 12597 5215 12631
rect 6561 12597 6595 12631
rect 7297 12597 7331 12631
rect 13737 12597 13771 12631
rect 14841 12597 14875 12631
rect 15853 12597 15887 12631
rect 16773 12597 16807 12631
rect 18061 12597 18095 12631
rect 2421 12393 2455 12427
rect 3801 12393 3835 12427
rect 7481 12393 7515 12427
rect 8125 12393 8159 12427
rect 10977 12393 11011 12427
rect 14657 12393 14691 12427
rect 15577 12393 15611 12427
rect 4629 12325 4663 12359
rect 6193 12325 6227 12359
rect 7297 12325 7331 12359
rect 11989 12325 12023 12359
rect 4537 12257 4571 12291
rect 9045 12257 9079 12291
rect 9137 12257 9171 12291
rect 9321 12257 9355 12291
rect 11345 12257 11379 12291
rect 11437 12257 11471 12291
rect 11805 12257 11839 12291
rect 2145 12189 2179 12223
rect 2283 12189 2317 12223
rect 2605 12189 2639 12223
rect 3985 12189 4019 12223
rect 4169 12189 4203 12223
rect 4287 12189 4321 12223
rect 4445 12189 4479 12223
rect 4721 12189 4755 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 5089 12189 5123 12223
rect 6377 12189 6411 12223
rect 6469 12189 6503 12223
rect 6597 12189 6631 12223
rect 6837 12189 6871 12223
rect 6929 12189 6963 12223
rect 7021 12189 7055 12223
rect 8033 12189 8067 12223
rect 8125 12189 8159 12223
rect 8309 12189 8343 12223
rect 9413 12189 9447 12223
rect 9525 12189 9559 12223
rect 9781 12189 9815 12223
rect 9873 12189 9907 12223
rect 11161 12189 11195 12223
rect 11529 12189 11563 12223
rect 11713 12189 11747 12223
rect 12081 12189 12115 12223
rect 12173 12189 12207 12223
rect 12357 12189 12391 12223
rect 12449 12189 12483 12223
rect 12909 12189 12943 12223
rect 13093 12189 13127 12223
rect 14381 12189 14415 12223
rect 14657 12189 14691 12223
rect 14841 12189 14875 12223
rect 14933 12189 14967 12223
rect 15301 12189 15335 12223
rect 15393 12189 15427 12223
rect 15945 12189 15979 12223
rect 16037 12189 16071 12223
rect 17877 12189 17911 12223
rect 4077 12121 4111 12155
rect 4997 12121 5031 12155
rect 6193 12121 6227 12155
rect 7205 12121 7239 12155
rect 7449 12121 7483 12155
rect 7665 12121 7699 12155
rect 8953 12121 8987 12155
rect 9689 12121 9723 12155
rect 11805 12121 11839 12155
rect 12587 12121 12621 12155
rect 12725 12121 12759 12155
rect 12817 12121 12851 12155
rect 15025 12121 15059 12155
rect 16313 12121 16347 12155
rect 2605 12053 2639 12087
rect 7849 12053 7883 12087
rect 10057 12053 10091 12087
rect 12357 12053 12391 12087
rect 15761 12053 15795 12087
rect 17785 12053 17819 12087
rect 17969 12053 18003 12087
rect 1961 11849 1995 11883
rect 2329 11849 2363 11883
rect 4077 11849 4111 11883
rect 5549 11849 5583 11883
rect 6561 11849 6595 11883
rect 9781 11849 9815 11883
rect 11805 11849 11839 11883
rect 12725 11849 12759 11883
rect 15393 11849 15427 11883
rect 15853 11849 15887 11883
rect 2697 11781 2731 11815
rect 15209 11781 15243 11815
rect 1869 11713 1903 11747
rect 2508 11713 2542 11747
rect 2605 11713 2639 11747
rect 2825 11713 2859 11747
rect 2973 11713 3007 11747
rect 4169 11713 4203 11747
rect 4261 11713 4295 11747
rect 4537 11713 4571 11747
rect 4992 11713 5026 11747
rect 5089 11713 5123 11747
rect 5181 11713 5215 11747
rect 5364 11713 5398 11747
rect 5457 11713 5491 11747
rect 5733 11713 5767 11747
rect 5917 11713 5951 11747
rect 6009 11713 6043 11747
rect 6377 11713 6411 11747
rect 6653 11713 6687 11747
rect 6929 11713 6963 11747
rect 7113 11713 7147 11747
rect 7389 11713 7423 11747
rect 9965 11713 9999 11747
rect 10057 11713 10091 11747
rect 10149 11713 10183 11747
rect 11529 11713 11563 11747
rect 12817 11713 12851 11747
rect 13185 11713 13219 11747
rect 13277 11713 13311 11747
rect 13369 11713 13403 11747
rect 13553 11713 13587 11747
rect 15485 11713 15519 11747
rect 16221 11713 16255 11747
rect 16681 11713 16715 11747
rect 17785 11713 17819 11747
rect 2053 11645 2087 11679
rect 10241 11645 10275 11679
rect 11621 11645 11655 11679
rect 11805 11645 11839 11679
rect 12909 11645 12943 11679
rect 13737 11645 13771 11679
rect 15853 11645 15887 11679
rect 15945 11645 15979 11679
rect 17509 11645 17543 11679
rect 4445 11577 4479 11611
rect 6377 11577 6411 11611
rect 7205 11577 7239 11611
rect 7297 11577 7331 11611
rect 15209 11577 15243 11611
rect 1501 11509 1535 11543
rect 4813 11509 4847 11543
rect 7573 11509 7607 11543
rect 13093 11509 13127 11543
rect 16129 11509 16163 11543
rect 16865 11509 16899 11543
rect 1501 11305 1535 11339
rect 1961 11305 1995 11339
rect 2145 11305 2179 11339
rect 4261 11305 4295 11339
rect 4445 11305 4479 11339
rect 7757 11305 7791 11339
rect 7941 11305 7975 11339
rect 13461 11305 13495 11339
rect 2789 11237 2823 11271
rect 4077 11237 4111 11271
rect 7389 11237 7423 11271
rect 8401 11237 8435 11271
rect 9045 11237 9079 11271
rect 14565 11237 14599 11271
rect 15025 11237 15059 11271
rect 2053 11169 2087 11203
rect 4629 11169 4663 11203
rect 6929 11169 6963 11203
rect 9137 11169 9171 11203
rect 13093 11169 13127 11203
rect 13185 11169 13219 11203
rect 13645 11169 13679 11203
rect 14657 11169 14691 11203
rect 16405 11169 16439 11203
rect 18153 11169 18187 11203
rect 1685 11101 1719 11135
rect 2513 11101 2547 11135
rect 2605 11101 2639 11135
rect 3801 11101 3835 11135
rect 4445 11101 4479 11135
rect 4813 11101 4847 11135
rect 7113 11101 7147 11135
rect 8125 11101 8159 11135
rect 8310 11101 8344 11135
rect 8493 11101 8527 11135
rect 8585 11101 8619 11135
rect 8953 11101 8987 11135
rect 9413 11101 9447 11135
rect 10057 11101 10091 11135
rect 10241 11101 10275 11135
rect 10333 11101 10367 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 13001 11101 13035 11135
rect 13277 11101 13311 11135
rect 13553 11101 13587 11135
rect 13737 11101 13771 11135
rect 14381 11101 14415 11135
rect 14749 11101 14783 11135
rect 14841 11101 14875 11135
rect 15025 11101 15059 11135
rect 15485 11101 15519 11135
rect 16313 11101 16347 11135
rect 2421 11033 2455 11067
rect 2789 11033 2823 11067
rect 4721 11033 4755 11067
rect 7481 11033 7515 11067
rect 7573 11033 7607 11067
rect 16681 11033 16715 11067
rect 2329 10965 2363 10999
rect 7773 10965 7807 10999
rect 8769 10965 8803 10999
rect 9229 10965 9263 10999
rect 9321 10965 9355 10999
rect 14197 10965 14231 10999
rect 15669 10965 15703 10999
rect 16129 10965 16163 10999
rect 3709 10761 3743 10795
rect 4905 10761 4939 10795
rect 5365 10761 5399 10795
rect 5641 10761 5675 10795
rect 14749 10761 14783 10795
rect 15301 10761 15335 10795
rect 15669 10761 15703 10795
rect 16681 10761 16715 10795
rect 7021 10693 7055 10727
rect 8125 10693 8159 10727
rect 11989 10693 12023 10727
rect 15025 10693 15059 10727
rect 17417 10693 17451 10727
rect 3525 10625 3559 10659
rect 3801 10625 3835 10659
rect 3893 10625 3927 10659
rect 4077 10625 4111 10659
rect 4169 10625 4203 10659
rect 4261 10625 4295 10659
rect 5549 10625 5583 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 6653 10625 6687 10659
rect 7838 10625 7872 10659
rect 7997 10625 8031 10659
rect 8217 10625 8251 10659
rect 8355 10625 8389 10659
rect 8861 10625 8895 10659
rect 11779 10625 11813 10659
rect 11897 10625 11931 10659
rect 12081 10625 12115 10659
rect 12265 10625 12299 10659
rect 13921 10625 13955 10659
rect 14013 10625 14047 10659
rect 14749 10625 14783 10659
rect 14933 10625 14967 10659
rect 15209 10625 15243 10659
rect 15393 10625 15427 10659
rect 15853 10625 15887 10659
rect 15945 10625 15979 10659
rect 16129 10625 16163 10659
rect 16221 10625 16255 10659
rect 16957 10625 16991 10659
rect 17049 10625 17083 10659
rect 17141 10625 17175 10659
rect 17325 10625 17359 10659
rect 17693 10625 17727 10659
rect 18153 10625 18187 10659
rect 5089 10557 5123 10591
rect 5181 10557 5215 10591
rect 5457 10557 5491 10591
rect 6561 10557 6595 10591
rect 6929 10557 6963 10591
rect 8585 10557 8619 10591
rect 8769 10557 8803 10591
rect 11621 10557 11655 10591
rect 15577 10557 15611 10591
rect 17509 10557 17543 10591
rect 8493 10489 8527 10523
rect 17877 10489 17911 10523
rect 17969 10489 18003 10523
rect 3341 10421 3375 10455
rect 4537 10421 4571 10455
rect 6377 10421 6411 10455
rect 8677 10421 8711 10455
rect 14105 10421 14139 10455
rect 14289 10421 14323 10455
rect 17417 10421 17451 10455
rect 9413 10217 9447 10251
rect 11437 10217 11471 10251
rect 12081 10217 12115 10251
rect 15577 10217 15611 10251
rect 16405 10217 16439 10251
rect 17693 10217 17727 10251
rect 6101 10149 6135 10183
rect 10057 10081 10091 10115
rect 10885 10081 10919 10115
rect 1685 10013 1719 10047
rect 3985 10013 4019 10047
rect 4077 10013 4111 10047
rect 4261 10013 4295 10047
rect 4353 10013 4387 10047
rect 5457 10013 5491 10047
rect 5550 10013 5584 10047
rect 5825 10013 5859 10047
rect 5963 10013 5997 10047
rect 7113 10013 7147 10047
rect 7205 10013 7239 10047
rect 7481 10013 7515 10047
rect 7573 10013 7607 10047
rect 8125 10013 8159 10047
rect 8401 10013 8435 10047
rect 9689 10013 9723 10047
rect 9781 10013 9815 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 10517 10013 10551 10047
rect 10793 10013 10827 10047
rect 10977 10013 11011 10047
rect 11345 10013 11379 10047
rect 11529 10013 11563 10047
rect 11989 10013 12023 10047
rect 12173 10013 12207 10047
rect 15393 10013 15427 10047
rect 15547 10013 15581 10047
rect 16497 10013 16531 10047
rect 16865 10013 16899 10047
rect 17049 10013 17083 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 17509 10013 17543 10047
rect 17877 10013 17911 10047
rect 17969 10013 18003 10047
rect 5733 9945 5767 9979
rect 6285 9945 6319 9979
rect 7389 9945 7423 9979
rect 7941 9945 7975 9979
rect 9873 9945 9907 9979
rect 10701 9945 10735 9979
rect 16037 9945 16071 9979
rect 16221 9945 16255 9979
rect 17141 9945 17175 9979
rect 17693 9945 17727 9979
rect 1501 9877 1535 9911
rect 3801 9877 3835 9911
rect 7757 9877 7791 9911
rect 8309 9877 8343 9911
rect 10333 9877 10367 9911
rect 16865 9877 16899 9911
rect 1501 9673 1535 9707
rect 5365 9673 5399 9707
rect 6377 9673 6411 9707
rect 9321 9673 9355 9707
rect 2329 9605 2363 9639
rect 3433 9605 3467 9639
rect 3985 9605 4019 9639
rect 17693 9605 17727 9639
rect 17877 9605 17911 9639
rect 3755 9571 3789 9605
rect 1869 9537 1903 9571
rect 1961 9537 1995 9571
rect 2513 9537 2547 9571
rect 2697 9537 2731 9571
rect 2789 9537 2823 9571
rect 3065 9537 3099 9571
rect 3157 9537 3191 9571
rect 4905 9537 4939 9571
rect 4997 9537 5031 9571
rect 5549 9537 5583 9571
rect 6009 9537 6043 9571
rect 6205 9537 6239 9571
rect 6561 9537 6595 9571
rect 7205 9537 7239 9571
rect 7481 9537 7515 9571
rect 7573 9537 7607 9571
rect 7757 9537 7791 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 9045 9537 9079 9571
rect 9597 9537 9631 9571
rect 9873 9537 9907 9571
rect 9965 9537 9999 9571
rect 11069 9537 11103 9571
rect 11253 9537 11287 9571
rect 12541 9537 12575 9571
rect 12737 9537 12771 9571
rect 13001 9537 13035 9571
rect 13185 9537 13219 9571
rect 13461 9537 13495 9571
rect 13737 9537 13771 9571
rect 13918 9537 13952 9571
rect 14381 9537 14415 9571
rect 17417 9537 17451 9571
rect 2145 9469 2179 9503
rect 3525 9469 3559 9503
rect 5181 9469 5215 9503
rect 6653 9469 6687 9503
rect 6745 9469 6779 9503
rect 6837 9469 6871 9503
rect 7297 9469 7331 9503
rect 8953 9469 8987 9503
rect 10057 9469 10091 9503
rect 10149 9469 10183 9503
rect 13553 9469 13587 9503
rect 13645 9469 13679 9503
rect 14289 9469 14323 9503
rect 16865 9469 16899 9503
rect 17509 9469 17543 9503
rect 3617 9401 3651 9435
rect 6009 9401 6043 9435
rect 11069 9401 11103 9435
rect 14013 9401 14047 9435
rect 17141 9401 17175 9435
rect 2881 9333 2915 9367
rect 3801 9333 3835 9367
rect 7849 9333 7883 9367
rect 9689 9333 9723 9367
rect 12725 9333 12759 9367
rect 12909 9333 12943 9367
rect 13277 9333 13311 9367
rect 14289 9333 14323 9367
rect 1685 9129 1719 9163
rect 2237 9129 2271 9163
rect 3433 9129 3467 9163
rect 3893 9129 3927 9163
rect 5181 9129 5215 9163
rect 5641 9129 5675 9163
rect 9045 9129 9079 9163
rect 11069 9129 11103 9163
rect 16773 9129 16807 9163
rect 17049 9129 17083 9163
rect 3295 9061 3329 9095
rect 6929 9061 6963 9095
rect 9597 9061 9631 9095
rect 11437 9061 11471 9095
rect 11713 9061 11747 9095
rect 11805 9061 11839 9095
rect 17325 9061 17359 9095
rect 4077 8993 4111 9027
rect 11621 8993 11655 9027
rect 13461 8993 13495 9027
rect 13645 8993 13679 9027
rect 15209 8993 15243 9027
rect 15577 8993 15611 9027
rect 16129 8993 16163 9027
rect 16221 8993 16255 9027
rect 1869 8925 1903 8959
rect 1961 8925 1995 8959
rect 2145 8925 2179 8959
rect 2329 8925 2363 8959
rect 2697 8925 2731 8959
rect 2789 8925 2823 8959
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 3157 8925 3191 8959
rect 3617 8925 3651 8959
rect 4261 8925 4295 8959
rect 4353 8925 4387 8959
rect 4813 8925 4847 8959
rect 4997 8925 5031 8959
rect 5089 8925 5123 8959
rect 5273 8925 5307 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 6377 8925 6411 8959
rect 6653 8925 6687 8959
rect 6929 8925 6963 8959
rect 8585 8925 8619 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9781 8925 9815 8959
rect 9873 8925 9907 8959
rect 9965 8925 9999 8959
rect 10057 8925 10091 8959
rect 10241 8925 10275 8959
rect 10333 8925 10367 8959
rect 10517 8925 10551 8959
rect 10609 8925 10643 8959
rect 11253 8925 11287 8959
rect 11529 8925 11563 8959
rect 11897 8925 11931 8959
rect 13369 8925 13403 8959
rect 13553 8925 13587 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 14841 8925 14875 8959
rect 14933 8925 14967 8959
rect 15485 8925 15519 8959
rect 15669 8925 15703 8959
rect 15761 8925 15795 8959
rect 16313 8925 16347 8959
rect 16405 8925 16439 8959
rect 16589 8925 16623 8959
rect 16773 8925 16807 8959
rect 16957 8925 16991 8959
rect 17509 8925 17543 8959
rect 17601 8925 17635 8959
rect 6193 8857 6227 8891
rect 7205 8857 7239 8891
rect 7481 8857 7515 8891
rect 8217 8857 8251 8891
rect 15301 8857 15335 8891
rect 2421 8789 2455 8823
rect 3617 8789 3651 8823
rect 4997 8789 5031 8823
rect 5917 8789 5951 8823
rect 8401 8789 8435 8823
rect 10793 8789 10827 8823
rect 13185 8789 13219 8823
rect 15945 8789 15979 8823
rect 17785 8789 17819 8823
rect 8309 8585 8343 8619
rect 9505 8585 9539 8619
rect 10517 8585 10551 8619
rect 12541 8585 12575 8619
rect 14565 8585 14599 8619
rect 15577 8585 15611 8619
rect 17693 8585 17727 8619
rect 7021 8517 7055 8551
rect 7849 8517 7883 8551
rect 9045 8517 9079 8551
rect 12449 8517 12483 8551
rect 14933 8517 14967 8551
rect 16037 8517 16071 8551
rect 16865 8517 16899 8551
rect 16957 8517 16991 8551
rect 1685 8449 1719 8483
rect 2053 8449 2087 8483
rect 4261 8449 4295 8483
rect 4353 8449 4387 8483
rect 4630 8449 4664 8483
rect 4721 8449 4755 8483
rect 4997 8449 5031 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 6837 8449 6871 8483
rect 7941 8449 7975 8483
rect 8125 8449 8159 8483
rect 8217 8449 8251 8483
rect 8954 8471 8988 8505
rect 9137 8449 9171 8483
rect 9255 8449 9289 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 9965 8449 9999 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 11069 8449 11103 8483
rect 11161 8449 11195 8483
rect 11345 8449 11379 8483
rect 11805 8449 11839 8483
rect 11897 8449 11931 8483
rect 11989 8449 12023 8483
rect 12173 8449 12207 8483
rect 12817 8449 12851 8483
rect 13829 8449 13863 8483
rect 14013 8449 14047 8483
rect 14749 8449 14783 8483
rect 15025 8449 15059 8483
rect 15117 8449 15151 8483
rect 15577 8449 15611 8483
rect 15945 8449 15979 8483
rect 16129 8449 16163 8483
rect 16497 8449 16531 8483
rect 16773 8449 16807 8483
rect 17141 8449 17175 8483
rect 17233 8449 17267 8483
rect 17325 8449 17359 8483
rect 17417 8449 17451 8483
rect 17785 8449 17819 8483
rect 4077 8381 4111 8415
rect 9413 8381 9447 8415
rect 15393 8381 15427 8415
rect 16681 8381 16715 8415
rect 1501 8313 1535 8347
rect 1869 8313 1903 8347
rect 4169 8313 4203 8347
rect 4905 8313 4939 8347
rect 6377 8313 6411 8347
rect 8125 8313 8159 8347
rect 8769 8313 8803 8347
rect 10149 8313 10183 8347
rect 11345 8313 11379 8347
rect 12725 8313 12759 8347
rect 12909 8313 12943 8347
rect 13829 8313 13863 8347
rect 17969 8313 18003 8347
rect 4445 8245 4479 8279
rect 11529 8245 11563 8279
rect 15255 8245 15289 8279
rect 16313 8245 16347 8279
rect 17325 8245 17359 8279
rect 1501 8041 1535 8075
rect 5641 8041 5675 8075
rect 7113 8041 7147 8075
rect 9597 8041 9631 8075
rect 10149 8041 10183 8075
rect 11483 8041 11517 8075
rect 15577 8041 15611 8075
rect 17233 8041 17267 8075
rect 7205 7973 7239 8007
rect 8493 7973 8527 8007
rect 9321 7973 9355 8007
rect 14657 7973 14691 8007
rect 17417 7973 17451 8007
rect 1961 7905 1995 7939
rect 2145 7905 2179 7939
rect 5273 7905 5307 7939
rect 6101 7905 6135 7939
rect 8769 7905 8803 7939
rect 11621 7905 11655 7939
rect 11713 7905 11747 7939
rect 11897 7905 11931 7939
rect 12909 7905 12943 7939
rect 13277 7905 13311 7939
rect 13921 7905 13955 7939
rect 15025 7905 15059 7939
rect 15117 7905 15151 7939
rect 15301 7905 15335 7939
rect 15761 7905 15795 7939
rect 1869 7837 1903 7871
rect 4077 7837 4111 7871
rect 4261 7837 4295 7871
rect 4353 7837 4387 7871
rect 4445 7837 4479 7871
rect 5089 7837 5123 7871
rect 5181 7837 5215 7871
rect 5365 7837 5399 7871
rect 5549 7837 5583 7871
rect 5826 7837 5860 7871
rect 5918 7837 5952 7871
rect 6193 7837 6227 7871
rect 6469 7837 6503 7871
rect 6562 7837 6596 7871
rect 6745 7837 6779 7871
rect 6975 7837 7009 7871
rect 7205 7837 7239 7871
rect 7389 7837 7423 7871
rect 7487 7837 7521 7871
rect 7665 7837 7699 7871
rect 7849 7837 7883 7871
rect 8033 7837 8067 7871
rect 8125 7815 8159 7849
rect 8287 7837 8321 7871
rect 8401 7837 8435 7871
rect 8585 7837 8619 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 9229 7837 9263 7871
rect 9413 7837 9447 7871
rect 9965 7837 9999 7871
rect 10149 7837 10183 7871
rect 11345 7837 11379 7871
rect 11805 7837 11839 7871
rect 12081 7837 12115 7871
rect 12173 7837 12207 7871
rect 12265 7837 12299 7871
rect 12357 7837 12391 7871
rect 12541 7837 12575 7871
rect 12725 7837 12759 7871
rect 12817 7837 12851 7871
rect 13093 7837 13127 7871
rect 13461 7837 13495 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 14473 7837 14507 7871
rect 14841 7837 14875 7871
rect 14933 7837 14967 7871
rect 15577 7837 15611 7871
rect 17877 7837 17911 7871
rect 6837 7769 6871 7803
rect 13553 7769 13587 7803
rect 14289 7769 14323 7803
rect 14381 7769 14415 7803
rect 15853 7769 15887 7803
rect 16865 7769 16899 7803
rect 4721 7701 4755 7735
rect 4905 7701 4939 7735
rect 7573 7701 7607 7735
rect 8033 7701 8067 7735
rect 15393 7701 15427 7735
rect 17242 7701 17276 7735
rect 18061 7701 18095 7735
rect 1961 7497 1995 7531
rect 5273 7497 5307 7531
rect 13645 7497 13679 7531
rect 15025 7497 15059 7531
rect 15209 7497 15243 7531
rect 2421 7429 2455 7463
rect 3893 7429 3927 7463
rect 10403 7429 10437 7463
rect 1869 7361 1903 7395
rect 2605 7361 2639 7395
rect 2706 7361 2740 7395
rect 2973 7361 3007 7395
rect 3065 7361 3099 7395
rect 3157 7361 3191 7395
rect 3341 7361 3375 7395
rect 4077 7361 4111 7395
rect 4353 7361 4387 7395
rect 4537 7361 4571 7395
rect 4813 7361 4847 7395
rect 4905 7361 4939 7395
rect 5089 7361 5123 7395
rect 5181 7361 5215 7395
rect 5457 7361 5491 7395
rect 5641 7361 5675 7395
rect 5733 7361 5767 7395
rect 10701 7361 10735 7395
rect 13277 7361 13311 7395
rect 14381 7361 14415 7395
rect 14565 7361 14599 7395
rect 14841 7361 14875 7395
rect 15209 7361 15243 7395
rect 15393 7361 15427 7395
rect 2145 7293 2179 7327
rect 4261 7293 4295 7327
rect 10517 7293 10551 7327
rect 13369 7293 13403 7327
rect 2789 7225 2823 7259
rect 4169 7225 4203 7259
rect 10333 7225 10367 7259
rect 14657 7225 14691 7259
rect 14749 7225 14783 7259
rect 1501 7157 1535 7191
rect 2421 7157 2455 7191
rect 4629 7157 4663 7191
rect 10609 7157 10643 7191
rect 13277 7157 13311 7191
rect 4445 6953 4479 6987
rect 6653 6953 6687 6987
rect 9505 6953 9539 6987
rect 9965 6953 9999 6987
rect 10241 6953 10275 6987
rect 10701 6953 10735 6987
rect 10977 6953 11011 6987
rect 2605 6817 2639 6851
rect 4721 6817 4755 6851
rect 4905 6817 4939 6851
rect 5181 6817 5215 6851
rect 5365 6817 5399 6851
rect 9781 6817 9815 6851
rect 11345 6817 11379 6851
rect 15577 6817 15611 6851
rect 15669 6817 15703 6851
rect 1685 6749 1719 6783
rect 2513 6749 2547 6783
rect 2697 6749 2731 6783
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 4353 6749 4387 6783
rect 4629 6749 4663 6783
rect 4813 6749 4847 6783
rect 5089 6749 5123 6783
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 6837 6749 6871 6783
rect 7113 6749 7147 6783
rect 7481 6749 7515 6783
rect 7573 6749 7607 6783
rect 7941 6749 7975 6783
rect 10057 6749 10091 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 10428 6749 10462 6783
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 11161 6749 11195 6783
rect 11253 6749 11287 6783
rect 11437 6749 11471 6783
rect 11621 6749 11655 6783
rect 14928 6749 14962 6783
rect 15245 6749 15279 6783
rect 15393 6749 15427 6783
rect 15853 6749 15887 6783
rect 15945 6749 15979 6783
rect 16497 6749 16531 6783
rect 16865 6749 16899 6783
rect 17049 6749 17083 6783
rect 9689 6681 9723 6715
rect 15025 6681 15059 6715
rect 15117 6681 15151 6715
rect 1501 6613 1535 6647
rect 7021 6613 7055 6647
rect 9321 6613 9355 6647
rect 9489 6613 9523 6647
rect 9781 6613 9815 6647
rect 14749 6613 14783 6647
rect 15485 6613 15519 6647
rect 16681 6613 16715 6647
rect 17049 6613 17083 6647
rect 5917 6409 5951 6443
rect 6009 6409 6043 6443
rect 11719 6409 11753 6443
rect 15669 6409 15703 6443
rect 17233 6409 17267 6443
rect 1685 6341 1719 6375
rect 1869 6341 1903 6375
rect 3157 6341 3191 6375
rect 3877 6341 3911 6375
rect 4077 6341 4111 6375
rect 8539 6341 8573 6375
rect 8677 6341 8711 6375
rect 11621 6341 11655 6375
rect 16865 6341 16899 6375
rect 1961 6273 1995 6307
rect 2329 6273 2363 6307
rect 2421 6273 2455 6307
rect 2513 6273 2547 6307
rect 2697 6273 2731 6307
rect 2973 6273 3007 6307
rect 3249 6273 3283 6307
rect 5825 6273 5859 6307
rect 6193 6273 6227 6307
rect 6837 6273 6871 6307
rect 7481 6273 7515 6307
rect 8769 6273 8803 6307
rect 8861 6273 8895 6307
rect 9413 6273 9447 6307
rect 9505 6273 9539 6307
rect 9597 6273 9631 6307
rect 9781 6273 9815 6307
rect 11805 6273 11839 6307
rect 11897 6273 11931 6307
rect 12817 6273 12851 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 13093 6273 13127 6307
rect 13277 6273 13311 6307
rect 13553 6273 13587 6307
rect 16313 6273 16347 6307
rect 16497 6273 16531 6307
rect 16681 6273 16715 6307
rect 16957 6273 16991 6307
rect 17049 6273 17083 6307
rect 17325 6273 17359 6307
rect 17417 6273 17451 6307
rect 17601 6273 17635 6307
rect 17693 6273 17727 6307
rect 8401 6205 8435 6239
rect 13369 6205 13403 6239
rect 13645 6205 13679 6239
rect 13737 6205 13771 6239
rect 13829 6205 13863 6239
rect 15853 6205 15887 6239
rect 15945 6205 15979 6239
rect 16037 6205 16071 6239
rect 16129 6205 16163 6239
rect 16405 6205 16439 6239
rect 2789 6137 2823 6171
rect 3709 6137 3743 6171
rect 5917 6137 5951 6171
rect 7665 6137 7699 6171
rect 1685 6069 1719 6103
rect 2053 6069 2087 6103
rect 3893 6069 3927 6103
rect 9045 6069 9079 6103
rect 9137 6069 9171 6103
rect 17877 6069 17911 6103
rect 1961 5865 1995 5899
rect 2421 5865 2455 5899
rect 3065 5865 3099 5899
rect 8585 5865 8619 5899
rect 8677 5865 8711 5899
rect 8953 5865 8987 5899
rect 11069 5865 11103 5899
rect 13277 5865 13311 5899
rect 14105 5865 14139 5899
rect 14841 5865 14875 5899
rect 15853 5865 15887 5899
rect 17417 5865 17451 5899
rect 7113 5797 7147 5831
rect 13461 5797 13495 5831
rect 15393 5797 15427 5831
rect 3801 5729 3835 5763
rect 3985 5729 4019 5763
rect 4261 5729 4295 5763
rect 5641 5729 5675 5763
rect 8769 5729 8803 5763
rect 9413 5729 9447 5763
rect 12725 5729 12759 5763
rect 14473 5729 14507 5763
rect 14565 5729 14599 5763
rect 17233 5729 17267 5763
rect 1685 5661 1719 5695
rect 1777 5661 1811 5695
rect 1961 5661 1995 5695
rect 2605 5661 2639 5695
rect 2789 5661 2823 5695
rect 2881 5661 2915 5695
rect 3249 5661 3283 5695
rect 3341 5661 3375 5695
rect 3433 5661 3467 5695
rect 3525 5661 3559 5695
rect 4077 5661 4111 5695
rect 4169 5661 4203 5695
rect 5089 5661 5123 5695
rect 5181 5661 5215 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 6669 5671 6703 5705
rect 6929 5661 6963 5695
rect 8493 5661 8527 5695
rect 9137 5661 9171 5695
rect 9321 5661 9355 5695
rect 10609 5661 10643 5695
rect 10885 5661 10919 5695
rect 10977 5661 11011 5695
rect 12449 5661 12483 5695
rect 12541 5661 12575 5695
rect 12817 5661 12851 5695
rect 13093 5661 13127 5695
rect 13369 5661 13403 5695
rect 13461 5661 13495 5695
rect 13737 5661 13771 5695
rect 14289 5661 14323 5695
rect 14381 5661 14415 5695
rect 15025 5661 15059 5695
rect 15117 5661 15151 5695
rect 15761 5661 15795 5695
rect 15945 5661 15979 5695
rect 16589 5661 16623 5695
rect 17049 5661 17083 5695
rect 17141 5661 17175 5695
rect 5365 5593 5399 5627
rect 10793 5593 10827 5627
rect 12909 5593 12943 5627
rect 13645 5593 13679 5627
rect 15393 5593 15427 5627
rect 16221 5593 16255 5627
rect 6745 5525 6779 5559
rect 10425 5525 10459 5559
rect 12265 5525 12299 5559
rect 15209 5525 15243 5559
rect 6377 5321 6411 5355
rect 7849 5321 7883 5355
rect 9229 5321 9263 5355
rect 10425 5321 10459 5355
rect 12817 5321 12851 5355
rect 14105 5321 14139 5355
rect 14933 5321 14967 5355
rect 15577 5321 15611 5355
rect 12449 5253 12483 5287
rect 13737 5253 13771 5287
rect 17141 5253 17175 5287
rect 3341 5185 3375 5219
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 5641 5185 5675 5219
rect 6101 5185 6135 5219
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 6883 5185 6917 5219
rect 7205 5185 7239 5219
rect 7353 5185 7387 5219
rect 7481 5185 7515 5219
rect 7573 5185 7607 5219
rect 7670 5185 7704 5219
rect 8217 5185 8251 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 9045 5185 9079 5219
rect 9965 5185 9999 5219
rect 10241 5185 10275 5219
rect 10609 5185 10643 5219
rect 10885 5185 10919 5219
rect 11989 5185 12023 5219
rect 12357 5185 12391 5219
rect 12541 5185 12575 5219
rect 12817 5185 12851 5219
rect 13001 5185 13035 5219
rect 13645 5185 13679 5219
rect 13921 5185 13955 5219
rect 14197 5185 14231 5219
rect 14381 5185 14415 5219
rect 14473 5185 14507 5219
rect 14565 5185 14599 5219
rect 15117 5185 15151 5219
rect 15301 5185 15335 5219
rect 15761 5185 15795 5219
rect 16957 5185 16991 5219
rect 17325 5185 17359 5219
rect 3709 5117 3743 5151
rect 4261 5117 4295 5151
rect 4353 5117 4387 5151
rect 4537 5117 4571 5151
rect 5365 5117 5399 5151
rect 7021 5117 7055 5151
rect 11804 5117 11838 5151
rect 11897 5117 11931 5151
rect 12081 5117 12115 5151
rect 12265 5117 12299 5151
rect 15393 5117 15427 5151
rect 4813 5049 4847 5083
rect 10057 5049 10091 5083
rect 10149 5049 10183 5083
rect 10701 5049 10735 5083
rect 10793 5049 10827 5083
rect 14841 5049 14875 5083
rect 4997 4981 5031 5015
rect 8033 4981 8067 5015
rect 9781 4981 9815 5015
rect 3341 4777 3375 4811
rect 5917 4777 5951 4811
rect 7389 4777 7423 4811
rect 7849 4777 7883 4811
rect 8769 4777 8803 4811
rect 8953 4777 8987 4811
rect 10057 4777 10091 4811
rect 10701 4777 10735 4811
rect 11621 4777 11655 4811
rect 11805 4777 11839 4811
rect 14197 4777 14231 4811
rect 14657 4777 14691 4811
rect 15301 4777 15335 4811
rect 15853 4777 15887 4811
rect 7481 4709 7515 4743
rect 7941 4709 7975 4743
rect 11161 4709 11195 4743
rect 6194 4641 6228 4675
rect 6377 4641 6411 4675
rect 10149 4641 10183 4675
rect 11345 4641 11379 4675
rect 11897 4641 11931 4675
rect 12173 4641 12207 4675
rect 3433 4573 3467 4607
rect 4077 4573 4111 4607
rect 4813 4573 4847 4607
rect 4905 4573 4939 4607
rect 5457 4573 5491 4607
rect 6101 4573 6135 4607
rect 6285 4573 6319 4607
rect 6745 4573 6779 4607
rect 6929 4573 6963 4607
rect 7021 4573 7055 4607
rect 7113 4573 7147 4607
rect 7205 4573 7239 4607
rect 7757 4573 7791 4607
rect 8033 4573 8067 4607
rect 8217 4573 8251 4607
rect 8493 4573 8527 4607
rect 9137 4573 9171 4607
rect 9229 4573 9263 4607
rect 9873 4573 9907 4607
rect 10517 4573 10551 4607
rect 10793 4573 10827 4607
rect 11069 4573 11103 4607
rect 11253 4573 11287 4607
rect 11529 4573 11563 4607
rect 11989 4573 12023 4607
rect 12081 4573 12115 4607
rect 12265 4573 12299 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 14841 4573 14875 4607
rect 15209 4573 15243 4607
rect 15393 4573 15427 4607
rect 15577 4573 15611 4607
rect 16405 4573 16439 4607
rect 16589 4573 16623 4607
rect 16957 4573 16991 4607
rect 17325 4573 17359 4607
rect 3617 4505 3651 4539
rect 4353 4505 4387 4539
rect 8769 4505 8803 4539
rect 9597 4505 9631 4539
rect 15117 4505 15151 4539
rect 8585 4437 8619 4471
rect 9689 4437 9723 4471
rect 10241 4437 10275 4471
rect 10885 4437 10919 4471
rect 15025 4437 15059 4471
rect 16865 4437 16899 4471
rect 6193 4233 6227 4267
rect 10241 4233 10275 4267
rect 11529 4233 11563 4267
rect 12541 4233 12575 4267
rect 13369 4233 13403 4267
rect 6009 4165 6043 4199
rect 8309 4165 8343 4199
rect 3617 4097 3651 4131
rect 4537 4097 4571 4131
rect 5825 4097 5859 4131
rect 6469 4097 6503 4131
rect 6837 4097 6871 4131
rect 8953 4097 8987 4131
rect 9413 4097 9447 4131
rect 10149 4097 10183 4131
rect 10517 4097 10551 4131
rect 13001 4097 13035 4131
rect 13829 4097 13863 4131
rect 14381 4097 14415 4131
rect 14565 4097 14599 4131
rect 16313 4097 16347 4131
rect 16405 4097 16439 4131
rect 16681 4097 16715 4131
rect 16774 4097 16808 4131
rect 5457 4029 5491 4063
rect 9689 4029 9723 4063
rect 10333 4029 10367 4063
rect 11989 4029 12023 4063
rect 8493 3961 8527 3995
rect 8677 3961 8711 3995
rect 9597 3961 9631 3995
rect 11713 3961 11747 3995
rect 12725 3961 12759 3995
rect 13461 3961 13495 3995
rect 14565 3961 14599 3995
rect 9505 3893 9539 3927
rect 10517 3893 10551 3927
rect 16865 3893 16899 3927
rect 7297 3689 7331 3723
rect 7389 3621 7423 3655
rect 7757 3553 7791 3587
rect 9137 2397 9171 2431
rect 11989 2397 12023 2431
rect 9321 2261 9355 2295
rect 11805 2261 11839 2295
<< metal1 >>
rect 1104 19066 18492 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 18492 19066
rect 1104 18992 18492 19014
rect 7742 18912 7748 18964
rect 7800 18952 7806 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 7800 18924 8493 18952
rect 7800 18912 7806 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 8481 18915 8539 18921
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 10137 18955 10195 18961
rect 10137 18952 10149 18955
rect 9732 18924 10149 18952
rect 9732 18912 9738 18924
rect 10137 18921 10149 18924
rect 10183 18921 10195 18955
rect 10137 18915 10195 18921
rect 11606 18912 11612 18964
rect 11664 18952 11670 18964
rect 11885 18955 11943 18961
rect 11885 18952 11897 18955
rect 11664 18924 11897 18952
rect 11664 18912 11670 18924
rect 11885 18921 11897 18924
rect 11931 18921 11943 18955
rect 11885 18915 11943 18921
rect 8938 18844 8944 18896
rect 8996 18884 9002 18896
rect 12618 18884 12624 18896
rect 8996 18856 12624 18884
rect 8996 18844 9002 18856
rect 12618 18844 12624 18856
rect 12676 18844 12682 18896
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 10318 18816 10324 18828
rect 7984 18788 10324 18816
rect 7984 18776 7990 18788
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 8018 18708 8024 18760
rect 8076 18748 8082 18760
rect 8297 18751 8355 18757
rect 8297 18748 8309 18751
rect 8076 18720 8309 18748
rect 8076 18708 8082 18720
rect 8297 18717 8309 18720
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 9398 18708 9404 18760
rect 9456 18748 9462 18760
rect 9953 18751 10011 18757
rect 9953 18748 9965 18751
rect 9456 18720 9965 18748
rect 9456 18708 9462 18720
rect 9953 18717 9965 18720
rect 9999 18717 10011 18751
rect 9953 18711 10011 18717
rect 11698 18708 11704 18760
rect 11756 18708 11762 18760
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 13964 18720 14657 18748
rect 13964 18708 13970 18720
rect 14645 18717 14657 18720
rect 14691 18748 14703 18751
rect 16574 18748 16580 18760
rect 14691 18720 16580 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 16574 18708 16580 18720
rect 16632 18708 16638 18760
rect 7282 18640 7288 18692
rect 7340 18680 7346 18692
rect 7745 18683 7803 18689
rect 7745 18680 7757 18683
rect 7340 18652 7757 18680
rect 7340 18640 7346 18652
rect 7745 18649 7757 18652
rect 7791 18649 7803 18683
rect 7745 18643 7803 18649
rect 8113 18683 8171 18689
rect 8113 18649 8125 18683
rect 8159 18649 8171 18683
rect 8113 18643 8171 18649
rect 8128 18612 8156 18643
rect 9582 18640 9588 18692
rect 9640 18640 9646 18692
rect 9769 18683 9827 18689
rect 9769 18649 9781 18683
rect 9815 18680 9827 18683
rect 16666 18680 16672 18692
rect 9815 18652 16672 18680
rect 9815 18649 9827 18652
rect 9769 18643 9827 18649
rect 16666 18640 16672 18652
rect 16724 18640 16730 18692
rect 11882 18612 11888 18624
rect 8128 18584 11888 18612
rect 11882 18572 11888 18584
rect 11940 18572 11946 18624
rect 14737 18615 14795 18621
rect 14737 18581 14749 18615
rect 14783 18612 14795 18615
rect 15378 18612 15384 18624
rect 14783 18584 15384 18612
rect 14783 18581 14795 18584
rect 14737 18575 14795 18581
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 1104 18522 18492 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 18492 18522
rect 1104 18448 18492 18470
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 2004 18380 7420 18408
rect 2004 18368 2010 18380
rect 2332 18312 7328 18340
rect 2332 18284 2360 18312
rect 7300 18284 7328 18312
rect 2314 18232 2320 18284
rect 2372 18232 2378 18284
rect 3789 18275 3847 18281
rect 3789 18241 3801 18275
rect 3835 18241 3847 18275
rect 3789 18235 3847 18241
rect 2222 18028 2228 18080
rect 2280 18028 2286 18080
rect 3602 18028 3608 18080
rect 3660 18028 3666 18080
rect 3804 18068 3832 18235
rect 7098 18232 7104 18284
rect 7156 18232 7162 18284
rect 7282 18232 7288 18284
rect 7340 18232 7346 18284
rect 7392 18272 7420 18380
rect 7834 18368 7840 18420
rect 7892 18368 7898 18420
rect 8018 18368 8024 18420
rect 8076 18368 8082 18420
rect 9398 18368 9404 18420
rect 9456 18368 9462 18420
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 13265 18411 13323 18417
rect 13265 18408 13277 18411
rect 10376 18380 10916 18408
rect 10376 18368 10382 18380
rect 7855 18312 9536 18340
rect 7855 18281 7883 18312
rect 7840 18275 7898 18281
rect 7840 18272 7852 18275
rect 7392 18244 7852 18272
rect 7840 18241 7852 18244
rect 7886 18241 7898 18275
rect 7840 18235 7898 18241
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 8076 18244 8493 18272
rect 8076 18232 8082 18244
rect 8481 18241 8493 18244
rect 8527 18272 8539 18275
rect 8757 18275 8815 18281
rect 8757 18272 8769 18275
rect 8527 18244 8769 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 8757 18241 8769 18244
rect 8803 18241 8815 18275
rect 8757 18235 8815 18241
rect 8938 18232 8944 18284
rect 8996 18232 9002 18284
rect 9508 18272 9536 18312
rect 9575 18275 9633 18281
rect 9575 18272 9587 18275
rect 9508 18244 9587 18272
rect 9575 18241 9587 18244
rect 9621 18241 9633 18275
rect 9575 18235 9633 18241
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18272 9919 18275
rect 9907 18244 10088 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 7193 18207 7251 18213
rect 7193 18173 7205 18207
rect 7239 18204 7251 18207
rect 7377 18207 7435 18213
rect 7377 18204 7389 18207
rect 7239 18176 7389 18204
rect 7239 18173 7251 18176
rect 7193 18167 7251 18173
rect 7377 18173 7389 18176
rect 7423 18173 7435 18207
rect 7377 18167 7435 18173
rect 8294 18164 8300 18216
rect 8352 18164 8358 18216
rect 8386 18164 8392 18216
rect 8444 18164 8450 18216
rect 8570 18164 8576 18216
rect 8628 18164 8634 18216
rect 7469 18139 7527 18145
rect 7469 18105 7481 18139
rect 7515 18136 7527 18139
rect 8113 18139 8171 18145
rect 8113 18136 8125 18139
rect 7515 18108 8125 18136
rect 7515 18105 7527 18108
rect 7469 18099 7527 18105
rect 8113 18105 8125 18108
rect 8159 18105 8171 18139
rect 8113 18099 8171 18105
rect 8956 18068 8984 18232
rect 9600 18204 9628 18235
rect 10060 18213 10088 18244
rect 10134 18232 10140 18284
rect 10192 18272 10198 18284
rect 10888 18281 10916 18380
rect 12406 18380 13277 18408
rect 11882 18300 11888 18352
rect 11940 18340 11946 18352
rect 12406 18340 12434 18380
rect 13265 18377 13277 18380
rect 13311 18377 13323 18411
rect 13265 18371 13323 18377
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 13412 18380 16436 18408
rect 13412 18368 13418 18380
rect 11940 18312 12434 18340
rect 11940 18300 11946 18312
rect 13722 18300 13728 18352
rect 13780 18300 13786 18352
rect 16408 18284 16436 18380
rect 10413 18275 10471 18281
rect 10413 18272 10425 18275
rect 10192 18244 10425 18272
rect 10192 18232 10198 18244
rect 10413 18241 10425 18244
rect 10459 18272 10471 18275
rect 10689 18275 10747 18281
rect 10689 18272 10701 18275
rect 10459 18244 10701 18272
rect 10459 18241 10471 18244
rect 10413 18235 10471 18241
rect 10689 18241 10701 18244
rect 10735 18241 10747 18275
rect 10689 18235 10747 18241
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12986 18272 12992 18284
rect 12529 18235 12587 18241
rect 12636 18244 12992 18272
rect 10045 18207 10103 18213
rect 9600 18176 9904 18204
rect 9677 18139 9735 18145
rect 9677 18105 9689 18139
rect 9723 18105 9735 18139
rect 9677 18099 9735 18105
rect 3804 18040 8984 18068
rect 9692 18068 9720 18099
rect 9766 18096 9772 18148
rect 9824 18096 9830 18148
rect 9876 18136 9904 18176
rect 10045 18173 10057 18207
rect 10091 18173 10103 18207
rect 10045 18167 10103 18173
rect 10226 18164 10232 18216
rect 10284 18164 10290 18216
rect 10318 18164 10324 18216
rect 10376 18164 10382 18216
rect 10505 18207 10563 18213
rect 10505 18173 10517 18207
rect 10551 18204 10563 18207
rect 11974 18204 11980 18216
rect 10551 18176 11980 18204
rect 10551 18173 10563 18176
rect 10505 18167 10563 18173
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 12544 18136 12572 18235
rect 12636 18213 12664 18244
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 13170 18232 13176 18284
rect 13228 18232 13234 18284
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18272 15347 18275
rect 15470 18272 15476 18284
rect 15335 18244 15476 18272
rect 15335 18241 15347 18244
rect 15289 18235 15347 18241
rect 15470 18232 15476 18244
rect 15528 18272 15534 18284
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15528 18244 15761 18272
rect 15528 18232 15534 18244
rect 15749 18241 15761 18244
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18272 15991 18275
rect 16022 18272 16028 18284
rect 15979 18244 16028 18272
rect 15979 18241 15991 18244
rect 15933 18235 15991 18241
rect 16022 18232 16028 18244
rect 16080 18272 16086 18284
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 16080 18244 16313 18272
rect 16080 18232 16086 18244
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 16301 18235 16359 18241
rect 16390 18232 16396 18284
rect 16448 18232 16454 18284
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16632 18244 16681 18272
rect 16632 18232 16638 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18173 12679 18207
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 12621 18167 12679 18173
rect 12912 18176 14749 18204
rect 12912 18145 12940 18176
rect 14737 18173 14749 18176
rect 14783 18173 14795 18207
rect 14737 18167 14795 18173
rect 15010 18164 15016 18216
rect 15068 18164 15074 18216
rect 15102 18164 15108 18216
rect 15160 18204 15166 18216
rect 15197 18207 15255 18213
rect 15197 18204 15209 18207
rect 15160 18176 15209 18204
rect 15160 18164 15166 18176
rect 15197 18173 15209 18176
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 9876 18108 12572 18136
rect 12897 18139 12955 18145
rect 12897 18105 12909 18139
rect 12943 18105 12955 18139
rect 12897 18099 12955 18105
rect 13173 18139 13231 18145
rect 13173 18105 13185 18139
rect 13219 18136 13231 18139
rect 15657 18139 15715 18145
rect 13219 18108 13768 18136
rect 13219 18105 13231 18108
rect 13173 18099 13231 18105
rect 10781 18071 10839 18077
rect 10781 18068 10793 18071
rect 9692 18040 10793 18068
rect 10781 18037 10793 18040
rect 10827 18037 10839 18071
rect 10781 18031 10839 18037
rect 11974 18028 11980 18080
rect 12032 18028 12038 18080
rect 13740 18068 13768 18108
rect 15657 18105 15669 18139
rect 15703 18136 15715 18139
rect 16206 18136 16212 18148
rect 15703 18108 16212 18136
rect 15703 18105 15715 18108
rect 15657 18099 15715 18105
rect 16206 18096 16212 18108
rect 16264 18096 16270 18148
rect 14366 18068 14372 18080
rect 13740 18040 14372 18068
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 16758 18028 16764 18080
rect 16816 18028 16822 18080
rect 1104 17978 18492 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 18492 17978
rect 1104 17904 18492 17926
rect 7098 17824 7104 17876
rect 7156 17824 7162 17876
rect 7653 17867 7711 17873
rect 7653 17833 7665 17867
rect 7699 17864 7711 17867
rect 7834 17864 7840 17876
rect 7699 17836 7840 17864
rect 7699 17833 7711 17836
rect 7653 17827 7711 17833
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 9030 17864 9036 17876
rect 7944 17836 9036 17864
rect 2406 17756 2412 17808
rect 2464 17796 2470 17808
rect 2464 17768 6684 17796
rect 2464 17756 2470 17768
rect 3602 17728 3608 17740
rect 3436 17700 3608 17728
rect 1670 17620 1676 17672
rect 1728 17620 1734 17672
rect 2590 17552 2596 17604
rect 2648 17592 2654 17604
rect 3436 17601 3464 17700
rect 3602 17688 3608 17700
rect 3660 17728 3666 17740
rect 6656 17728 6684 17768
rect 6730 17756 6736 17808
rect 6788 17796 6794 17808
rect 7944 17796 7972 17836
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 10045 17867 10103 17873
rect 10045 17864 10057 17867
rect 9824 17836 10057 17864
rect 9824 17824 9830 17836
rect 10045 17833 10057 17836
rect 10091 17833 10103 17867
rect 10045 17827 10103 17833
rect 10226 17824 10232 17876
rect 10284 17864 10290 17876
rect 10781 17867 10839 17873
rect 10781 17864 10793 17867
rect 10284 17836 10793 17864
rect 10284 17824 10290 17836
rect 10781 17833 10793 17836
rect 10827 17833 10839 17867
rect 10781 17827 10839 17833
rect 11333 17867 11391 17873
rect 11333 17833 11345 17867
rect 11379 17864 11391 17867
rect 11698 17864 11704 17876
rect 11379 17836 11704 17864
rect 11379 17833 11391 17836
rect 11333 17827 11391 17833
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 12805 17867 12863 17873
rect 12805 17833 12817 17867
rect 12851 17833 12863 17867
rect 12805 17827 12863 17833
rect 8294 17796 8300 17808
rect 6788 17768 7972 17796
rect 8036 17768 8300 17796
rect 6788 17756 6794 17768
rect 8036 17728 8064 17768
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 8389 17799 8447 17805
rect 8389 17765 8401 17799
rect 8435 17765 8447 17799
rect 12345 17799 12403 17805
rect 12345 17796 12357 17799
rect 8389 17759 8447 17765
rect 11992 17768 12357 17796
rect 8404 17728 8432 17759
rect 10689 17731 10747 17737
rect 10689 17728 10701 17731
rect 3660 17700 4108 17728
rect 6656 17700 7328 17728
rect 3660 17688 3666 17700
rect 3878 17620 3884 17672
rect 3936 17620 3942 17672
rect 4080 17669 4108 17700
rect 7300 17672 7328 17700
rect 7852 17700 8064 17728
rect 8220 17700 8432 17728
rect 10244 17700 10701 17728
rect 4065 17663 4123 17669
rect 4065 17629 4077 17663
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 5166 17620 5172 17672
rect 5224 17620 5230 17672
rect 7282 17620 7288 17672
rect 7340 17620 7346 17672
rect 7558 17620 7564 17672
rect 7616 17620 7622 17672
rect 7852 17669 7880 17700
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17660 7987 17663
rect 8110 17660 8116 17672
rect 7975 17632 8116 17660
rect 7975 17629 7987 17632
rect 7929 17623 7987 17629
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 8220 17669 8248 17700
rect 10244 17672 10272 17700
rect 10689 17697 10701 17700
rect 10735 17697 10747 17731
rect 10689 17691 10747 17697
rect 10778 17688 10784 17740
rect 10836 17728 10842 17740
rect 11992 17737 12020 17768
rect 12345 17765 12357 17768
rect 12391 17765 12403 17799
rect 12820 17796 12848 17827
rect 12986 17824 12992 17876
rect 13044 17824 13050 17876
rect 13081 17867 13139 17873
rect 13081 17833 13093 17867
rect 13127 17864 13139 17867
rect 13170 17864 13176 17876
rect 13127 17836 13176 17864
rect 13127 17833 13139 17836
rect 13081 17827 13139 17833
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 13722 17824 13728 17876
rect 13780 17864 13786 17876
rect 13817 17867 13875 17873
rect 13817 17864 13829 17867
rect 13780 17836 13829 17864
rect 13780 17824 13786 17836
rect 13817 17833 13829 17836
rect 13863 17833 13875 17867
rect 14458 17864 14464 17876
rect 13817 17827 13875 17833
rect 13924 17836 14464 17864
rect 13262 17796 13268 17808
rect 12820 17768 13268 17796
rect 12345 17759 12403 17765
rect 13262 17756 13268 17768
rect 13320 17756 13326 17808
rect 11149 17731 11207 17737
rect 10836 17700 11100 17728
rect 10836 17688 10842 17700
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 8297 17663 8355 17669
rect 8297 17629 8309 17663
rect 8343 17660 8355 17663
rect 8478 17660 8484 17672
rect 8343 17632 8484 17660
rect 8343 17629 8355 17632
rect 8297 17623 8355 17629
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8662 17620 8668 17672
rect 8720 17620 8726 17672
rect 9214 17620 9220 17672
rect 9272 17620 9278 17672
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17660 9551 17663
rect 9950 17660 9956 17672
rect 9539 17632 9956 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 9950 17620 9956 17632
rect 10008 17620 10014 17672
rect 10226 17620 10232 17672
rect 10284 17620 10290 17672
rect 10410 17620 10416 17672
rect 10468 17620 10474 17672
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17660 10563 17663
rect 10594 17660 10600 17672
rect 10551 17632 10600 17660
rect 10551 17629 10563 17632
rect 10505 17623 10563 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 10870 17620 10876 17672
rect 10928 17620 10934 17672
rect 10962 17620 10968 17672
rect 11020 17620 11026 17672
rect 11072 17669 11100 17700
rect 11149 17697 11161 17731
rect 11195 17728 11207 17731
rect 11977 17731 12035 17737
rect 11195 17700 11652 17728
rect 11195 17697 11207 17700
rect 11149 17691 11207 17697
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11238 17620 11244 17672
rect 11296 17620 11302 17672
rect 11514 17620 11520 17672
rect 11572 17620 11578 17672
rect 11624 17660 11652 17700
rect 11977 17697 11989 17731
rect 12023 17697 12035 17731
rect 13924 17728 13952 17836
rect 14458 17824 14464 17836
rect 14516 17864 14522 17876
rect 15102 17864 15108 17876
rect 14516 17836 15108 17864
rect 14516 17824 14522 17836
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 11977 17691 12035 17697
rect 13372 17700 13952 17728
rect 12069 17663 12127 17669
rect 12069 17660 12081 17663
rect 11624 17632 12081 17660
rect 12069 17629 12081 17632
rect 12115 17629 12127 17663
rect 12069 17623 12127 17629
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 12710 17660 12716 17672
rect 12391 17632 12716 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 3421 17595 3479 17601
rect 3421 17592 3433 17595
rect 2648 17564 3433 17592
rect 2648 17552 2654 17564
rect 3421 17561 3433 17564
rect 3467 17561 3479 17595
rect 3421 17555 3479 17561
rect 3605 17595 3663 17601
rect 3605 17561 3617 17595
rect 3651 17592 3663 17595
rect 3786 17592 3792 17604
rect 3651 17564 3792 17592
rect 3651 17561 3663 17564
rect 3605 17555 3663 17561
rect 3786 17552 3792 17564
rect 3844 17552 3850 17604
rect 7190 17552 7196 17604
rect 7248 17592 7254 17604
rect 7742 17592 7748 17604
rect 7248 17564 7748 17592
rect 7248 17552 7254 17564
rect 7742 17552 7748 17564
rect 7800 17592 7806 17604
rect 8018 17592 8024 17604
rect 7800 17564 8024 17592
rect 7800 17552 7806 17564
rect 8018 17552 8024 17564
rect 8076 17552 8082 17604
rect 8389 17595 8447 17601
rect 8389 17561 8401 17595
rect 8435 17592 8447 17595
rect 8435 17564 8708 17592
rect 8435 17561 8447 17564
rect 8389 17555 8447 17561
rect 1486 17484 1492 17536
rect 1544 17484 1550 17536
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 3694 17524 3700 17536
rect 3292 17496 3700 17524
rect 3292 17484 3298 17496
rect 3694 17484 3700 17496
rect 3752 17484 3758 17536
rect 4062 17484 4068 17536
rect 4120 17484 4126 17536
rect 4798 17484 4804 17536
rect 4856 17524 4862 17536
rect 4985 17527 5043 17533
rect 4985 17524 4997 17527
rect 4856 17496 4997 17524
rect 4856 17484 4862 17496
rect 4985 17493 4997 17496
rect 5031 17493 5043 17527
rect 4985 17487 5043 17493
rect 7469 17527 7527 17533
rect 7469 17493 7481 17527
rect 7515 17524 7527 17527
rect 7650 17524 7656 17536
rect 7515 17496 7656 17524
rect 7515 17493 7527 17496
rect 7469 17487 7527 17493
rect 7650 17484 7656 17496
rect 7708 17524 7714 17536
rect 8573 17527 8631 17533
rect 8573 17524 8585 17527
rect 7708 17496 8585 17524
rect 7708 17484 7714 17496
rect 8573 17493 8585 17496
rect 8619 17493 8631 17527
rect 8680 17524 8708 17564
rect 8754 17552 8760 17604
rect 8812 17592 8818 17604
rect 9677 17595 9735 17601
rect 8812 17564 9444 17592
rect 8812 17552 8818 17564
rect 8846 17524 8852 17536
rect 8680 17496 8852 17524
rect 8573 17487 8631 17493
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 9306 17484 9312 17536
rect 9364 17484 9370 17536
rect 9416 17524 9444 17564
rect 9677 17561 9689 17595
rect 9723 17592 9735 17595
rect 11609 17595 11667 17601
rect 11609 17592 11621 17595
rect 9723 17564 11621 17592
rect 9723 17561 9735 17564
rect 9677 17555 9735 17561
rect 11609 17561 11621 17564
rect 11655 17561 11667 17595
rect 11609 17555 11667 17561
rect 11698 17552 11704 17604
rect 11756 17552 11762 17604
rect 11819 17595 11877 17601
rect 11819 17561 11831 17595
rect 11865 17561 11877 17595
rect 11819 17555 11877 17561
rect 10502 17524 10508 17536
rect 9416 17496 10508 17524
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 10594 17484 10600 17536
rect 10652 17524 10658 17536
rect 10962 17524 10968 17536
rect 10652 17496 10968 17524
rect 10652 17484 10658 17496
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 11834 17524 11862 17555
rect 11974 17552 11980 17604
rect 12032 17592 12038 17604
rect 12360 17592 12388 17623
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 13372 17669 13400 17700
rect 14366 17688 14372 17740
rect 14424 17688 14430 17740
rect 15010 17688 15016 17740
rect 15068 17728 15074 17740
rect 15933 17731 15991 17737
rect 15933 17728 15945 17731
rect 15068 17700 15945 17728
rect 15068 17688 15074 17700
rect 15933 17697 15945 17700
rect 15979 17697 15991 17731
rect 15933 17691 15991 17697
rect 16206 17688 16212 17740
rect 16264 17688 16270 17740
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 12852 17635 13369 17660
rect 12851 17632 13369 17635
rect 12851 17629 12909 17632
rect 12032 17564 12388 17592
rect 12032 17552 12038 17564
rect 12618 17552 12624 17604
rect 12676 17552 12682 17604
rect 12851 17595 12863 17629
rect 12897 17595 12909 17629
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 13357 17623 13415 17629
rect 13906 17620 13912 17672
rect 13964 17620 13970 17672
rect 14090 17620 14096 17672
rect 14148 17620 14154 17672
rect 12851 17589 12909 17595
rect 13081 17595 13139 17601
rect 13081 17561 13093 17595
rect 13127 17592 13139 17595
rect 14642 17592 14648 17604
rect 13127 17564 14648 17592
rect 13127 17561 13139 17564
rect 13081 17555 13139 17561
rect 11388 17496 11862 17524
rect 12161 17527 12219 17533
rect 11388 17484 11394 17496
rect 12161 17493 12173 17527
rect 12207 17524 12219 17527
rect 12250 17524 12256 17536
rect 12207 17496 12256 17524
rect 12207 17493 12219 17496
rect 12161 17487 12219 17493
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12636 17524 12664 17552
rect 13096 17524 13124 17555
rect 14642 17552 14648 17564
rect 14700 17552 14706 17604
rect 15378 17552 15384 17604
rect 15436 17552 15442 17604
rect 16758 17552 16764 17604
rect 16816 17552 16822 17604
rect 12636 17496 13124 17524
rect 13262 17484 13268 17536
rect 13320 17484 13326 17536
rect 15841 17527 15899 17533
rect 15841 17493 15853 17527
rect 15887 17524 15899 17527
rect 15930 17524 15936 17536
rect 15887 17496 15936 17524
rect 15887 17493 15899 17496
rect 15841 17487 15899 17493
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 17678 17484 17684 17536
rect 17736 17484 17742 17536
rect 1104 17434 18492 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 18492 17434
rect 1104 17360 18492 17382
rect 5810 17280 5816 17332
rect 5868 17320 5874 17332
rect 5868 17292 7236 17320
rect 5868 17280 5874 17292
rect 2593 17255 2651 17261
rect 2593 17221 2605 17255
rect 2639 17252 2651 17255
rect 3234 17252 3240 17264
rect 2639 17224 3240 17252
rect 2639 17221 2651 17224
rect 2593 17215 2651 17221
rect 3234 17212 3240 17224
rect 3292 17212 3298 17264
rect 3436 17224 4660 17252
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17184 1915 17187
rect 1946 17184 1952 17196
rect 1903 17156 1952 17184
rect 1903 17153 1915 17156
rect 1857 17147 1915 17153
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 3326 17144 3332 17196
rect 3384 17144 3390 17196
rect 3436 17193 3464 17224
rect 4632 17196 4660 17224
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 3513 17187 3571 17193
rect 3513 17153 3525 17187
rect 3559 17153 3571 17187
rect 3513 17147 3571 17153
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17184 3755 17187
rect 3786 17184 3792 17196
rect 3743 17156 3792 17184
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 2148 17048 2176 17079
rect 2682 17076 2688 17128
rect 2740 17116 2746 17128
rect 3528 17116 3556 17147
rect 2740 17088 3556 17116
rect 3712 17116 3740 17147
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 4614 17144 4620 17196
rect 4672 17144 4678 17196
rect 4798 17144 4804 17196
rect 4856 17144 4862 17196
rect 5718 17144 5724 17196
rect 5776 17144 5782 17196
rect 6270 17144 6276 17196
rect 6328 17184 6334 17196
rect 6917 17187 6975 17193
rect 6917 17184 6929 17187
rect 6328 17156 6929 17184
rect 6328 17144 6334 17156
rect 6917 17153 6929 17156
rect 6963 17153 6975 17187
rect 6917 17147 6975 17153
rect 7098 17144 7104 17196
rect 7156 17144 7162 17196
rect 7208 17193 7236 17292
rect 7650 17280 7656 17332
rect 7708 17280 7714 17332
rect 8294 17280 8300 17332
rect 8352 17280 8358 17332
rect 9214 17320 9220 17332
rect 8496 17292 9220 17320
rect 7837 17255 7895 17261
rect 7837 17221 7849 17255
rect 7883 17252 7895 17255
rect 8496 17252 8524 17292
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 9677 17323 9735 17329
rect 9677 17320 9689 17323
rect 9364 17292 9689 17320
rect 9364 17280 9370 17292
rect 9677 17289 9689 17292
rect 9723 17289 9735 17323
rect 9677 17283 9735 17289
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 9824 17292 10456 17320
rect 9824 17280 9830 17292
rect 7883 17224 8524 17252
rect 8573 17255 8631 17261
rect 7883 17221 7895 17224
rect 7837 17215 7895 17221
rect 8573 17221 8585 17255
rect 8619 17252 8631 17255
rect 8619 17224 9352 17252
rect 8619 17221 8631 17224
rect 8573 17215 8631 17221
rect 9324 17196 9352 17224
rect 9416 17224 10272 17252
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 7745 17187 7803 17193
rect 7745 17184 7757 17187
rect 7432 17156 7757 17184
rect 7432 17144 7438 17156
rect 7745 17153 7757 17156
rect 7791 17153 7803 17187
rect 7745 17147 7803 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 8481 17187 8539 17193
rect 8481 17153 8493 17187
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17153 8723 17187
rect 8665 17147 8723 17153
rect 6730 17116 6736 17128
rect 3712 17088 6736 17116
rect 2740 17076 2746 17088
rect 2406 17048 2412 17060
rect 2148 17020 2412 17048
rect 2406 17008 2412 17020
rect 2464 17008 2470 17060
rect 3528 17048 3556 17088
rect 6730 17076 6736 17088
rect 6788 17076 6794 17128
rect 7466 17076 7472 17128
rect 7524 17076 7530 17128
rect 7558 17076 7564 17128
rect 7616 17076 7622 17128
rect 7944 17116 7972 17147
rect 7668 17088 7972 17116
rect 8496 17116 8524 17147
rect 8570 17116 8576 17128
rect 8496 17088 8576 17116
rect 7190 17048 7196 17060
rect 3528 17020 7196 17048
rect 7190 17008 7196 17020
rect 7248 17008 7254 17060
rect 7484 17048 7512 17076
rect 7668 17048 7696 17088
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 8680 17116 8708 17147
rect 8846 17144 8852 17196
rect 8904 17144 8910 17196
rect 8938 17144 8944 17196
rect 8996 17144 9002 17196
rect 9030 17144 9036 17196
rect 9088 17144 9094 17196
rect 9214 17193 9220 17196
rect 9181 17187 9220 17193
rect 9181 17153 9193 17187
rect 9181 17147 9220 17153
rect 9214 17144 9220 17147
rect 9272 17144 9278 17196
rect 9306 17144 9312 17196
rect 9364 17144 9370 17196
rect 9416 17193 9444 17224
rect 10244 17196 10272 17224
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17153 9459 17187
rect 9401 17147 9459 17153
rect 9539 17187 9597 17193
rect 9539 17153 9551 17187
rect 9585 17184 9597 17187
rect 9766 17184 9772 17196
rect 9585 17156 9772 17184
rect 9585 17153 9597 17156
rect 9539 17147 9597 17153
rect 9416 17116 9444 17147
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 9876 17156 10149 17184
rect 8680 17088 9444 17116
rect 8680 17048 8708 17088
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 9876 17116 9904 17156
rect 10137 17153 10149 17156
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 10226 17144 10232 17196
rect 10284 17144 10290 17196
rect 10428 17193 10456 17292
rect 12250 17280 12256 17332
rect 12308 17280 12314 17332
rect 14090 17280 14096 17332
rect 14148 17320 14154 17332
rect 15010 17320 15016 17332
rect 14148 17292 15016 17320
rect 14148 17280 14154 17292
rect 13262 17252 13268 17264
rect 11716 17224 13268 17252
rect 11716 17196 11744 17224
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 14752 17261 14780 17292
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 16390 17280 16396 17332
rect 16448 17320 16454 17332
rect 17773 17323 17831 17329
rect 17773 17320 17785 17323
rect 16448 17292 17785 17320
rect 16448 17280 16454 17292
rect 17773 17289 17785 17292
rect 17819 17289 17831 17323
rect 17773 17283 17831 17289
rect 14737 17255 14795 17261
rect 14737 17221 14749 17255
rect 14783 17221 14795 17255
rect 14737 17215 14795 17221
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17153 10471 17187
rect 10413 17147 10471 17153
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 11793 17187 11851 17193
rect 11793 17153 11805 17187
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 9732 17088 9904 17116
rect 9953 17119 10011 17125
rect 9732 17076 9738 17088
rect 9953 17085 9965 17119
rect 9999 17085 10011 17119
rect 9953 17079 10011 17085
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 10318 17116 10324 17128
rect 10091 17088 10324 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 7484 17020 7696 17048
rect 8404 17020 8708 17048
rect 8404 16992 8432 17020
rect 9122 17008 9128 17060
rect 9180 17048 9186 17060
rect 9769 17051 9827 17057
rect 9769 17048 9781 17051
rect 9180 17020 9781 17048
rect 9180 17008 9186 17020
rect 9769 17017 9781 17020
rect 9815 17017 9827 17051
rect 9769 17011 9827 17017
rect 1673 16983 1731 16989
rect 1673 16949 1685 16983
rect 1719 16980 1731 16983
rect 1854 16980 1860 16992
rect 1719 16952 1860 16980
rect 1719 16949 1731 16952
rect 1673 16943 1731 16949
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 2038 16940 2044 16992
rect 2096 16940 2102 16992
rect 3050 16940 3056 16992
rect 3108 16940 3114 16992
rect 4985 16983 5043 16989
rect 4985 16949 4997 16983
rect 5031 16980 5043 16983
rect 5074 16980 5080 16992
rect 5031 16952 5080 16980
rect 5031 16949 5043 16952
rect 4985 16943 5043 16949
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 5442 16940 5448 16992
rect 5500 16980 5506 16992
rect 5629 16983 5687 16989
rect 5629 16980 5641 16983
rect 5500 16952 5641 16980
rect 5500 16940 5506 16952
rect 5629 16949 5641 16952
rect 5675 16980 5687 16983
rect 6178 16980 6184 16992
rect 5675 16952 6184 16980
rect 5675 16949 5687 16952
rect 5629 16943 5687 16949
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6917 16983 6975 16989
rect 6917 16949 6929 16983
rect 6963 16980 6975 16983
rect 7006 16980 7012 16992
rect 6963 16952 7012 16980
rect 6963 16949 6975 16952
rect 6917 16943 6975 16949
rect 7006 16940 7012 16952
rect 7064 16940 7070 16992
rect 7282 16940 7288 16992
rect 7340 16940 7346 16992
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 8386 16980 8392 16992
rect 7616 16952 8392 16980
rect 7616 16940 7622 16952
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9582 16940 9588 16992
rect 9640 16980 9646 16992
rect 9674 16980 9680 16992
rect 9640 16952 9680 16980
rect 9640 16940 9646 16952
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 9968 16980 9996 17079
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 11808 17116 11836 17147
rect 11974 17144 11980 17196
rect 12032 17144 12038 17196
rect 12066 17144 12072 17196
rect 12124 17144 12130 17196
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17184 14151 17187
rect 14182 17184 14188 17196
rect 14139 17156 14188 17184
rect 14139 17153 14151 17156
rect 14093 17147 14151 17153
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 14550 17144 14556 17196
rect 14608 17184 14614 17196
rect 14608 17156 16344 17184
rect 14608 17144 14614 17156
rect 16316 17128 16344 17156
rect 16482 17144 16488 17196
rect 16540 17144 16546 17196
rect 16666 17144 16672 17196
rect 16724 17144 16730 17196
rect 17678 17144 17684 17196
rect 17736 17144 17742 17196
rect 12802 17116 12808 17128
rect 11808 17088 12808 17116
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 16298 17076 16304 17128
rect 16356 17116 16362 17128
rect 16945 17119 17003 17125
rect 16945 17116 16957 17119
rect 16356 17088 16957 17116
rect 16356 17076 16362 17088
rect 16945 17085 16957 17088
rect 16991 17085 17003 17119
rect 16945 17079 17003 17085
rect 11606 17008 11612 17060
rect 11664 17048 11670 17060
rect 11974 17048 11980 17060
rect 11664 17020 11980 17048
rect 11664 17008 11670 17020
rect 11974 17008 11980 17020
rect 12032 17048 12038 17060
rect 12032 17020 14504 17048
rect 12032 17008 12038 17020
rect 9916 16952 9996 16980
rect 9916 16940 9922 16952
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10597 16983 10655 16989
rect 10597 16980 10609 16983
rect 10284 16952 10609 16980
rect 10284 16940 10290 16952
rect 10597 16949 10609 16952
rect 10643 16980 10655 16983
rect 10686 16980 10692 16992
rect 10643 16952 10692 16980
rect 10643 16949 10655 16952
rect 10597 16943 10655 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 14476 16989 14504 17020
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13596 16952 13921 16980
rect 13596 16940 13602 16952
rect 13909 16949 13921 16952
rect 13955 16949 13967 16983
rect 13909 16943 13967 16949
rect 14461 16983 14519 16989
rect 14461 16949 14473 16983
rect 14507 16980 14519 16983
rect 14918 16980 14924 16992
rect 14507 16952 14924 16980
rect 14507 16949 14519 16952
rect 14461 16943 14519 16949
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 1104 16890 18492 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 18492 16890
rect 1104 16816 18492 16838
rect 1489 16779 1547 16785
rect 1489 16745 1501 16779
rect 1535 16776 1547 16779
rect 1670 16776 1676 16788
rect 1535 16748 1676 16776
rect 1535 16745 1547 16748
rect 1489 16739 1547 16745
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 3418 16776 3424 16788
rect 2792 16748 3424 16776
rect 2792 16717 2820 16748
rect 3418 16736 3424 16748
rect 3476 16736 3482 16788
rect 3510 16736 3516 16788
rect 3568 16776 3574 16788
rect 3878 16776 3884 16788
rect 3568 16748 3884 16776
rect 3568 16736 3574 16748
rect 3878 16736 3884 16748
rect 3936 16736 3942 16788
rect 4433 16779 4491 16785
rect 4433 16745 4445 16779
rect 4479 16776 4491 16779
rect 5718 16776 5724 16788
rect 4479 16748 5724 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 7098 16776 7104 16788
rect 5828 16748 7104 16776
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16677 2835 16711
rect 2777 16671 2835 16677
rect 2869 16711 2927 16717
rect 2869 16677 2881 16711
rect 2915 16708 2927 16711
rect 3142 16708 3148 16720
rect 2915 16680 3148 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 3326 16668 3332 16720
rect 3384 16708 3390 16720
rect 3602 16708 3608 16720
rect 3384 16680 3608 16708
rect 3384 16668 3390 16680
rect 3602 16668 3608 16680
rect 3660 16708 3666 16720
rect 4798 16708 4804 16720
rect 3660 16680 4804 16708
rect 3660 16668 3666 16680
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 2498 16640 2504 16652
rect 2179 16612 2504 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3160 16612 3801 16640
rect 1854 16532 1860 16584
rect 1912 16532 1918 16584
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 2314 16572 2320 16584
rect 1995 16544 2320 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 2314 16532 2320 16544
rect 2372 16532 2378 16584
rect 2682 16532 2688 16584
rect 2740 16532 2746 16584
rect 3160 16581 3188 16612
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 4290 16640 4318 16680
rect 4798 16668 4804 16680
rect 4856 16668 4862 16720
rect 5828 16708 5856 16748
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 7374 16736 7380 16788
rect 7432 16736 7438 16788
rect 9122 16736 9128 16788
rect 9180 16776 9186 16788
rect 9217 16779 9275 16785
rect 9217 16776 9229 16779
rect 9180 16748 9229 16776
rect 9180 16736 9186 16748
rect 9217 16745 9229 16748
rect 9263 16745 9275 16779
rect 9217 16739 9275 16745
rect 9306 16736 9312 16788
rect 9364 16776 9370 16788
rect 9585 16779 9643 16785
rect 9585 16776 9597 16779
rect 9364 16748 9597 16776
rect 9364 16736 9370 16748
rect 9585 16745 9597 16748
rect 9631 16745 9643 16779
rect 9585 16739 9643 16745
rect 10410 16736 10416 16788
rect 10468 16736 10474 16788
rect 10502 16736 10508 16788
rect 10560 16776 10566 16788
rect 11609 16779 11667 16785
rect 11609 16776 11621 16779
rect 10560 16748 11621 16776
rect 10560 16736 10566 16748
rect 11609 16745 11621 16748
rect 11655 16745 11667 16779
rect 11609 16739 11667 16745
rect 11977 16779 12035 16785
rect 11977 16745 11989 16779
rect 12023 16776 12035 16779
rect 12066 16776 12072 16788
rect 12023 16748 12072 16776
rect 12023 16745 12035 16748
rect 11977 16739 12035 16745
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 12802 16736 12808 16788
rect 12860 16736 12866 16788
rect 14829 16779 14887 16785
rect 14829 16745 14841 16779
rect 14875 16776 14887 16779
rect 15730 16779 15788 16785
rect 15730 16776 15742 16779
rect 14875 16748 15742 16776
rect 14875 16745 14887 16748
rect 14829 16739 14887 16745
rect 15730 16745 15742 16748
rect 15776 16745 15788 16779
rect 15730 16739 15788 16745
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 17221 16779 17279 16785
rect 17221 16776 17233 16779
rect 16816 16748 17233 16776
rect 16816 16736 16822 16748
rect 17221 16745 17233 16748
rect 17267 16745 17279 16779
rect 17221 16739 17279 16745
rect 4908 16680 5856 16708
rect 4290 16612 4384 16640
rect 3789 16603 3847 16609
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16541 3019 16575
rect 2961 16535 3019 16541
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16541 3203 16575
rect 3145 16535 3203 16541
rect 2976 16504 3004 16535
rect 3234 16532 3240 16584
rect 3292 16572 3298 16584
rect 3510 16572 3516 16584
rect 3292 16544 3516 16572
rect 3292 16532 3298 16544
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 3602 16532 3608 16584
rect 3660 16532 3666 16584
rect 3694 16532 3700 16584
rect 3752 16572 3758 16584
rect 4356 16581 4384 16612
rect 3973 16575 4031 16581
rect 3973 16572 3985 16575
rect 3752 16544 3985 16572
rect 3752 16532 3758 16544
rect 3973 16541 3985 16544
rect 4019 16541 4031 16575
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 3973 16535 4031 16541
rect 4080 16544 4261 16572
rect 2976 16476 3648 16504
rect 2130 16396 2136 16448
rect 2188 16436 2194 16448
rect 2501 16439 2559 16445
rect 2501 16436 2513 16439
rect 2188 16408 2513 16436
rect 2188 16396 2194 16408
rect 2501 16405 2513 16408
rect 2547 16405 2559 16439
rect 3620 16436 3648 16476
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 4080 16504 4108 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4341 16575 4399 16581
rect 4341 16541 4353 16575
rect 4387 16541 4399 16575
rect 4341 16535 4399 16541
rect 4796 16575 4854 16581
rect 4796 16541 4808 16575
rect 4842 16572 4854 16575
rect 4908 16572 4936 16680
rect 7006 16668 7012 16720
rect 7064 16668 7070 16720
rect 8938 16668 8944 16720
rect 8996 16708 9002 16720
rect 12342 16708 12348 16720
rect 8996 16680 12348 16708
rect 8996 16668 9002 16680
rect 12342 16668 12348 16680
rect 12400 16668 12406 16720
rect 14737 16711 14795 16717
rect 14737 16677 14749 16711
rect 14783 16708 14795 16711
rect 14921 16711 14979 16717
rect 14921 16708 14933 16711
rect 14783 16680 14933 16708
rect 14783 16677 14795 16680
rect 14737 16671 14795 16677
rect 14921 16677 14933 16680
rect 14967 16677 14979 16711
rect 14921 16671 14979 16677
rect 6273 16643 6331 16649
rect 6273 16640 6285 16643
rect 4842 16544 4936 16572
rect 5000 16612 6285 16640
rect 4842 16541 4854 16544
rect 4796 16535 4854 16541
rect 3936 16476 4108 16504
rect 3936 16464 3942 16476
rect 4154 16464 4160 16516
rect 4212 16504 4218 16516
rect 4212 16476 4844 16504
rect 4212 16464 4218 16476
rect 4617 16439 4675 16445
rect 4617 16436 4629 16439
rect 3620 16408 4629 16436
rect 2501 16399 2559 16405
rect 4617 16405 4629 16408
rect 4663 16405 4675 16439
rect 4816 16436 4844 16476
rect 4890 16464 4896 16516
rect 4948 16464 4954 16516
rect 5000 16513 5028 16612
rect 6273 16609 6285 16612
rect 6319 16609 6331 16643
rect 6273 16603 6331 16609
rect 6656 16612 7696 16640
rect 5074 16532 5080 16584
rect 5132 16581 5138 16584
rect 5132 16575 5171 16581
rect 5159 16541 5171 16575
rect 5132 16535 5171 16541
rect 5261 16575 5319 16581
rect 5261 16541 5273 16575
rect 5307 16572 5319 16575
rect 5626 16572 5632 16584
rect 5307 16544 5632 16572
rect 5307 16541 5319 16544
rect 5261 16535 5319 16541
rect 5132 16532 5138 16535
rect 5626 16532 5632 16544
rect 5684 16532 5690 16584
rect 5905 16575 5963 16581
rect 5905 16541 5917 16575
rect 5951 16541 5963 16575
rect 5905 16535 5963 16541
rect 4985 16507 5043 16513
rect 4985 16473 4997 16507
rect 5031 16473 5043 16507
rect 5920 16504 5948 16535
rect 6178 16532 6184 16584
rect 6236 16532 6242 16584
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 6656 16581 6684 16612
rect 6641 16575 6699 16581
rect 6641 16572 6653 16575
rect 6420 16544 6653 16572
rect 6420 16532 6426 16544
rect 6641 16541 6653 16544
rect 6687 16541 6699 16575
rect 6641 16535 6699 16541
rect 6730 16532 6736 16584
rect 6788 16532 6794 16584
rect 6917 16575 6975 16581
rect 6917 16541 6929 16575
rect 6963 16541 6975 16575
rect 6917 16535 6975 16541
rect 6454 16504 6460 16516
rect 5920 16476 6460 16504
rect 4985 16467 5043 16473
rect 5000 16436 5028 16467
rect 6454 16464 6460 16476
rect 6512 16464 6518 16516
rect 4816 16408 5028 16436
rect 6932 16436 6960 16535
rect 7006 16532 7012 16584
rect 7064 16572 7070 16584
rect 7101 16575 7159 16581
rect 7101 16572 7113 16575
rect 7064 16544 7113 16572
rect 7064 16532 7070 16544
rect 7101 16541 7113 16544
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16572 7251 16575
rect 7558 16572 7564 16584
rect 7239 16544 7564 16572
rect 7239 16541 7251 16544
rect 7193 16535 7251 16541
rect 7116 16504 7144 16535
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 7668 16572 7696 16612
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 8628 16612 10180 16640
rect 8628 16600 8634 16612
rect 7668 16544 8984 16572
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 7116 16476 7481 16504
rect 7469 16473 7481 16476
rect 7515 16473 7527 16507
rect 7469 16467 7527 16473
rect 7834 16464 7840 16516
rect 7892 16504 7898 16516
rect 8021 16507 8079 16513
rect 8021 16504 8033 16507
rect 7892 16476 8033 16504
rect 7892 16464 7898 16476
rect 8021 16473 8033 16476
rect 8067 16473 8079 16507
rect 8021 16467 8079 16473
rect 8205 16507 8263 16513
rect 8205 16473 8217 16507
rect 8251 16504 8263 16507
rect 8846 16504 8852 16516
rect 8251 16476 8852 16504
rect 8251 16473 8263 16476
rect 8205 16467 8263 16473
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 8956 16504 8984 16544
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 9309 16575 9367 16581
rect 9309 16572 9321 16575
rect 9272 16544 9321 16572
rect 9272 16532 9278 16544
rect 9309 16541 9321 16544
rect 9355 16541 9367 16575
rect 9309 16535 9367 16541
rect 9490 16532 9496 16584
rect 9548 16532 9554 16584
rect 9674 16532 9680 16584
rect 9732 16532 9738 16584
rect 10152 16581 10180 16612
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 11296 16612 11744 16640
rect 11296 16600 11302 16612
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16541 10103 16575
rect 10045 16535 10103 16541
rect 10137 16575 10195 16581
rect 10137 16541 10149 16575
rect 10183 16541 10195 16575
rect 10137 16535 10195 16541
rect 9692 16504 9720 16532
rect 8956 16476 9720 16504
rect 9766 16464 9772 16516
rect 9824 16464 9830 16516
rect 10060 16504 10088 16535
rect 10226 16532 10232 16584
rect 10284 16532 10290 16584
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16572 10471 16575
rect 10686 16572 10692 16584
rect 10459 16544 10692 16572
rect 10459 16541 10471 16544
rect 10413 16535 10471 16541
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16541 11575 16575
rect 11716 16572 11744 16612
rect 11790 16600 11796 16652
rect 11848 16600 11854 16652
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 11974 16640 11980 16652
rect 11931 16612 11980 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 12492 16612 13492 16640
rect 12492 16600 12498 16612
rect 12069 16575 12127 16581
rect 12069 16572 12081 16575
rect 11716 16544 12081 16572
rect 11517 16535 11575 16541
rect 12069 16541 12081 16544
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12250 16572 12256 16584
rect 12207 16544 12256 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 10244 16504 10272 16532
rect 10060 16476 10272 16504
rect 11532 16504 11560 16535
rect 12176 16504 12204 16535
rect 12250 16532 12256 16544
rect 12308 16532 12314 16584
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 11532 16476 12204 16504
rect 13096 16504 13124 16535
rect 13170 16532 13176 16584
rect 13228 16532 13234 16584
rect 13262 16532 13268 16584
rect 13320 16532 13326 16584
rect 13464 16581 13492 16612
rect 13906 16600 13912 16652
rect 13964 16640 13970 16652
rect 14369 16643 14427 16649
rect 14369 16640 14381 16643
rect 13964 16612 14381 16640
rect 13964 16600 13970 16612
rect 14369 16609 14381 16612
rect 14415 16640 14427 16643
rect 14458 16640 14464 16652
rect 14415 16612 14464 16640
rect 14415 16609 14427 16612
rect 14369 16603 14427 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16640 15531 16643
rect 15838 16640 15844 16652
rect 15519 16612 15844 16640
rect 15519 16609 15531 16612
rect 15473 16603 15531 16609
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 16816 16612 17540 16640
rect 16816 16600 16822 16612
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16541 13507 16575
rect 13449 16535 13507 16541
rect 14918 16532 14924 16584
rect 14976 16572 14982 16584
rect 15105 16575 15163 16581
rect 15105 16572 15117 16575
rect 14976 16544 15117 16572
rect 14976 16532 14982 16544
rect 15105 16541 15117 16544
rect 15151 16541 15163 16575
rect 15105 16535 15163 16541
rect 15378 16532 15384 16584
rect 15436 16532 15442 16584
rect 17512 16581 17540 16612
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16541 17555 16575
rect 17497 16535 17555 16541
rect 14182 16504 14188 16516
rect 13096 16476 14188 16504
rect 14182 16464 14188 16476
rect 14240 16464 14246 16516
rect 17405 16507 17463 16513
rect 17405 16504 17417 16507
rect 16974 16476 17417 16504
rect 17405 16473 17417 16476
rect 17451 16473 17463 16507
rect 17405 16467 17463 16473
rect 7190 16436 7196 16448
rect 6932 16408 7196 16436
rect 4617 16399 4675 16405
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 9858 16436 9864 16448
rect 9916 16445 9922 16448
rect 9825 16408 9864 16436
rect 9858 16396 9864 16408
rect 9916 16399 9925 16445
rect 9953 16439 10011 16445
rect 9953 16405 9965 16439
rect 9999 16436 10011 16439
rect 10042 16436 10048 16448
rect 9999 16408 10048 16436
rect 9999 16405 10011 16408
rect 9953 16399 10011 16405
rect 9916 16396 9922 16399
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 10229 16439 10287 16445
rect 10229 16405 10241 16439
rect 10275 16436 10287 16439
rect 10318 16436 10324 16448
rect 10275 16408 10324 16436
rect 10275 16405 10287 16408
rect 10229 16399 10287 16405
rect 10318 16396 10324 16408
rect 10376 16436 10382 16448
rect 10502 16436 10508 16448
rect 10376 16408 10508 16436
rect 10376 16396 10382 16408
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 11698 16396 11704 16448
rect 11756 16436 11762 16448
rect 11793 16439 11851 16445
rect 11793 16436 11805 16439
rect 11756 16408 11805 16436
rect 11756 16396 11762 16408
rect 11793 16405 11805 16408
rect 11839 16405 11851 16439
rect 11793 16399 11851 16405
rect 13998 16396 14004 16448
rect 14056 16436 14062 16448
rect 14550 16436 14556 16448
rect 14056 16408 14556 16436
rect 14056 16396 14062 16408
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 15286 16396 15292 16448
rect 15344 16396 15350 16448
rect 1104 16346 18492 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 18492 16346
rect 1104 16272 18492 16294
rect 1854 16192 1860 16244
rect 1912 16232 1918 16244
rect 1949 16235 2007 16241
rect 1949 16232 1961 16235
rect 1912 16204 1961 16232
rect 1912 16192 1918 16204
rect 1949 16201 1961 16204
rect 1995 16201 2007 16235
rect 1949 16195 2007 16201
rect 2498 16192 2504 16244
rect 2556 16192 2562 16244
rect 4154 16232 4160 16244
rect 2700 16204 4160 16232
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 1857 16099 1915 16105
rect 1857 16096 1869 16099
rect 1820 16068 1869 16096
rect 1820 16056 1826 16068
rect 1857 16065 1869 16068
rect 1903 16096 1915 16099
rect 2314 16096 2320 16108
rect 1903 16068 2320 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 2700 16105 2728 16204
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 4264 16204 8892 16232
rect 2866 16124 2872 16176
rect 2924 16164 2930 16176
rect 3418 16164 3424 16176
rect 2924 16136 3424 16164
rect 2924 16124 2930 16136
rect 3418 16124 3424 16136
rect 3476 16164 3482 16176
rect 4264 16164 4292 16204
rect 5350 16164 5356 16176
rect 3476 16136 4292 16164
rect 4356 16136 5356 16164
rect 3476 16124 3482 16136
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16065 2743 16099
rect 2685 16059 2743 16065
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16096 3019 16099
rect 3050 16096 3056 16108
rect 3007 16068 3056 16096
rect 3007 16065 3019 16068
rect 2961 16059 3019 16065
rect 3050 16056 3056 16068
rect 3108 16056 3114 16108
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4157 16059 4215 16065
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 4356 16096 4384 16136
rect 4295 16068 4384 16096
rect 4433 16099 4491 16105
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 4433 16065 4445 16099
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 4525 16099 4583 16105
rect 4525 16065 4537 16099
rect 4571 16096 4583 16099
rect 4798 16096 4804 16108
rect 4571 16068 4804 16096
rect 4571 16065 4583 16068
rect 4525 16059 4583 16065
rect 2130 15988 2136 16040
rect 2188 15988 2194 16040
rect 2777 16031 2835 16037
rect 2777 16028 2789 16031
rect 2240 16000 2789 16028
rect 1854 15920 1860 15972
rect 1912 15960 1918 15972
rect 2038 15960 2044 15972
rect 1912 15932 2044 15960
rect 1912 15920 1918 15932
rect 2038 15920 2044 15932
rect 2096 15960 2102 15972
rect 2240 15960 2268 16000
rect 2777 15997 2789 16000
rect 2823 15997 2835 16031
rect 2777 15991 2835 15997
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 16028 2927 16031
rect 4062 16028 4068 16040
rect 2915 16000 4068 16028
rect 2915 15997 2927 16000
rect 2869 15991 2927 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 2096 15932 2268 15960
rect 2096 15920 2102 15932
rect 3694 15920 3700 15972
rect 3752 15960 3758 15972
rect 4172 15960 4200 16059
rect 4448 16028 4476 16059
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 5074 16056 5080 16108
rect 5132 16096 5138 16108
rect 5184 16105 5212 16136
rect 5350 16124 5356 16136
rect 5408 16124 5414 16176
rect 7193 16167 7251 16173
rect 5920 16136 7052 16164
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 5132 16068 5181 16096
rect 5132 16056 5138 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5169 16059 5227 16065
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 5534 16096 5540 16108
rect 5316 16068 5540 16096
rect 5316 16056 5322 16068
rect 5534 16056 5540 16068
rect 5592 16096 5598 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5592 16068 5733 16096
rect 5592 16056 5598 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 5721 16059 5779 16065
rect 5810 16056 5816 16108
rect 5868 16096 5874 16108
rect 5920 16105 5948 16136
rect 5905 16099 5963 16105
rect 5905 16096 5917 16099
rect 5868 16068 5917 16096
rect 5868 16056 5874 16068
rect 5905 16065 5917 16068
rect 5951 16065 5963 16099
rect 5905 16059 5963 16065
rect 6178 16056 6184 16108
rect 6236 16096 6242 16108
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 6236 16068 6377 16096
rect 6236 16056 6242 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 6914 16056 6920 16108
rect 6972 16056 6978 16108
rect 7024 16105 7052 16136
rect 7193 16133 7205 16167
rect 7239 16164 7251 16167
rect 8754 16164 8760 16176
rect 7239 16136 8760 16164
rect 7239 16133 7251 16136
rect 7193 16127 7251 16133
rect 7009 16099 7067 16105
rect 7009 16065 7021 16099
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 6270 16028 6276 16040
rect 4448 16000 6276 16028
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 7208 16028 7236 16127
rect 8754 16124 8760 16136
rect 8812 16124 8818 16176
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16065 7435 16099
rect 8864 16096 8892 16204
rect 9784 16204 10732 16232
rect 9306 16124 9312 16176
rect 9364 16164 9370 16176
rect 9784 16164 9812 16204
rect 9364 16136 9812 16164
rect 9364 16124 9370 16136
rect 9125 16099 9183 16105
rect 9125 16096 9137 16099
rect 8864 16068 9137 16096
rect 7377 16059 7435 16065
rect 9125 16065 9137 16068
rect 9171 16065 9183 16099
rect 9125 16059 9183 16065
rect 6380 16000 7236 16028
rect 3752 15932 4200 15960
rect 3752 15920 3758 15932
rect 1489 15895 1547 15901
rect 1489 15861 1501 15895
rect 1535 15892 1547 15895
rect 1670 15892 1676 15904
rect 1535 15864 1676 15892
rect 1535 15861 1547 15864
rect 1489 15855 1547 15861
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 3142 15852 3148 15904
rect 3200 15892 3206 15904
rect 3973 15895 4031 15901
rect 3973 15892 3985 15895
rect 3200 15864 3985 15892
rect 3200 15852 3206 15864
rect 3973 15861 3985 15864
rect 4019 15861 4031 15895
rect 4172 15892 4200 15932
rect 5718 15920 5724 15972
rect 5776 15920 5782 15972
rect 5994 15920 6000 15972
rect 6052 15960 6058 15972
rect 6380 15960 6408 16000
rect 6052 15932 6408 15960
rect 6052 15920 6058 15932
rect 6822 15920 6828 15972
rect 6880 15920 6886 15972
rect 7006 15920 7012 15972
rect 7064 15960 7070 15972
rect 7392 15960 7420 16059
rect 9490 16056 9496 16108
rect 9548 16056 9554 16108
rect 9784 16105 9812 16136
rect 10318 16124 10324 16176
rect 10376 16164 10382 16176
rect 10376 16136 10645 16164
rect 10376 16124 10382 16136
rect 9769 16099 9827 16105
rect 9769 16065 9781 16099
rect 9815 16065 9827 16099
rect 9769 16059 9827 16065
rect 9950 16056 9956 16108
rect 10008 16096 10014 16108
rect 10617 16105 10645 16136
rect 10137 16099 10195 16105
rect 10137 16096 10149 16099
rect 10008 16068 10149 16096
rect 10008 16056 10014 16068
rect 10137 16065 10149 16068
rect 10183 16065 10195 16099
rect 10137 16059 10195 16065
rect 10230 16099 10288 16105
rect 10230 16065 10242 16099
rect 10276 16065 10288 16099
rect 10230 16059 10288 16065
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 10505 16099 10563 16105
rect 10505 16065 10517 16099
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 10602 16099 10660 16105
rect 10602 16065 10614 16099
rect 10648 16065 10660 16099
rect 10704 16096 10732 16204
rect 10778 16192 10784 16244
rect 10836 16192 10842 16244
rect 11330 16192 11336 16244
rect 11388 16192 11394 16244
rect 11514 16192 11520 16244
rect 11572 16192 11578 16244
rect 13081 16235 13139 16241
rect 11900 16204 12204 16232
rect 10870 16124 10876 16176
rect 10928 16124 10934 16176
rect 11422 16124 11428 16176
rect 11480 16164 11486 16176
rect 11900 16164 11928 16204
rect 11480 16136 11928 16164
rect 11480 16124 11486 16136
rect 11146 16096 11152 16108
rect 10704 16068 11152 16096
rect 10602 16059 10660 16065
rect 10042 15988 10048 16040
rect 10100 16028 10106 16040
rect 10244 16028 10272 16059
rect 10100 16000 10272 16028
rect 10100 15988 10106 16000
rect 10428 15972 10456 16059
rect 10520 16028 10548 16059
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 11330 16056 11336 16108
rect 11388 16096 11394 16108
rect 11900 16105 11928 16136
rect 12066 16124 12072 16176
rect 12124 16124 12130 16176
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 11388 16068 11805 16096
rect 11388 16056 11394 16068
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12084 16096 12112 16124
rect 12023 16068 12112 16096
rect 12176 16096 12204 16204
rect 13081 16201 13093 16235
rect 13127 16232 13139 16235
rect 13262 16232 13268 16244
rect 13127 16204 13268 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13262 16192 13268 16204
rect 13320 16192 13326 16244
rect 13906 16192 13912 16244
rect 13964 16232 13970 16244
rect 14093 16235 14151 16241
rect 14093 16232 14105 16235
rect 13964 16204 14105 16232
rect 13964 16192 13970 16204
rect 14093 16201 14105 16204
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 14550 16192 14556 16244
rect 14608 16232 14614 16244
rect 14608 16204 16804 16232
rect 14608 16192 14614 16204
rect 16776 16176 16804 16204
rect 12342 16124 12348 16176
rect 12400 16164 12406 16176
rect 13633 16167 13691 16173
rect 13633 16164 13645 16167
rect 12400 16136 13645 16164
rect 12400 16124 12406 16136
rect 13280 16105 13308 16136
rect 13633 16133 13645 16136
rect 13679 16133 13691 16167
rect 13633 16127 13691 16133
rect 13817 16167 13875 16173
rect 13817 16133 13829 16167
rect 13863 16164 13875 16167
rect 13998 16164 14004 16176
rect 13863 16136 14004 16164
rect 13863 16133 13875 16136
rect 13817 16127 13875 16133
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 14231 16133 14289 16139
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 12176 16068 12449 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 10778 16028 10784 16040
rect 10520 16000 10784 16028
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 11020 16000 11069 16028
rect 11020 15988 11026 16000
rect 11057 15997 11069 16000
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 12066 15988 12072 16040
rect 12124 16028 12130 16040
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 12124 16000 12173 16028
rect 12124 15988 12130 16000
rect 12161 15997 12173 16000
rect 12207 15997 12219 16031
rect 12452 16028 12480 16059
rect 13446 16056 13452 16108
rect 13504 16056 13510 16108
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14231 16099 14243 16133
rect 14277 16130 14289 16133
rect 14277 16099 14304 16130
rect 14458 16124 14464 16176
rect 14516 16124 14522 16176
rect 15378 16164 15384 16176
rect 14568 16136 15384 16164
rect 14231 16096 14304 16099
rect 14568 16096 14596 16136
rect 15378 16124 15384 16136
rect 15436 16164 15442 16176
rect 15436 16136 16160 16164
rect 15436 16124 15442 16136
rect 13964 16068 14596 16096
rect 13964 16056 13970 16068
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 14700 16068 15669 16096
rect 14700 16056 14706 16068
rect 15657 16065 15669 16068
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 15930 16056 15936 16108
rect 15988 16056 15994 16108
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16065 16083 16099
rect 16132 16096 16160 16136
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 16853 16167 16911 16173
rect 16853 16164 16865 16167
rect 16816 16136 16865 16164
rect 16816 16124 16822 16136
rect 16853 16133 16865 16136
rect 16899 16133 16911 16167
rect 17681 16167 17739 16173
rect 17681 16164 17693 16167
rect 16853 16127 16911 16133
rect 16960 16136 17693 16164
rect 16960 16096 16988 16136
rect 17681 16133 17693 16136
rect 17727 16133 17739 16167
rect 17681 16127 17739 16133
rect 16132 16068 16988 16096
rect 17497 16099 17555 16105
rect 16025 16059 16083 16065
rect 17497 16065 17509 16099
rect 17543 16065 17555 16099
rect 17497 16059 17555 16065
rect 15470 16028 15476 16040
rect 12452 16000 15476 16028
rect 12161 15991 12219 15997
rect 15470 15988 15476 16000
rect 15528 15988 15534 16040
rect 16040 16028 16068 16059
rect 15948 16000 16068 16028
rect 15948 15972 15976 16000
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 17313 16031 17371 16037
rect 17313 16028 17325 16031
rect 17000 16000 17325 16028
rect 17000 15988 17006 16000
rect 17313 15997 17325 16000
rect 17359 15997 17371 16031
rect 17313 15991 17371 15997
rect 7064 15932 7420 15960
rect 7561 15963 7619 15969
rect 7064 15920 7070 15932
rect 7561 15929 7573 15963
rect 7607 15960 7619 15963
rect 10410 15960 10416 15972
rect 7607 15932 10416 15960
rect 7607 15929 7619 15932
rect 7561 15923 7619 15929
rect 10410 15920 10416 15932
rect 10468 15920 10474 15972
rect 12621 15963 12679 15969
rect 12621 15960 12633 15963
rect 11782 15932 12633 15960
rect 5258 15892 5264 15904
rect 4172 15864 5264 15892
rect 3973 15855 4031 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 6086 15852 6092 15904
rect 6144 15892 6150 15904
rect 6454 15892 6460 15904
rect 6144 15864 6460 15892
rect 6144 15852 6150 15864
rect 6454 15852 6460 15864
rect 6512 15892 6518 15904
rect 8018 15892 8024 15904
rect 6512 15864 8024 15892
rect 6512 15852 6518 15864
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 9309 15895 9367 15901
rect 9309 15861 9321 15895
rect 9355 15892 9367 15895
rect 9766 15892 9772 15904
rect 9355 15864 9772 15892
rect 9355 15861 9367 15864
rect 9309 15855 9367 15861
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 9858 15852 9864 15904
rect 9916 15852 9922 15904
rect 10045 15895 10103 15901
rect 10045 15861 10057 15895
rect 10091 15892 10103 15895
rect 10686 15892 10692 15904
rect 10091 15864 10692 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 11782 15892 11810 15932
rect 12621 15929 12633 15932
rect 12667 15929 12679 15963
rect 12621 15923 12679 15929
rect 13538 15920 13544 15972
rect 13596 15960 13602 15972
rect 15286 15960 15292 15972
rect 13596 15932 15292 15960
rect 13596 15920 13602 15932
rect 11195 15864 11810 15892
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 12253 15895 12311 15901
rect 12253 15892 12265 15895
rect 12216 15864 12265 15892
rect 12216 15852 12222 15864
rect 12253 15861 12265 15864
rect 12299 15861 12311 15895
rect 12253 15855 12311 15861
rect 13998 15852 14004 15904
rect 14056 15852 14062 15904
rect 14292 15901 14320 15932
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 15930 15920 15936 15972
rect 15988 15920 15994 15972
rect 17221 15963 17279 15969
rect 17221 15960 17233 15963
rect 16224 15932 17233 15960
rect 14277 15895 14335 15901
rect 14277 15861 14289 15895
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 15194 15892 15200 15904
rect 14967 15864 15200 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 16224 15901 16252 15932
rect 17221 15929 17233 15932
rect 17267 15929 17279 15963
rect 17221 15923 17279 15929
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 15620 15864 16221 15892
rect 15620 15852 15626 15864
rect 16209 15861 16221 15864
rect 16255 15861 16267 15895
rect 16209 15855 16267 15861
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17512 15892 17540 16059
rect 16908 15864 17540 15892
rect 16908 15852 16914 15864
rect 1104 15802 18492 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 18492 15802
rect 1104 15728 18492 15750
rect 1302 15648 1308 15700
rect 1360 15688 1366 15700
rect 1489 15691 1547 15697
rect 1489 15688 1501 15691
rect 1360 15660 1501 15688
rect 1360 15648 1366 15660
rect 1489 15657 1501 15660
rect 1535 15657 1547 15691
rect 1489 15651 1547 15657
rect 3513 15691 3571 15697
rect 3513 15657 3525 15691
rect 3559 15688 3571 15691
rect 3878 15688 3884 15700
rect 3559 15660 3884 15688
rect 3559 15657 3571 15660
rect 3513 15651 3571 15657
rect 3878 15648 3884 15660
rect 3936 15648 3942 15700
rect 4249 15691 4307 15697
rect 4249 15657 4261 15691
rect 4295 15688 4307 15691
rect 4706 15688 4712 15700
rect 4295 15660 4712 15688
rect 4295 15657 4307 15660
rect 4249 15651 4307 15657
rect 2958 15580 2964 15632
rect 3016 15620 3022 15632
rect 4264 15620 4292 15651
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 5166 15648 5172 15700
rect 5224 15688 5230 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 5224 15660 5457 15688
rect 5224 15648 5230 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 5445 15651 5503 15657
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 5684 15660 6776 15688
rect 5684 15648 5690 15660
rect 6086 15620 6092 15632
rect 3016 15592 4292 15620
rect 4356 15592 6092 15620
rect 3016 15580 3022 15592
rect 3234 15552 3240 15564
rect 2976 15524 3240 15552
rect 1670 15444 1676 15496
rect 1728 15444 1734 15496
rect 2222 15444 2228 15496
rect 2280 15444 2286 15496
rect 2774 15444 2780 15496
rect 2832 15444 2838 15496
rect 2976 15493 3004 15524
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 3605 15555 3663 15561
rect 3605 15521 3617 15555
rect 3651 15552 3663 15555
rect 3878 15552 3884 15564
rect 3651 15524 3884 15552
rect 3651 15521 3663 15524
rect 3605 15515 3663 15521
rect 3878 15512 3884 15524
rect 3936 15552 3942 15564
rect 4356 15552 4384 15592
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 6546 15580 6552 15632
rect 6604 15580 6610 15632
rect 6748 15620 6776 15660
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 7374 15688 7380 15700
rect 6880 15660 7380 15688
rect 6880 15648 6886 15660
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 7984 15660 8033 15688
rect 7984 15648 7990 15660
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 8386 15648 8392 15700
rect 8444 15688 8450 15700
rect 8754 15688 8760 15700
rect 8444 15660 8760 15688
rect 8444 15648 8450 15660
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 9769 15691 9827 15697
rect 9769 15688 9781 15691
rect 9548 15660 9781 15688
rect 9548 15648 9554 15660
rect 9769 15657 9781 15660
rect 9815 15657 9827 15691
rect 9769 15651 9827 15657
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 10229 15691 10287 15697
rect 10229 15688 10241 15691
rect 10100 15660 10241 15688
rect 10100 15648 10106 15660
rect 10229 15657 10241 15660
rect 10275 15657 10287 15691
rect 10229 15651 10287 15657
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 10870 15688 10876 15700
rect 10459 15660 10876 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 12158 15648 12164 15700
rect 12216 15648 12222 15700
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 12308 15660 13032 15688
rect 12308 15648 12314 15660
rect 7834 15620 7840 15632
rect 6748 15592 7840 15620
rect 7834 15580 7840 15592
rect 7892 15580 7898 15632
rect 8266 15592 9618 15620
rect 3936 15524 4384 15552
rect 3936 15512 3942 15524
rect 5074 15512 5080 15564
rect 5132 15512 5138 15564
rect 6178 15552 6184 15564
rect 5552 15524 6184 15552
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15453 3019 15487
rect 2961 15447 3019 15453
rect 3050 15444 3056 15496
rect 3108 15444 3114 15496
rect 3326 15444 3332 15496
rect 3384 15444 3390 15496
rect 3418 15444 3424 15496
rect 3476 15444 3482 15496
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15453 5227 15487
rect 5169 15447 5227 15453
rect 2792 15416 2820 15444
rect 3602 15416 3608 15428
rect 2792 15388 3608 15416
rect 3602 15376 3608 15388
rect 3660 15376 3666 15428
rect 4356 15416 4384 15447
rect 4706 15416 4712 15428
rect 4356 15388 4712 15416
rect 4706 15376 4712 15388
rect 4764 15416 4770 15428
rect 5184 15416 5212 15447
rect 5350 15444 5356 15496
rect 5408 15484 5414 15496
rect 5552 15493 5580 15524
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 6270 15512 6276 15564
rect 6328 15512 6334 15564
rect 6564 15552 6592 15580
rect 6914 15552 6920 15564
rect 6564 15524 6920 15552
rect 6914 15512 6920 15524
rect 6972 15552 6978 15564
rect 8266 15552 8294 15592
rect 6972 15524 7052 15552
rect 6972 15512 6978 15524
rect 5537 15487 5595 15493
rect 5537 15484 5549 15487
rect 5408 15456 5549 15484
rect 5408 15444 5414 15456
rect 5537 15453 5549 15456
rect 5583 15453 5595 15487
rect 5537 15447 5595 15453
rect 5626 15444 5632 15496
rect 5684 15444 5690 15496
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 6288 15484 6316 15512
rect 5859 15456 6316 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 5828 15416 5856 15447
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 7024 15493 7052 15524
rect 7760 15524 8294 15552
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6788 15456 6837 15484
rect 6788 15444 6794 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 7466 15444 7472 15496
rect 7524 15444 7530 15496
rect 7558 15444 7564 15496
rect 7616 15444 7622 15496
rect 7650 15444 7656 15496
rect 7708 15484 7714 15496
rect 7760 15493 7788 15524
rect 9122 15512 9128 15564
rect 9180 15552 9186 15564
rect 9309 15555 9367 15561
rect 9309 15552 9321 15555
rect 9180 15524 9321 15552
rect 9180 15512 9186 15524
rect 9309 15521 9321 15524
rect 9355 15521 9367 15555
rect 9309 15515 9367 15521
rect 9490 15512 9496 15564
rect 9548 15512 9554 15564
rect 9590 15552 9618 15592
rect 9674 15580 9680 15632
rect 9732 15620 9738 15632
rect 9858 15620 9864 15632
rect 9732 15592 9864 15620
rect 9732 15580 9738 15592
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 13004 15620 13032 15660
rect 13078 15648 13084 15700
rect 13136 15688 13142 15700
rect 15841 15691 15899 15697
rect 15841 15688 15853 15691
rect 13136 15660 15853 15688
rect 13136 15648 13142 15660
rect 15841 15657 15853 15660
rect 15887 15688 15899 15691
rect 15930 15688 15936 15700
rect 15887 15660 15936 15688
rect 15887 15657 15899 15660
rect 15841 15651 15899 15657
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 13004 15592 13952 15620
rect 11422 15552 11428 15564
rect 9590 15524 11428 15552
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 12253 15555 12311 15561
rect 12253 15552 12265 15555
rect 11716 15524 12265 15552
rect 11716 15496 11744 15524
rect 12253 15521 12265 15524
rect 12299 15521 12311 15555
rect 12253 15515 12311 15521
rect 13924 15552 13952 15592
rect 15102 15552 15108 15564
rect 13924 15524 15108 15552
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 7708 15456 7757 15484
rect 7708 15444 7714 15456
rect 7745 15453 7757 15456
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 7834 15444 7840 15496
rect 7892 15444 7898 15496
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 8481 15487 8539 15493
rect 8481 15484 8493 15487
rect 8444 15456 8493 15484
rect 8444 15444 8450 15456
rect 8481 15453 8493 15456
rect 8527 15484 8539 15487
rect 8938 15484 8944 15496
rect 8527 15456 8944 15484
rect 8527 15453 8539 15456
rect 8481 15447 8539 15453
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9398 15444 9404 15496
rect 9456 15444 9462 15496
rect 9585 15487 9643 15493
rect 9585 15453 9597 15487
rect 9631 15484 9643 15487
rect 9674 15484 9680 15496
rect 9631 15456 9680 15484
rect 9631 15453 9643 15456
rect 9585 15447 9643 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10318 15484 10324 15496
rect 10060 15456 10324 15484
rect 4764 15388 5856 15416
rect 6089 15419 6147 15425
rect 4764 15376 4770 15388
rect 6089 15385 6101 15419
rect 6135 15416 6147 15419
rect 6362 15416 6368 15428
rect 6135 15388 6368 15416
rect 6135 15385 6147 15388
rect 6089 15379 6147 15385
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 7098 15416 7104 15428
rect 7024 15388 7104 15416
rect 1946 15308 1952 15360
rect 2004 15348 2010 15360
rect 2041 15351 2099 15357
rect 2041 15348 2053 15351
rect 2004 15320 2053 15348
rect 2004 15308 2010 15320
rect 2041 15317 2053 15320
rect 2087 15348 2099 15351
rect 2130 15348 2136 15360
rect 2087 15320 2136 15348
rect 2087 15317 2099 15320
rect 2041 15311 2099 15317
rect 2130 15308 2136 15320
rect 2188 15308 2194 15360
rect 5166 15308 5172 15360
rect 5224 15348 5230 15360
rect 5994 15348 6000 15360
rect 5224 15320 6000 15348
rect 5224 15308 5230 15320
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 6733 15351 6791 15357
rect 6733 15317 6745 15351
rect 6779 15348 6791 15351
rect 6914 15348 6920 15360
rect 6779 15320 6920 15348
rect 6779 15317 6791 15320
rect 6733 15311 6791 15317
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 7024 15357 7052 15388
rect 7098 15376 7104 15388
rect 7156 15416 7162 15428
rect 9416 15416 9444 15444
rect 10060 15425 10088 15456
rect 10318 15444 10324 15456
rect 10376 15484 10382 15496
rect 10870 15484 10876 15496
rect 10376 15456 10876 15484
rect 10376 15444 10382 15456
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 11514 15484 11520 15496
rect 11112 15456 11520 15484
rect 11112 15444 11118 15456
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 11698 15444 11704 15496
rect 11756 15444 11762 15496
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 10045 15419 10103 15425
rect 7156 15388 9628 15416
rect 7156 15376 7162 15388
rect 9600 15360 9628 15388
rect 10045 15385 10057 15419
rect 10091 15385 10103 15419
rect 10045 15379 10103 15385
rect 10152 15388 10364 15416
rect 7009 15351 7067 15357
rect 7009 15317 7021 15351
rect 7055 15317 7067 15351
rect 7009 15311 7067 15317
rect 8110 15308 8116 15360
rect 8168 15348 8174 15360
rect 8389 15351 8447 15357
rect 8389 15348 8401 15351
rect 8168 15320 8401 15348
rect 8168 15308 8174 15320
rect 8389 15317 8401 15320
rect 8435 15348 8447 15351
rect 9030 15348 9036 15360
rect 8435 15320 9036 15348
rect 8435 15317 8447 15320
rect 8389 15311 8447 15317
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 9582 15308 9588 15360
rect 9640 15308 9646 15360
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 10152 15348 10180 15388
rect 10008 15320 10180 15348
rect 10008 15308 10014 15320
rect 10226 15308 10232 15360
rect 10284 15357 10290 15360
rect 10284 15351 10303 15357
rect 10291 15317 10303 15351
rect 10336 15348 10364 15388
rect 10410 15376 10416 15428
rect 10468 15416 10474 15428
rect 11238 15416 11244 15428
rect 10468 15388 11244 15416
rect 10468 15376 10474 15388
rect 11238 15376 11244 15388
rect 11296 15416 11302 15428
rect 11808 15416 11836 15447
rect 11882 15444 11888 15496
rect 11940 15444 11946 15496
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12437 15487 12495 15493
rect 12437 15484 12449 15487
rect 12216 15456 12449 15484
rect 12216 15444 12222 15456
rect 12437 15453 12449 15456
rect 12483 15453 12495 15487
rect 12437 15447 12495 15453
rect 12713 15487 12771 15493
rect 12713 15453 12725 15487
rect 12759 15484 12771 15487
rect 13354 15484 13360 15496
rect 12759 15456 13360 15484
rect 12759 15453 12771 15456
rect 12713 15447 12771 15453
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 13924 15493 13952 15524
rect 15102 15512 15108 15524
rect 15160 15512 15166 15564
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 16850 15552 16856 15564
rect 15712 15524 16856 15552
rect 15712 15512 15718 15524
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15453 13967 15487
rect 13909 15447 13967 15453
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 15933 15487 15991 15493
rect 15933 15484 15945 15487
rect 15896 15456 15945 15484
rect 15896 15444 15902 15456
rect 15933 15453 15945 15456
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 11296 15388 11836 15416
rect 11296 15376 11302 15388
rect 12526 15376 12532 15428
rect 12584 15416 12590 15428
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 12584 15388 14381 15416
rect 12584 15376 12590 15388
rect 14369 15385 14381 15388
rect 14415 15385 14427 15419
rect 14369 15379 14427 15385
rect 15378 15376 15384 15428
rect 15436 15376 15442 15428
rect 16206 15376 16212 15428
rect 16264 15376 16270 15428
rect 17862 15416 17868 15428
rect 17434 15388 17868 15416
rect 17862 15376 17868 15388
rect 17920 15376 17926 15428
rect 12250 15348 12256 15360
rect 10336 15320 12256 15348
rect 10284 15311 10303 15317
rect 10284 15308 10290 15311
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 12621 15351 12679 15357
rect 12621 15317 12633 15351
rect 12667 15348 12679 15351
rect 12894 15348 12900 15360
rect 12667 15320 12900 15348
rect 12667 15317 12679 15320
rect 12621 15311 12679 15317
rect 12894 15308 12900 15320
rect 12952 15348 12958 15360
rect 13446 15348 13452 15360
rect 12952 15320 13452 15348
rect 12952 15308 12958 15320
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 13817 15351 13875 15357
rect 13817 15317 13829 15351
rect 13863 15348 13875 15351
rect 14734 15348 14740 15360
rect 13863 15320 14740 15348
rect 13863 15317 13875 15320
rect 13817 15311 13875 15317
rect 14734 15308 14740 15320
rect 14792 15308 14798 15360
rect 17678 15308 17684 15360
rect 17736 15308 17742 15360
rect 1104 15258 18492 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 18492 15258
rect 1104 15184 18492 15206
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 5166 15144 5172 15156
rect 4120 15116 5172 15144
rect 4120 15104 4126 15116
rect 5166 15104 5172 15116
rect 5224 15104 5230 15156
rect 5350 15104 5356 15156
rect 5408 15104 5414 15156
rect 5994 15104 6000 15156
rect 6052 15144 6058 15156
rect 6822 15144 6828 15156
rect 6052 15116 6828 15144
rect 6052 15104 6058 15116
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7616 15116 7849 15144
rect 7616 15104 7622 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 9490 15104 9496 15156
rect 9548 15104 9554 15156
rect 9674 15104 9680 15156
rect 9732 15104 9738 15156
rect 10042 15104 10048 15156
rect 10100 15104 10106 15156
rect 10870 15144 10876 15156
rect 10152 15116 10876 15144
rect 4706 15036 4712 15088
rect 4764 15036 4770 15088
rect 8849 15079 8907 15085
rect 8849 15076 8861 15079
rect 5552 15048 8248 15076
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1636 14980 1685 15008
rect 1636 14968 1642 14980
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 2682 14968 2688 15020
rect 2740 14968 2746 15020
rect 2866 14968 2872 15020
rect 2924 14968 2930 15020
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 14977 3571 15011
rect 3513 14971 3571 14977
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 5258 15008 5264 15020
rect 4571 14980 5264 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 2406 14900 2412 14952
rect 2464 14940 2470 14952
rect 3528 14940 3556 14971
rect 2464 14912 3556 14940
rect 3712 14940 3740 14971
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 5552 15017 5580 15048
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 7006 15008 7012 15020
rect 6595 14980 7012 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 7006 14968 7012 14980
rect 7064 14968 7070 15020
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7282 15008 7288 15020
rect 7239 14980 7288 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 8110 14968 8116 15020
rect 8168 14968 8174 15020
rect 8220 14952 8248 15048
rect 8404 15048 8861 15076
rect 8404 15020 8432 15048
rect 8849 15045 8861 15048
rect 8895 15045 8907 15079
rect 8849 15039 8907 15045
rect 9122 15036 9128 15088
rect 9180 15076 9186 15088
rect 10152 15076 10180 15116
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14182 15144 14188 15156
rect 14139 15116 14188 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 14642 15104 14648 15156
rect 14700 15104 14706 15156
rect 16850 15104 16856 15156
rect 16908 15104 16914 15156
rect 12526 15076 12532 15088
rect 9180 15048 10180 15076
rect 10245 15048 12532 15076
rect 9180 15036 9186 15048
rect 8386 14968 8392 15020
rect 8444 14968 8450 15020
rect 8757 15011 8815 15017
rect 8757 15008 8769 15011
rect 8496 14980 8769 15008
rect 4154 14940 4160 14952
rect 3712 14912 4160 14940
rect 2464 14900 2470 14912
rect 3528 14872 3556 14912
rect 4154 14900 4160 14912
rect 4212 14940 4218 14952
rect 4798 14940 4804 14952
rect 4212 14912 4804 14940
rect 4212 14900 4218 14912
rect 4798 14900 4804 14912
rect 4856 14940 4862 14952
rect 6641 14943 6699 14949
rect 6641 14940 6653 14943
rect 4856 14912 6653 14940
rect 4856 14900 4862 14912
rect 6641 14909 6653 14912
rect 6687 14940 6699 14943
rect 6822 14940 6828 14952
rect 6687 14912 6828 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7742 14940 7748 14952
rect 6972 14912 7748 14940
rect 6972 14900 6978 14912
rect 7742 14900 7748 14912
rect 7800 14940 7806 14952
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 7800 14912 7849 14940
rect 7800 14900 7806 14912
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 8496 14940 8524 14980
rect 8757 14977 8769 14980
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 15008 8999 15011
rect 9309 15011 9367 15017
rect 8987 14980 9021 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 9309 14977 9321 15011
rect 9355 14977 9367 15011
rect 9309 14971 9367 14977
rect 8260 14912 8524 14940
rect 8665 14943 8723 14949
rect 8260 14900 8266 14912
rect 8665 14909 8677 14943
rect 8711 14940 8723 14943
rect 8956 14940 8984 14971
rect 9122 14940 9128 14952
rect 8711 14912 9128 14940
rect 8711 14909 8723 14912
rect 8665 14903 8723 14909
rect 9122 14900 9128 14912
rect 9180 14900 9186 14952
rect 9324 14884 9352 14971
rect 9490 14968 9496 15020
rect 9548 14968 9554 15020
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 9674 15008 9680 15020
rect 9631 14980 9680 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 15008 9827 15011
rect 9858 15008 9864 15020
rect 9815 14980 9864 15008
rect 9815 14977 9827 14980
rect 9769 14971 9827 14977
rect 9858 14968 9864 14980
rect 9916 14968 9922 15020
rect 10245 15017 10273 15048
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 13265 15079 13323 15085
rect 13265 15045 13277 15079
rect 13311 15076 13323 15079
rect 16868 15076 16896 15104
rect 13311 15048 13584 15076
rect 16868 15048 17356 15076
rect 13311 15045 13323 15048
rect 13265 15039 13323 15045
rect 10229 15011 10287 15017
rect 10229 14977 10241 15011
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 5077 14875 5135 14881
rect 3528 14844 4384 14872
rect 842 14764 848 14816
rect 900 14804 906 14816
rect 1489 14807 1547 14813
rect 1489 14804 1501 14807
rect 900 14776 1501 14804
rect 900 14764 906 14776
rect 1489 14773 1501 14776
rect 1535 14773 1547 14807
rect 1489 14767 1547 14773
rect 2866 14764 2872 14816
rect 2924 14764 2930 14816
rect 3418 14764 3424 14816
rect 3476 14804 3482 14816
rect 3513 14807 3571 14813
rect 3513 14804 3525 14807
rect 3476 14776 3525 14804
rect 3476 14764 3482 14776
rect 3513 14773 3525 14776
rect 3559 14773 3571 14807
rect 3513 14767 3571 14773
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 3660 14776 4261 14804
rect 3660 14764 3666 14776
rect 4249 14773 4261 14776
rect 4295 14773 4307 14807
rect 4356 14804 4384 14844
rect 5077 14841 5089 14875
rect 5123 14872 5135 14875
rect 5350 14872 5356 14884
rect 5123 14844 5356 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 5350 14832 5356 14844
rect 5408 14832 5414 14884
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 6546 14872 6552 14884
rect 5776 14844 6552 14872
rect 5776 14832 5782 14844
rect 6546 14832 6552 14844
rect 6604 14832 6610 14884
rect 6656 14844 7328 14872
rect 5736 14804 5764 14832
rect 6656 14813 6684 14844
rect 4356 14776 5764 14804
rect 6641 14807 6699 14813
rect 4249 14767 4307 14773
rect 6641 14773 6653 14807
rect 6687 14773 6699 14807
rect 6641 14767 6699 14773
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 6917 14807 6975 14813
rect 6917 14804 6929 14807
rect 6788 14776 6929 14804
rect 6788 14764 6794 14776
rect 6917 14773 6929 14776
rect 6963 14773 6975 14807
rect 6917 14767 6975 14773
rect 7190 14764 7196 14816
rect 7248 14764 7254 14816
rect 7300 14804 7328 14844
rect 7374 14832 7380 14884
rect 7432 14872 7438 14884
rect 7432 14844 8616 14872
rect 7432 14832 7438 14844
rect 7742 14804 7748 14816
rect 7300 14776 7748 14804
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 8588 14813 8616 14844
rect 9306 14832 9312 14884
rect 9364 14872 9370 14884
rect 10244 14872 10272 14971
rect 10318 14968 10324 15020
rect 10376 14968 10382 15020
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 12158 15008 12164 15020
rect 10643 14980 12164 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 12158 14968 12164 14980
rect 12216 15008 12222 15020
rect 12802 15008 12808 15020
rect 12216 14980 12808 15008
rect 12216 14968 12222 14980
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 13078 14968 13084 15020
rect 13136 14968 13142 15020
rect 13556 15017 13584 15048
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11698 14940 11704 14952
rect 10744 14912 11704 14940
rect 10744 14900 10750 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 12894 14900 12900 14952
rect 12952 14900 12958 14952
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 9364 14844 10272 14872
rect 10336 14844 12112 14872
rect 9364 14832 9370 14844
rect 8021 14807 8079 14813
rect 8021 14773 8033 14807
rect 8067 14804 8079 14807
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 8067 14776 8217 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 8573 14807 8631 14813
rect 8573 14773 8585 14807
rect 8619 14804 8631 14807
rect 10336 14804 10364 14844
rect 8619 14776 10364 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 11054 14804 11060 14816
rect 10468 14776 11060 14804
rect 10468 14764 10474 14776
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 12084 14804 12112 14844
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 13004 14872 13032 14903
rect 13446 14900 13452 14952
rect 13504 14940 13510 14952
rect 14292 14940 14320 14971
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 14424 14980 14565 15008
rect 14424 14968 14430 14980
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 13504 14912 14320 14940
rect 13504 14900 13510 14912
rect 14292 14872 14320 14912
rect 14458 14900 14464 14952
rect 14516 14900 14522 14952
rect 14568 14940 14596 14971
rect 14918 14968 14924 15020
rect 14976 15008 14982 15020
rect 15013 15011 15071 15017
rect 15013 15008 15025 15011
rect 14976 14980 15025 15008
rect 14976 14968 14982 14980
rect 15013 14977 15025 14980
rect 15059 14977 15071 15011
rect 15013 14971 15071 14977
rect 15841 15011 15899 15017
rect 15841 14977 15853 15011
rect 15887 15008 15899 15011
rect 16022 15008 16028 15020
rect 15887 14980 16028 15008
rect 15887 14977 15899 14980
rect 15841 14971 15899 14977
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 16942 15017 16948 15020
rect 16911 15011 16948 15017
rect 16911 14977 16923 15011
rect 16911 14971 16948 14977
rect 16942 14968 16948 14971
rect 17000 14968 17006 15020
rect 17328 15017 17356 15048
rect 17313 15011 17371 15017
rect 17313 14977 17325 15011
rect 17359 14977 17371 15011
rect 17313 14971 17371 14977
rect 15657 14943 15715 14949
rect 15657 14940 15669 14943
rect 14568 14912 15669 14940
rect 15657 14909 15669 14912
rect 15703 14909 15715 14943
rect 15657 14903 15715 14909
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 17221 14943 17279 14949
rect 17221 14940 17233 14943
rect 16816 14912 17233 14940
rect 16816 14900 16822 14912
rect 17221 14909 17233 14912
rect 17267 14909 17279 14943
rect 17221 14903 17279 14909
rect 15562 14872 15568 14884
rect 12216 14844 14228 14872
rect 14292 14844 15568 14872
rect 12216 14832 12222 14844
rect 12342 14804 12348 14816
rect 12084 14776 12348 14804
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 12676 14776 13369 14804
rect 12676 14764 12682 14776
rect 13357 14773 13369 14776
rect 13403 14773 13415 14807
rect 14200 14804 14228 14844
rect 15562 14832 15568 14844
rect 15620 14832 15626 14884
rect 16666 14832 16672 14884
rect 16724 14832 16730 14884
rect 14458 14804 14464 14816
rect 14200 14776 14464 14804
rect 13357 14767 13415 14773
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 1104 14714 18492 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 18492 14714
rect 1104 14640 18492 14662
rect 1578 14560 1584 14612
rect 1636 14560 1642 14612
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 3384 14572 3433 14600
rect 3384 14560 3390 14572
rect 3421 14569 3433 14572
rect 3467 14569 3479 14603
rect 3421 14563 3479 14569
rect 3528 14572 4660 14600
rect 1946 14492 1952 14544
rect 2004 14532 2010 14544
rect 2133 14535 2191 14541
rect 2133 14532 2145 14535
rect 2004 14504 2145 14532
rect 2004 14492 2010 14504
rect 2133 14501 2145 14504
rect 2179 14501 2191 14535
rect 2133 14495 2191 14501
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14464 2099 14467
rect 2498 14464 2504 14476
rect 2087 14436 2504 14464
rect 2087 14433 2099 14436
rect 2041 14427 2099 14433
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 2866 14464 2872 14476
rect 2792 14436 2872 14464
rect 1762 14356 1768 14408
rect 1820 14356 1826 14408
rect 1854 14356 1860 14408
rect 1912 14396 1918 14408
rect 1949 14399 2007 14405
rect 1949 14396 1961 14399
rect 1912 14368 1961 14396
rect 1912 14356 1918 14368
rect 1949 14365 1961 14368
rect 1995 14365 2007 14399
rect 2406 14396 2412 14408
rect 1949 14359 2007 14365
rect 2240 14368 2412 14396
rect 2130 14288 2136 14340
rect 2188 14288 2194 14340
rect 2038 14220 2044 14272
rect 2096 14260 2102 14272
rect 2240 14260 2268 14368
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2792 14405 2820 14436
rect 2866 14424 2872 14436
rect 2924 14464 2930 14476
rect 3528 14464 3556 14572
rect 3970 14492 3976 14544
rect 4028 14532 4034 14544
rect 4430 14532 4436 14544
rect 4028 14504 4436 14532
rect 4028 14492 4034 14504
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 4632 14532 4660 14572
rect 4706 14560 4712 14612
rect 4764 14560 4770 14612
rect 6365 14603 6423 14609
rect 6365 14569 6377 14603
rect 6411 14600 6423 14603
rect 7282 14600 7288 14612
rect 6411 14572 7288 14600
rect 6411 14569 6423 14572
rect 6365 14563 6423 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14569 7435 14603
rect 7377 14563 7435 14569
rect 4798 14532 4804 14544
rect 4632 14504 4804 14532
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 5077 14535 5135 14541
rect 5077 14501 5089 14535
rect 5123 14532 5135 14535
rect 5350 14532 5356 14544
rect 5123 14504 5356 14532
rect 5123 14501 5135 14504
rect 5077 14495 5135 14501
rect 5350 14492 5356 14504
rect 5408 14492 5414 14544
rect 2924 14436 3556 14464
rect 2924 14424 2930 14436
rect 3602 14424 3608 14476
rect 3660 14464 3666 14476
rect 3786 14464 3792 14476
rect 3660 14436 3792 14464
rect 3660 14424 3666 14436
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 4157 14467 4215 14473
rect 4157 14464 4169 14467
rect 3896 14436 4169 14464
rect 2777 14399 2835 14405
rect 2777 14365 2789 14399
rect 2823 14365 2835 14399
rect 2777 14359 2835 14365
rect 2958 14356 2964 14408
rect 3016 14356 3022 14408
rect 3050 14356 3056 14408
rect 3108 14356 3114 14408
rect 3142 14356 3148 14408
rect 3200 14356 3206 14408
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14365 3295 14399
rect 3237 14359 3295 14365
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14396 3387 14399
rect 3896 14396 3924 14436
rect 4157 14433 4169 14436
rect 4203 14464 4215 14467
rect 6457 14467 6515 14473
rect 4203 14436 4384 14464
rect 4203 14433 4215 14436
rect 4157 14427 4215 14433
rect 3375 14368 3924 14396
rect 3973 14399 4031 14405
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 2866 14288 2872 14340
rect 2924 14328 2930 14340
rect 3068 14328 3096 14356
rect 2924 14300 3096 14328
rect 3252 14328 3280 14359
rect 3789 14331 3847 14337
rect 3789 14328 3801 14331
rect 3252 14300 3801 14328
rect 2924 14288 2930 14300
rect 3789 14297 3801 14300
rect 3835 14297 3847 14331
rect 3789 14291 3847 14297
rect 3878 14288 3884 14340
rect 3936 14328 3942 14340
rect 3988 14328 4016 14359
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4172 14368 4261 14396
rect 3936 14300 4016 14328
rect 3936 14288 3942 14300
rect 2096 14232 2268 14260
rect 2096 14220 2102 14232
rect 2314 14220 2320 14272
rect 2372 14220 2378 14272
rect 2590 14220 2596 14272
rect 2648 14220 2654 14272
rect 3605 14263 3663 14269
rect 3605 14229 3617 14263
rect 3651 14260 3663 14263
rect 4172 14260 4200 14368
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 3651 14232 4200 14260
rect 4356 14260 4384 14436
rect 6457 14433 6469 14467
rect 6503 14464 6515 14467
rect 7006 14464 7012 14476
rect 6503 14436 7012 14464
rect 6503 14433 6515 14436
rect 6457 14427 6515 14433
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 7190 14424 7196 14476
rect 7248 14424 7254 14476
rect 7392 14464 7420 14563
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7524 14572 7665 14600
rect 7524 14560 7530 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 10134 14600 10140 14612
rect 10091 14572 10140 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10962 14560 10968 14612
rect 11020 14560 11026 14612
rect 12066 14560 12072 14612
rect 12124 14560 12130 14612
rect 14645 14603 14703 14609
rect 14645 14569 14657 14603
rect 14691 14600 14703 14603
rect 15378 14600 15384 14612
rect 14691 14572 15384 14600
rect 14691 14569 14703 14572
rect 14645 14563 14703 14569
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 16482 14600 16488 14612
rect 15795 14572 16488 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 16482 14560 16488 14572
rect 16540 14560 16546 14612
rect 17862 14560 17868 14612
rect 17920 14560 17926 14612
rect 7561 14535 7619 14541
rect 7561 14501 7573 14535
rect 7607 14532 7619 14535
rect 7607 14504 8432 14532
rect 7607 14501 7619 14504
rect 7561 14495 7619 14501
rect 8404 14473 8432 14504
rect 8478 14492 8484 14544
rect 8536 14492 8542 14544
rect 8573 14535 8631 14541
rect 8573 14501 8585 14535
rect 8619 14532 8631 14535
rect 11606 14532 11612 14544
rect 8619 14504 11612 14532
rect 8619 14501 8631 14504
rect 8573 14495 8631 14501
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 12437 14535 12495 14541
rect 12437 14501 12449 14535
rect 12483 14532 12495 14535
rect 12621 14535 12679 14541
rect 12621 14532 12633 14535
rect 12483 14504 12633 14532
rect 12483 14501 12495 14504
rect 12437 14495 12495 14501
rect 12621 14501 12633 14504
rect 12667 14501 12679 14535
rect 12621 14495 12679 14501
rect 12802 14492 12808 14544
rect 12860 14532 12866 14544
rect 12860 14504 12940 14532
rect 12860 14492 12866 14504
rect 12912 14473 12940 14504
rect 14826 14492 14832 14544
rect 14884 14492 14890 14544
rect 8389 14467 8447 14473
rect 7392 14436 8248 14464
rect 4430 14356 4436 14408
rect 4488 14356 4494 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 4856 14368 5764 14396
rect 4856 14356 4862 14368
rect 4709 14331 4767 14337
rect 4709 14297 4721 14331
rect 4755 14328 4767 14331
rect 5626 14328 5632 14340
rect 4755 14300 5632 14328
rect 4755 14297 4767 14300
rect 4709 14291 4767 14297
rect 5626 14288 5632 14300
rect 5684 14288 5690 14340
rect 5736 14328 5764 14368
rect 5994 14356 6000 14408
rect 6052 14356 6058 14408
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 7466 14396 7472 14408
rect 7423 14368 7472 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 7944 14405 7972 14436
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 6917 14331 6975 14337
rect 6917 14328 6929 14331
rect 5736 14300 6929 14328
rect 6917 14297 6929 14300
rect 6963 14297 6975 14331
rect 6917 14291 6975 14297
rect 4522 14260 4528 14272
rect 4356 14232 4528 14260
rect 3651 14229 3663 14232
rect 3605 14223 3663 14229
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 5258 14220 5264 14272
rect 5316 14260 5322 14272
rect 5721 14263 5779 14269
rect 5721 14260 5733 14263
rect 5316 14232 5733 14260
rect 5316 14220 5322 14232
rect 5721 14229 5733 14232
rect 5767 14229 5779 14263
rect 5721 14223 5779 14229
rect 6086 14220 6092 14272
rect 6144 14220 6150 14272
rect 6181 14263 6239 14269
rect 6181 14229 6193 14263
rect 6227 14260 6239 14263
rect 6454 14260 6460 14272
rect 6227 14232 6460 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6454 14220 6460 14232
rect 6512 14220 6518 14272
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 8036 14260 8064 14359
rect 8110 14356 8116 14408
rect 8168 14356 8174 14408
rect 8220 14328 8248 14436
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 12897 14467 12955 14473
rect 8389 14427 8447 14433
rect 8588 14436 12664 14464
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8478 14396 8484 14408
rect 8343 14368 8484 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 8588 14328 8616 14436
rect 12636 14408 12664 14436
rect 12897 14433 12909 14467
rect 12943 14464 12955 14467
rect 12986 14464 12992 14476
rect 12943 14436 12992 14464
rect 12943 14433 12955 14436
rect 12897 14427 12955 14433
rect 12986 14424 12992 14436
rect 13044 14424 13050 14476
rect 16574 14464 16580 14476
rect 14568 14436 16580 14464
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 8754 14396 8760 14408
rect 8711 14368 8760 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 9490 14356 9496 14408
rect 9548 14396 9554 14408
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 9548 14368 10241 14396
rect 9548 14356 9554 14368
rect 10229 14365 10241 14368
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 8220 14300 8616 14328
rect 9030 14288 9036 14340
rect 9088 14288 9094 14340
rect 9950 14288 9956 14340
rect 10008 14328 10014 14340
rect 10336 14328 10364 14359
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 10502 14356 10508 14408
rect 10560 14356 10566 14408
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14396 10839 14399
rect 11330 14396 11336 14408
rect 10827 14368 11336 14396
rect 10827 14365 10839 14368
rect 10781 14359 10839 14365
rect 10704 14328 10732 14359
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 12250 14356 12256 14408
rect 12308 14356 12314 14408
rect 12342 14356 12348 14408
rect 12400 14396 12406 14408
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 12400 14368 12541 14396
rect 12400 14356 12406 14368
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12618 14356 12624 14408
rect 12676 14356 12682 14408
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14396 12771 14399
rect 12802 14396 12808 14408
rect 12759 14368 12808 14396
rect 12759 14365 12771 14368
rect 12713 14359 12771 14365
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 14568 14405 14596 14436
rect 16574 14424 16580 14436
rect 16632 14464 16638 14476
rect 16632 14436 17816 14464
rect 16632 14424 16638 14436
rect 17788 14408 17816 14436
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 17770 14356 17776 14408
rect 17828 14356 17834 14408
rect 10008 14300 10732 14328
rect 10008 14288 10014 14300
rect 10962 14288 10968 14340
rect 11020 14288 11026 14340
rect 11146 14288 11152 14340
rect 11204 14328 11210 14340
rect 14090 14328 14096 14340
rect 11204 14300 14096 14328
rect 11204 14288 11210 14300
rect 14090 14288 14096 14300
rect 14148 14288 14154 14340
rect 15010 14288 15016 14340
rect 15068 14288 15074 14340
rect 15197 14331 15255 14337
rect 15197 14297 15209 14331
rect 15243 14328 15255 14331
rect 16574 14328 16580 14340
rect 15243 14300 16580 14328
rect 15243 14297 15255 14300
rect 15197 14291 15255 14297
rect 16574 14288 16580 14300
rect 16632 14288 16638 14340
rect 17037 14331 17095 14337
rect 17037 14297 17049 14331
rect 17083 14328 17095 14331
rect 17954 14328 17960 14340
rect 17083 14300 17960 14328
rect 17083 14297 17095 14300
rect 17037 14291 17095 14297
rect 17954 14288 17960 14300
rect 18012 14288 18018 14340
rect 6788 14232 8064 14260
rect 6788 14220 6794 14232
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 8846 14260 8852 14272
rect 8536 14232 8852 14260
rect 8536 14220 8542 14232
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9122 14220 9128 14272
rect 9180 14220 9186 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 11422 14260 11428 14272
rect 9272 14232 11428 14260
rect 9272 14220 9278 14232
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 11514 14220 11520 14272
rect 11572 14260 11578 14272
rect 13170 14260 13176 14272
rect 11572 14232 13176 14260
rect 11572 14220 11578 14232
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 1104 14170 18492 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 18492 14170
rect 1104 14096 18492 14118
rect 1946 14016 1952 14068
rect 2004 14016 2010 14068
rect 2777 14059 2835 14065
rect 2777 14025 2789 14059
rect 2823 14056 2835 14059
rect 3142 14056 3148 14068
rect 2823 14028 3148 14056
rect 2823 14025 2835 14028
rect 2777 14019 2835 14025
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 6089 14059 6147 14065
rect 3804 14028 5120 14056
rect 1857 13991 1915 13997
rect 1857 13957 1869 13991
rect 1903 13988 1915 13991
rect 2130 13988 2136 14000
rect 1903 13960 2136 13988
rect 1903 13957 1915 13960
rect 1857 13951 1915 13957
rect 2130 13948 2136 13960
rect 2188 13948 2194 14000
rect 2406 13948 2412 14000
rect 2464 13948 2470 14000
rect 2625 13991 2683 13997
rect 2625 13957 2637 13991
rect 2671 13988 2683 13991
rect 2958 13988 2964 14000
rect 2671 13960 2964 13988
rect 2671 13957 2683 13960
rect 2625 13951 2683 13957
rect 2958 13948 2964 13960
rect 3016 13948 3022 14000
rect 3234 13988 3240 14000
rect 3068 13960 3240 13988
rect 2314 13880 2320 13932
rect 2372 13920 2378 13932
rect 3068 13929 3096 13960
rect 3234 13948 3240 13960
rect 3292 13948 3298 14000
rect 3697 13991 3755 13997
rect 3697 13988 3709 13991
rect 3344 13960 3709 13988
rect 3344 13932 3372 13960
rect 3697 13957 3709 13960
rect 3743 13957 3755 13991
rect 3697 13951 3755 13957
rect 3053 13923 3111 13929
rect 2372 13892 2728 13920
rect 2372 13880 2378 13892
rect 1854 13812 1860 13864
rect 1912 13852 1918 13864
rect 2038 13852 2044 13864
rect 1912 13824 2044 13852
rect 1912 13812 1918 13824
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 2590 13852 2596 13864
rect 2179 13824 2596 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 2700 13852 2728 13892
rect 3053 13889 3065 13923
rect 3099 13889 3111 13923
rect 3053 13883 3111 13889
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3191 13892 3280 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3252 13852 3280 13892
rect 3326 13880 3332 13932
rect 3384 13880 3390 13932
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13920 3479 13923
rect 3510 13920 3516 13932
rect 3467 13892 3516 13920
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 3510 13880 3516 13892
rect 3568 13920 3574 13932
rect 3804 13920 3832 14028
rect 4706 13988 4712 14000
rect 4448 13960 4712 13988
rect 3568 13892 3832 13920
rect 3568 13880 3574 13892
rect 3878 13880 3884 13932
rect 3936 13880 3942 13932
rect 4062 13880 4068 13932
rect 4120 13880 4126 13932
rect 4448 13929 4476 13960
rect 4706 13948 4712 13960
rect 4764 13948 4770 14000
rect 5092 13932 5120 14028
rect 6089 14025 6101 14059
rect 6135 14056 6147 14059
rect 6270 14056 6276 14068
rect 6135 14028 6276 14056
rect 6135 14025 6147 14028
rect 6089 14019 6147 14025
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 7190 14056 7196 14068
rect 6880 14028 7196 14056
rect 6880 14016 6886 14028
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 7469 14059 7527 14065
rect 7469 14025 7481 14059
rect 7515 14056 7527 14059
rect 8110 14056 8116 14068
rect 7515 14028 8116 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 8573 14059 8631 14065
rect 8573 14056 8585 14059
rect 8352 14028 8585 14056
rect 8352 14016 8358 14028
rect 8573 14025 8585 14028
rect 8619 14025 8631 14059
rect 8573 14019 8631 14025
rect 9858 14016 9864 14068
rect 9916 14016 9922 14068
rect 9950 14016 9956 14068
rect 10008 14016 10014 14068
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 10560 14028 11345 14056
rect 10560 14016 10566 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 11606 14016 11612 14068
rect 11664 14016 11670 14068
rect 11977 14059 12035 14065
rect 11977 14025 11989 14059
rect 12023 14056 12035 14059
rect 12066 14056 12072 14068
rect 12023 14028 12072 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 12066 14016 12072 14028
rect 12124 14056 12130 14068
rect 12342 14056 12348 14068
rect 12124 14028 12348 14056
rect 12124 14016 12130 14028
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12894 14016 12900 14068
rect 12952 14016 12958 14068
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 13964 14028 14105 14056
rect 13964 14016 13970 14028
rect 14093 14025 14105 14028
rect 14139 14025 14151 14059
rect 14093 14019 14151 14025
rect 14274 14016 14280 14068
rect 14332 14016 14338 14068
rect 15749 14059 15807 14065
rect 15749 14025 15761 14059
rect 15795 14056 15807 14059
rect 16206 14056 16212 14068
rect 15795 14028 16212 14056
rect 15795 14025 15807 14028
rect 15749 14019 15807 14025
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 17770 14016 17776 14068
rect 17828 14016 17834 14068
rect 6641 13991 6699 13997
rect 6641 13988 6653 13991
rect 6104 13960 6653 13988
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 2700 13824 3280 13852
rect 2869 13787 2927 13793
rect 2869 13784 2881 13787
rect 2746 13756 2881 13784
rect 1489 13719 1547 13725
rect 1489 13685 1501 13719
rect 1535 13716 1547 13719
rect 1670 13716 1676 13728
rect 1535 13688 1676 13716
rect 1535 13685 1547 13688
rect 1489 13679 1547 13685
rect 1670 13676 1676 13688
rect 1728 13676 1734 13728
rect 2593 13719 2651 13725
rect 2593 13685 2605 13719
rect 2639 13716 2651 13719
rect 2746 13716 2774 13756
rect 2869 13753 2881 13756
rect 2915 13753 2927 13787
rect 3252 13784 3280 13824
rect 3602 13812 3608 13864
rect 3660 13852 3666 13864
rect 4264 13852 4292 13883
rect 4522 13880 4528 13932
rect 4580 13920 4586 13932
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4580 13892 4905 13920
rect 4580 13880 4586 13892
rect 4893 13889 4905 13892
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5074 13880 5080 13932
rect 5132 13880 5138 13932
rect 5905 13923 5963 13929
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 5994 13920 6000 13932
rect 5951 13892 6000 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 6104 13864 6132 13960
rect 6641 13957 6653 13960
rect 6687 13957 6699 13991
rect 6641 13951 6699 13957
rect 6730 13948 6736 14000
rect 6788 13948 6794 14000
rect 8478 13988 8484 14000
rect 6840 13960 8484 13988
rect 6178 13880 6184 13932
rect 6236 13880 6242 13932
rect 6544 13923 6602 13929
rect 6544 13889 6556 13923
rect 6590 13920 6602 13923
rect 6840 13920 6868 13960
rect 8478 13948 8484 13960
rect 8536 13948 8542 14000
rect 8941 13991 8999 13997
rect 8941 13988 8953 13991
rect 8588 13960 8953 13988
rect 6590 13892 6868 13920
rect 6916 13923 6974 13929
rect 6590 13889 6602 13892
rect 6544 13883 6602 13889
rect 6916 13889 6928 13923
rect 6962 13889 6974 13923
rect 6916 13883 6974 13889
rect 3660 13824 4292 13852
rect 4617 13855 4675 13861
rect 3660 13812 3666 13824
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 4706 13852 4712 13864
rect 4663 13824 4712 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 4706 13812 4712 13824
rect 4764 13852 4770 13864
rect 4985 13855 5043 13861
rect 4764 13824 4936 13852
rect 4764 13812 4770 13824
rect 4798 13784 4804 13796
rect 3252 13756 4804 13784
rect 2869 13747 2927 13753
rect 4798 13744 4804 13756
rect 4856 13744 4862 13796
rect 4908 13784 4936 13824
rect 4985 13821 4997 13855
rect 5031 13852 5043 13855
rect 5626 13852 5632 13864
rect 5031 13824 5632 13852
rect 5031 13821 5043 13824
rect 4985 13815 5043 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 5718 13812 5724 13864
rect 5776 13812 5782 13864
rect 6086 13812 6092 13864
rect 6144 13812 6150 13864
rect 6931 13796 6959 13883
rect 7006 13880 7012 13932
rect 7064 13880 7070 13932
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13920 7159 13923
rect 7742 13920 7748 13932
rect 7147 13892 7748 13920
rect 7147 13889 7159 13892
rect 7101 13883 7159 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8588 13920 8616 13960
rect 8941 13957 8953 13960
rect 8987 13957 8999 13991
rect 9876 13988 9904 14016
rect 12250 13988 12256 14000
rect 9876 13960 9996 13988
rect 8941 13951 8999 13957
rect 9968 13932 9996 13960
rect 10060 13960 12256 13988
rect 10060 13932 10088 13960
rect 12250 13948 12256 13960
rect 12308 13948 12314 14000
rect 13170 13948 13176 14000
rect 13228 13988 13234 14000
rect 15381 13991 15439 13997
rect 15381 13988 15393 13991
rect 13228 13960 15393 13988
rect 13228 13948 13234 13960
rect 15381 13957 15393 13960
rect 15427 13988 15439 13991
rect 16390 13988 16396 14000
rect 15427 13960 16396 13988
rect 15427 13957 15439 13960
rect 15381 13951 15439 13957
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 18046 13948 18052 14000
rect 18104 13948 18110 14000
rect 8168 13892 8616 13920
rect 8168 13880 8174 13892
rect 8754 13880 8760 13932
rect 8812 13880 8818 13932
rect 9030 13880 9036 13932
rect 9088 13880 9094 13932
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 9585 13923 9643 13929
rect 9585 13920 9597 13923
rect 9180 13892 9597 13920
rect 9180 13880 9186 13892
rect 9585 13889 9597 13892
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 9858 13880 9864 13932
rect 9916 13880 9922 13932
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 10042 13880 10048 13932
rect 10100 13880 10106 13932
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13920 10195 13923
rect 10778 13920 10784 13932
rect 10183 13892 10784 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 11054 13880 11060 13932
rect 11112 13880 11118 13932
rect 11514 13920 11520 13932
rect 11348 13892 11520 13920
rect 7193 13855 7251 13861
rect 7193 13821 7205 13855
rect 7239 13852 7251 13855
rect 7558 13852 7564 13864
rect 7239 13824 7564 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 7760 13824 10364 13852
rect 4908 13756 6776 13784
rect 2639 13688 2774 13716
rect 2639 13685 2651 13688
rect 2593 13679 2651 13685
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 6362 13716 6368 13728
rect 5868 13688 6368 13716
rect 5868 13676 5874 13688
rect 6362 13676 6368 13688
rect 6420 13676 6426 13728
rect 6748 13716 6776 13756
rect 6914 13744 6920 13796
rect 6972 13744 6978 13796
rect 7760 13784 7788 13824
rect 7020 13756 7788 13784
rect 6822 13716 6828 13728
rect 6748 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13716 6886 13728
rect 7020 13716 7048 13756
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 9858 13784 9864 13796
rect 8076 13756 9864 13784
rect 8076 13744 8082 13756
rect 9858 13744 9864 13756
rect 9916 13784 9922 13796
rect 10226 13784 10232 13796
rect 9916 13756 10232 13784
rect 9916 13744 9922 13756
rect 10226 13744 10232 13756
rect 10284 13744 10290 13796
rect 10336 13784 10364 13824
rect 10410 13812 10416 13864
rect 10468 13812 10474 13864
rect 11348 13861 11376 13892
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 11698 13880 11704 13932
rect 11756 13880 11762 13932
rect 12158 13880 12164 13932
rect 12216 13880 12222 13932
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13920 12587 13923
rect 12618 13920 12624 13932
rect 12575 13892 12624 13920
rect 12575 13889 12587 13892
rect 12529 13883 12587 13889
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13889 12771 13923
rect 12713 13883 12771 13889
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 12342 13812 12348 13864
rect 12400 13812 12406 13864
rect 12728 13852 12756 13883
rect 12802 13880 12808 13932
rect 12860 13880 12866 13932
rect 12986 13880 12992 13932
rect 13044 13880 13050 13932
rect 13998 13880 14004 13932
rect 14056 13880 14062 13932
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13920 14427 13923
rect 14458 13920 14464 13932
rect 14415 13892 14464 13920
rect 14415 13889 14427 13892
rect 14369 13883 14427 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 15286 13880 15292 13932
rect 15344 13880 15350 13932
rect 15470 13880 15476 13932
rect 15528 13880 15534 13932
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13889 15715 13923
rect 15657 13883 15715 13889
rect 13004 13852 13032 13880
rect 12728 13824 13032 13852
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 14918 13852 14924 13864
rect 14240 13824 14924 13852
rect 14240 13812 14246 13824
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 15672 13852 15700 13883
rect 16758 13880 16764 13932
rect 16816 13880 16822 13932
rect 17589 13923 17647 13929
rect 17589 13920 17601 13923
rect 16960 13892 17601 13920
rect 16850 13852 16856 13864
rect 15068 13824 16856 13852
rect 15068 13812 15074 13824
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 12360 13784 12388 13812
rect 10336 13756 12388 13784
rect 12434 13744 12440 13796
rect 12492 13784 12498 13796
rect 13078 13784 13084 13796
rect 12492 13756 13084 13784
rect 12492 13744 12498 13756
rect 13078 13744 13084 13756
rect 13136 13784 13142 13796
rect 13814 13784 13820 13796
rect 13136 13756 13820 13784
rect 13136 13744 13142 13756
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 13906 13744 13912 13796
rect 13964 13784 13970 13796
rect 14550 13784 14556 13796
rect 13964 13756 14556 13784
rect 13964 13744 13970 13756
rect 14550 13744 14556 13756
rect 14608 13744 14614 13796
rect 15562 13744 15568 13796
rect 15620 13784 15626 13796
rect 16960 13784 16988 13892
rect 17589 13889 17601 13892
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 15620 13756 16988 13784
rect 15620 13744 15626 13756
rect 6880 13688 7048 13716
rect 6880 13676 6886 13688
rect 7282 13676 7288 13728
rect 7340 13676 7346 13728
rect 8294 13676 8300 13728
rect 8352 13716 8358 13728
rect 9309 13719 9367 13725
rect 9309 13716 9321 13719
rect 8352 13688 9321 13716
rect 8352 13676 8358 13688
rect 9309 13685 9321 13688
rect 9355 13685 9367 13719
rect 9309 13679 9367 13685
rect 11146 13676 11152 13728
rect 11204 13676 11210 13728
rect 12158 13676 12164 13728
rect 12216 13716 12222 13728
rect 12342 13716 12348 13728
rect 12216 13688 12348 13716
rect 12216 13676 12222 13688
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12618 13676 12624 13728
rect 12676 13716 12682 13728
rect 13630 13716 13636 13728
rect 12676 13688 13636 13716
rect 12676 13676 12682 13688
rect 13630 13676 13636 13688
rect 13688 13716 13694 13728
rect 14458 13716 14464 13728
rect 13688 13688 14464 13716
rect 13688 13676 13694 13688
rect 14458 13676 14464 13688
rect 14516 13716 14522 13728
rect 17129 13719 17187 13725
rect 17129 13716 17141 13719
rect 14516 13688 17141 13716
rect 14516 13676 14522 13688
rect 17129 13685 17141 13688
rect 17175 13685 17187 13719
rect 17129 13679 17187 13685
rect 1104 13626 18492 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 18492 13626
rect 1104 13552 18492 13574
rect 1302 13472 1308 13524
rect 1360 13512 1366 13524
rect 1489 13515 1547 13521
rect 1489 13512 1501 13515
rect 1360 13484 1501 13512
rect 1360 13472 1366 13484
rect 1489 13481 1501 13484
rect 1535 13481 1547 13515
rect 1489 13475 1547 13481
rect 2406 13472 2412 13524
rect 2464 13472 2470 13524
rect 3142 13472 3148 13524
rect 3200 13512 3206 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3200 13484 3801 13512
rect 3200 13472 3206 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 3789 13475 3847 13481
rect 4172 13484 5948 13512
rect 4172 13444 4200 13484
rect 4706 13444 4712 13456
rect 2746 13416 4200 13444
rect 4264 13416 4712 13444
rect 1670 13268 1676 13320
rect 1728 13268 1734 13320
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13308 2651 13311
rect 2746 13308 2774 13416
rect 3786 13336 3792 13388
rect 3844 13376 3850 13388
rect 3970 13376 3976 13388
rect 3844 13348 3976 13376
rect 3844 13336 3850 13348
rect 3970 13336 3976 13348
rect 4028 13336 4034 13388
rect 4264 13376 4292 13416
rect 4706 13404 4712 13416
rect 4764 13404 4770 13456
rect 4172 13348 4292 13376
rect 4433 13379 4491 13385
rect 2639 13280 2774 13308
rect 2869 13311 2927 13317
rect 2639 13277 2651 13280
rect 2593 13271 2651 13277
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 3142 13308 3148 13320
rect 2915 13280 3148 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3234 13268 3240 13320
rect 3292 13308 3298 13320
rect 4172 13317 4200 13348
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4798 13376 4804 13388
rect 4479 13348 4804 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 4798 13336 4804 13348
rect 4856 13376 4862 13388
rect 5442 13376 5448 13388
rect 4856 13348 5448 13376
rect 4856 13336 4862 13348
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 5920 13376 5948 13484
rect 5994 13472 6000 13524
rect 6052 13472 6058 13524
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13512 6423 13515
rect 6914 13512 6920 13524
rect 6411 13484 6920 13512
rect 6411 13481 6423 13484
rect 6365 13475 6423 13481
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 8754 13472 8760 13524
rect 8812 13472 8818 13524
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 9088 13484 9505 13512
rect 9088 13472 9094 13484
rect 9493 13481 9505 13484
rect 9539 13481 9551 13515
rect 9493 13475 9551 13481
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 10318 13512 10324 13524
rect 9824 13484 10324 13512
rect 9824 13472 9830 13484
rect 10318 13472 10324 13484
rect 10376 13512 10382 13524
rect 13725 13515 13783 13521
rect 10376 13484 13676 13512
rect 10376 13472 10382 13484
rect 6270 13404 6276 13456
rect 6328 13444 6334 13456
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 6328 13416 6561 13444
rect 6328 13404 6334 13416
rect 6549 13413 6561 13416
rect 6595 13413 6607 13447
rect 6549 13407 6607 13413
rect 8202 13404 8208 13456
rect 8260 13444 8266 13456
rect 10410 13444 10416 13456
rect 8260 13416 10416 13444
rect 8260 13404 8266 13416
rect 6454 13376 6460 13388
rect 5920 13348 6460 13376
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 8386 13336 8392 13388
rect 8444 13376 8450 13388
rect 8444 13348 9168 13376
rect 8444 13336 8450 13348
rect 4157 13311 4215 13317
rect 3292 13280 4108 13308
rect 3292 13268 3298 13280
rect 2774 13200 2780 13252
rect 2832 13240 2838 13252
rect 3510 13240 3516 13252
rect 2832 13212 3516 13240
rect 2832 13200 2838 13212
rect 3510 13200 3516 13212
rect 3568 13200 3574 13252
rect 3694 13200 3700 13252
rect 3752 13240 3758 13252
rect 3970 13240 3976 13252
rect 3752 13212 3976 13240
rect 3752 13200 3758 13212
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 4080 13240 4108 13280
rect 4157 13277 4169 13311
rect 4203 13277 4215 13311
rect 5905 13311 5963 13317
rect 5905 13308 5917 13311
rect 4157 13271 4215 13277
rect 4264 13280 5917 13308
rect 4264 13249 4292 13280
rect 5905 13277 5917 13280
rect 5951 13308 5963 13311
rect 6086 13308 6092 13320
rect 5951 13280 6092 13308
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 6181 13311 6239 13317
rect 6181 13277 6193 13311
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 4249 13243 4307 13249
rect 4249 13240 4261 13243
rect 4080 13212 4261 13240
rect 4249 13209 4261 13212
rect 4295 13209 4307 13243
rect 4249 13203 4307 13209
rect 4706 13200 4712 13252
rect 4764 13240 4770 13252
rect 6196 13240 6224 13271
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 6730 13308 6736 13320
rect 6420 13280 6736 13308
rect 6420 13268 6426 13280
rect 6730 13268 6736 13280
rect 6788 13268 6794 13320
rect 8294 13268 8300 13320
rect 8352 13268 8358 13320
rect 8478 13268 8484 13320
rect 8536 13268 8542 13320
rect 8570 13268 8576 13320
rect 8628 13268 8634 13320
rect 9140 13317 9168 13348
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 9309 13379 9367 13385
rect 9309 13376 9321 13379
rect 9272 13348 9321 13376
rect 9272 13336 9278 13348
rect 9309 13345 9321 13348
rect 9355 13345 9367 13379
rect 9309 13339 9367 13345
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 8956 13240 8984 13271
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 9876 13317 9904 13416
rect 10410 13404 10416 13416
rect 10468 13404 10474 13456
rect 11072 13416 13584 13444
rect 11072 13385 11100 13416
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 11057 13379 11115 13385
rect 10183 13348 11008 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10042 13317 10048 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9640 13280 9689 13308
rect 9640 13268 9646 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9861 13311 9919 13317
rect 9861 13277 9873 13311
rect 9907 13277 9919 13311
rect 9861 13271 9919 13277
rect 9999 13311 10048 13317
rect 9999 13277 10011 13311
rect 10045 13277 10048 13311
rect 9999 13271 10048 13277
rect 10042 13268 10048 13271
rect 10100 13268 10106 13320
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 10980 13308 11008 13348
rect 11057 13345 11069 13379
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 13446 13376 13452 13388
rect 12492 13348 12664 13376
rect 12492 13336 12498 13348
rect 10980 13280 12020 13308
rect 9766 13240 9772 13252
rect 4764 13212 6224 13240
rect 8312 13212 8984 13240
rect 9140 13212 9772 13240
rect 4764 13200 4770 13212
rect 8312 13184 8340 13212
rect 9140 13184 9168 13212
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 5074 13132 5080 13184
rect 5132 13172 5138 13184
rect 5902 13172 5908 13184
rect 5132 13144 5908 13172
rect 5132 13132 5138 13144
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 8294 13132 8300 13184
rect 8352 13132 8358 13184
rect 9122 13132 9128 13184
rect 9180 13132 9186 13184
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 10870 13172 10876 13184
rect 9272 13144 10876 13172
rect 9272 13132 9278 13144
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11790 13132 11796 13184
rect 11848 13172 11854 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11848 13144 11897 13172
rect 11848 13132 11854 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 11992 13172 12020 13280
rect 12066 13268 12072 13320
rect 12124 13268 12130 13320
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 12636 13317 12664 13348
rect 12820 13348 13452 13376
rect 12820 13317 12848 13348
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 12308 13280 12357 13308
rect 12308 13268 12314 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 13262 13268 13268 13320
rect 13320 13308 13326 13320
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 13320 13280 13369 13308
rect 13320 13268 13326 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 12437 13243 12495 13249
rect 12437 13209 12449 13243
rect 12483 13209 12495 13243
rect 13556 13240 13584 13416
rect 13648 13385 13676 13484
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13771 13484 14105 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 15654 13444 15660 13456
rect 13872 13416 15660 13444
rect 13872 13404 13878 13416
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13345 13691 13379
rect 14430 13376 14458 13416
rect 15654 13404 15660 13416
rect 15712 13404 15718 13456
rect 16942 13376 16948 13388
rect 13633 13339 13691 13345
rect 14384 13348 14458 13376
rect 14752 13348 16948 13376
rect 14384 13317 14412 13348
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14458 13268 14464 13320
rect 14516 13268 14522 13320
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 14752 13317 14780 13348
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13308 16451 13311
rect 16482 13308 16488 13320
rect 16439 13280 16488 13308
rect 16439 13277 16451 13280
rect 16393 13271 16451 13277
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 15010 13240 15016 13252
rect 13556 13212 15016 13240
rect 12437 13203 12495 13209
rect 12158 13172 12164 13184
rect 11992 13144 12164 13172
rect 11885 13135 11943 13141
rect 12158 13132 12164 13144
rect 12216 13172 12222 13184
rect 12253 13175 12311 13181
rect 12253 13172 12265 13175
rect 12216 13144 12265 13172
rect 12216 13132 12222 13144
rect 12253 13141 12265 13144
rect 12299 13172 12311 13175
rect 12452 13172 12480 13203
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 12299 13144 12480 13172
rect 12299 13141 12311 13144
rect 12253 13135 12311 13141
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 13538 13172 13544 13184
rect 12768 13144 13544 13172
rect 12768 13132 12774 13144
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 13906 13132 13912 13184
rect 13964 13132 13970 13184
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 15286 13172 15292 13184
rect 14056 13144 15292 13172
rect 14056 13132 14062 13144
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 17681 13175 17739 13181
rect 17681 13172 17693 13175
rect 15896 13144 17693 13172
rect 15896 13132 15902 13144
rect 17681 13141 17693 13144
rect 17727 13141 17739 13175
rect 17681 13135 17739 13141
rect 1104 13082 18492 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 18492 13082
rect 1104 13008 18492 13030
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 5166 12968 5172 12980
rect 4672 12940 5172 12968
rect 4672 12928 4678 12940
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 6454 12928 6460 12980
rect 6512 12968 6518 12980
rect 6917 12971 6975 12977
rect 6917 12968 6929 12971
rect 6512 12940 6929 12968
rect 6512 12928 6518 12940
rect 6917 12937 6929 12940
rect 6963 12968 6975 12971
rect 8018 12968 8024 12980
rect 6963 12940 8024 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 8570 12928 8576 12980
rect 8628 12928 8634 12980
rect 9674 12968 9680 12980
rect 8864 12940 9680 12968
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 3237 12903 3295 12909
rect 3237 12900 3249 12903
rect 2924 12872 3249 12900
rect 2924 12860 2930 12872
rect 3237 12869 3249 12872
rect 3283 12900 3295 12903
rect 4706 12900 4712 12912
rect 3283 12872 4712 12900
rect 3283 12869 3295 12872
rect 3237 12863 3295 12869
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 5810 12900 5816 12912
rect 4908 12872 5816 12900
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3142 12832 3148 12844
rect 3099 12804 3148 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3326 12792 3332 12844
rect 3384 12792 3390 12844
rect 3602 12792 3608 12844
rect 3660 12832 3666 12844
rect 3786 12832 3792 12844
rect 3660 12804 3792 12832
rect 3660 12792 3666 12804
rect 3786 12792 3792 12804
rect 3844 12832 3850 12844
rect 4908 12841 4936 12872
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 4617 12835 4675 12841
rect 4617 12832 4629 12835
rect 3844 12804 4629 12832
rect 3844 12792 3850 12804
rect 4617 12801 4629 12804
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12801 5043 12835
rect 4985 12795 5043 12801
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 5994 12832 6000 12844
rect 5215 12804 6000 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 5000 12764 5028 12795
rect 5994 12792 6000 12804
rect 6052 12832 6058 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6052 12804 6561 12832
rect 6052 12792 6058 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 8202 12832 8208 12844
rect 7147 12804 8208 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12832 8447 12835
rect 8570 12832 8576 12844
rect 8435 12804 8576 12832
rect 8435 12801 8447 12804
rect 8389 12795 8447 12801
rect 5074 12764 5080 12776
rect 4571 12736 5080 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5074 12724 5080 12736
rect 5132 12764 5138 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 5132 12736 6653 12764
rect 5132 12724 5138 12736
rect 6641 12733 6653 12736
rect 6687 12764 6699 12767
rect 8404 12764 8432 12795
rect 8570 12792 8576 12804
rect 8628 12792 8634 12844
rect 8864 12841 8892 12940
rect 9674 12928 9680 12940
rect 9732 12968 9738 12980
rect 10042 12968 10048 12980
rect 9732 12940 10048 12968
rect 9732 12928 9738 12940
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 10928 12940 13860 12968
rect 10928 12928 10934 12940
rect 11054 12900 11060 12912
rect 8956 12872 11060 12900
rect 8956 12841 8984 12872
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 12342 12900 12348 12912
rect 12124 12872 12348 12900
rect 12124 12860 12130 12872
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 12805 12903 12863 12909
rect 12805 12869 12817 12903
rect 12851 12900 12863 12903
rect 13832 12900 13860 12940
rect 13906 12928 13912 12980
rect 13964 12928 13970 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 14884 12940 15792 12968
rect 14884 12928 14890 12940
rect 14274 12900 14280 12912
rect 12851 12872 13400 12900
rect 13832 12872 14280 12900
rect 12851 12869 12863 12872
rect 12805 12863 12863 12869
rect 8849 12835 8907 12841
rect 8849 12801 8861 12835
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9048 12764 9076 12795
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 9398 12764 9404 12776
rect 6687 12736 8432 12764
rect 8680 12736 9404 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 2958 12656 2964 12708
rect 3016 12696 3022 12708
rect 3053 12699 3111 12705
rect 3053 12696 3065 12699
rect 3016 12668 3065 12696
rect 3016 12656 3022 12668
rect 3053 12665 3065 12668
rect 3099 12665 3111 12699
rect 3053 12659 3111 12665
rect 3160 12668 7420 12696
rect 3160 12640 3188 12668
rect 3142 12588 3148 12640
rect 3200 12588 3206 12640
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 4614 12628 4620 12640
rect 4120 12600 4620 12628
rect 4120 12588 4126 12600
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5166 12588 5172 12640
rect 5224 12588 5230 12640
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6144 12600 6561 12628
rect 6144 12588 6150 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 7285 12631 7343 12637
rect 7285 12628 7297 12631
rect 7248 12600 7297 12628
rect 7248 12588 7254 12600
rect 7285 12597 7297 12600
rect 7331 12597 7343 12631
rect 7392 12628 7420 12668
rect 8294 12656 8300 12708
rect 8352 12656 8358 12708
rect 8386 12656 8392 12708
rect 8444 12696 8450 12708
rect 8680 12696 8708 12736
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 10612 12764 10640 12795
rect 10778 12792 10784 12844
rect 10836 12792 10842 12844
rect 10870 12792 10876 12844
rect 10928 12792 10934 12844
rect 12710 12792 12716 12844
rect 12768 12792 12774 12844
rect 12894 12792 12900 12844
rect 12952 12792 12958 12844
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 13004 12804 13185 12832
rect 11330 12764 11336 12776
rect 10612 12736 11336 12764
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 13004 12764 13032 12804
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 13262 12792 13268 12844
rect 13320 12792 13326 12844
rect 13372 12841 13400 12872
rect 14274 12860 14280 12872
rect 14332 12860 14338 12912
rect 15102 12900 15108 12912
rect 14660 12872 15108 12900
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 13906 12832 13912 12844
rect 13771 12804 13912 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12832 14059 12835
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 14047 12804 14197 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 12584 12736 13032 12764
rect 12584 12724 12590 12736
rect 13078 12724 13084 12776
rect 13136 12724 13142 12776
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14384 12764 14412 12795
rect 14458 12792 14464 12844
rect 14516 12792 14522 12844
rect 14660 12841 14688 12872
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 15764 12909 15792 12940
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 16816 12940 17141 12968
rect 16816 12928 16822 12940
rect 17129 12937 17141 12940
rect 17175 12937 17187 12971
rect 17129 12931 17187 12937
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12869 15807 12903
rect 15749 12863 15807 12869
rect 17497 12903 17555 12909
rect 17497 12869 17509 12903
rect 17543 12900 17555 12903
rect 17678 12900 17684 12912
rect 17543 12872 17684 12900
rect 17543 12869 17555 12872
rect 17497 12863 17555 12869
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 14734 12792 14740 12844
rect 14792 12792 14798 12844
rect 15194 12792 15200 12844
rect 15252 12792 15258 12844
rect 16666 12792 16672 12844
rect 16724 12792 16730 12844
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16908 12804 16957 12832
rect 16908 12792 16914 12804
rect 16945 12801 16957 12804
rect 16991 12832 17003 12835
rect 17310 12832 17316 12844
rect 16991 12804 17316 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 14826 12764 14832 12776
rect 13872 12736 14832 12764
rect 13872 12724 13878 12736
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12733 15347 12767
rect 15289 12727 15347 12733
rect 8444 12668 8708 12696
rect 8444 12656 8450 12668
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 9858 12696 9864 12708
rect 8812 12668 9864 12696
rect 8812 12656 8818 12668
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 10410 12656 10416 12708
rect 10468 12656 10474 12708
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 12066 12696 12072 12708
rect 10836 12668 12072 12696
rect 10836 12656 10842 12668
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 13541 12699 13599 12705
rect 13541 12665 13553 12699
rect 13587 12696 13599 12699
rect 15304 12696 15332 12727
rect 15378 12724 15384 12776
rect 15436 12724 15442 12776
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 17880 12764 17908 12795
rect 15528 12736 17908 12764
rect 15528 12724 15534 12736
rect 13587 12668 15332 12696
rect 13587 12665 13599 12668
rect 13541 12659 13599 12665
rect 13725 12631 13783 12637
rect 13725 12628 13737 12631
rect 7392 12600 13737 12628
rect 7285 12591 7343 12597
rect 13725 12597 13737 12600
rect 13771 12597 13783 12631
rect 13725 12591 13783 12597
rect 14274 12588 14280 12640
rect 14332 12628 14338 12640
rect 14550 12628 14556 12640
rect 14332 12600 14556 12628
rect 14332 12588 14338 12600
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 14829 12631 14887 12637
rect 14829 12628 14841 12631
rect 14700 12600 14841 12628
rect 14700 12588 14706 12600
rect 14829 12597 14841 12600
rect 14875 12597 14887 12631
rect 14829 12591 14887 12597
rect 14918 12588 14924 12640
rect 14976 12628 14982 12640
rect 15841 12631 15899 12637
rect 15841 12628 15853 12631
rect 14976 12600 15853 12628
rect 14976 12588 14982 12600
rect 15841 12597 15853 12600
rect 15887 12597 15899 12631
rect 15841 12591 15899 12597
rect 16758 12588 16764 12640
rect 16816 12588 16822 12640
rect 18046 12588 18052 12640
rect 18104 12588 18110 12640
rect 1104 12538 18492 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 18492 12538
rect 1104 12464 18492 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2222 12424 2228 12436
rect 2004 12396 2228 12424
rect 2004 12384 2010 12396
rect 2222 12384 2228 12396
rect 2280 12424 2286 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2280 12396 2421 12424
rect 2280 12384 2286 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 2409 12387 2467 12393
rect 3326 12384 3332 12436
rect 3384 12424 3390 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3384 12396 3801 12424
rect 3384 12384 3390 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 5258 12424 5264 12436
rect 3789 12387 3847 12393
rect 3896 12396 5264 12424
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 3896 12356 3924 12396
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 7432 12396 7481 12424
rect 7432 12384 7438 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 7469 12387 7527 12393
rect 8113 12427 8171 12433
rect 8113 12393 8125 12427
rect 8159 12424 8171 12427
rect 9030 12424 9036 12436
rect 8159 12396 9036 12424
rect 8159 12393 8171 12396
rect 8113 12387 8171 12393
rect 9030 12384 9036 12396
rect 9088 12424 9094 12436
rect 10226 12424 10232 12436
rect 9088 12396 10232 12424
rect 9088 12384 9094 12396
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 10652 12396 10977 12424
rect 10652 12384 10658 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 12710 12424 12716 12436
rect 10965 12387 11023 12393
rect 11440 12396 12716 12424
rect 3292 12328 3924 12356
rect 3292 12316 3298 12328
rect 4338 12316 4344 12368
rect 4396 12316 4402 12368
rect 4430 12316 4436 12368
rect 4488 12356 4494 12368
rect 4617 12359 4675 12365
rect 4617 12356 4629 12359
rect 4488 12328 4629 12356
rect 4488 12316 4494 12328
rect 4617 12325 4629 12328
rect 4663 12325 4675 12359
rect 4617 12319 4675 12325
rect 4706 12316 4712 12368
rect 4764 12316 4770 12368
rect 4982 12316 4988 12368
rect 5040 12356 5046 12368
rect 6181 12359 6239 12365
rect 6181 12356 6193 12359
rect 5040 12328 6193 12356
rect 5040 12316 5046 12328
rect 6181 12325 6193 12328
rect 6227 12325 6239 12359
rect 7285 12359 7343 12365
rect 7285 12356 7297 12359
rect 6181 12319 6239 12325
rect 6656 12328 7297 12356
rect 2774 12288 2780 12300
rect 2148 12260 2780 12288
rect 2148 12229 2176 12260
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 4062 12288 4068 12300
rect 3988 12260 4068 12288
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2271 12223 2329 12229
rect 2271 12189 2283 12223
rect 2317 12189 2329 12223
rect 2271 12183 2329 12189
rect 2286 12152 2314 12183
rect 2590 12180 2596 12232
rect 2648 12220 2654 12232
rect 3326 12220 3332 12232
rect 2648 12192 3332 12220
rect 2648 12180 2654 12192
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 3988 12229 4016 12260
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4356 12288 4384 12316
rect 4172 12260 4384 12288
rect 4525 12291 4583 12297
rect 4172 12229 4200 12260
rect 4525 12257 4537 12291
rect 4571 12288 4583 12291
rect 4724 12288 4752 12316
rect 5534 12288 5540 12300
rect 4571 12260 4752 12288
rect 4908 12260 5540 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 4246 12180 4252 12232
rect 4304 12229 4310 12232
rect 4304 12223 4333 12229
rect 4321 12189 4333 12223
rect 4304 12183 4333 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4614 12220 4620 12232
rect 4479 12192 4620 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4304 12180 4310 12183
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 4908 12229 4936 12260
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 6656 12288 6684 12328
rect 7285 12325 7297 12328
rect 7331 12356 7343 12359
rect 8754 12356 8760 12368
rect 7331 12328 8760 12356
rect 7331 12325 7343 12328
rect 7285 12319 7343 12325
rect 8754 12316 8760 12328
rect 8812 12316 8818 12368
rect 11440 12356 11468 12396
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 14645 12427 14703 12433
rect 14645 12393 14657 12427
rect 14691 12424 14703 12427
rect 14691 12396 15056 12424
rect 14691 12393 14703 12396
rect 14645 12387 14703 12393
rect 9600 12328 11468 12356
rect 7190 12288 7196 12300
rect 6600 12260 6684 12288
rect 6840 12260 7196 12288
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 3878 12152 3884 12164
rect 2286 12124 3884 12152
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 4065 12155 4123 12161
rect 4065 12121 4077 12155
rect 4111 12152 4123 12155
rect 4522 12152 4528 12164
rect 4111 12124 4528 12152
rect 4111 12121 4123 12124
rect 4065 12115 4123 12121
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12084 2651 12087
rect 2682 12084 2688 12096
rect 2639 12056 2688 12084
rect 2639 12053 2651 12056
rect 2593 12047 2651 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 4724 12084 4752 12183
rect 4816 12152 4844 12183
rect 5074 12180 5080 12232
rect 5132 12180 5138 12232
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 5994 12220 6000 12232
rect 5776 12192 6000 12220
rect 5776 12180 5782 12192
rect 5994 12180 6000 12192
rect 6052 12220 6058 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 6052 12192 6377 12220
rect 6052 12180 6058 12192
rect 6365 12189 6377 12192
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 6454 12180 6460 12232
rect 6512 12180 6518 12232
rect 6600 12229 6628 12260
rect 6840 12229 6868 12260
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 7926 12248 7932 12300
rect 7984 12288 7990 12300
rect 7984 12260 8156 12288
rect 7984 12248 7990 12260
rect 8128 12229 8156 12260
rect 8938 12248 8944 12300
rect 8996 12288 9002 12300
rect 9033 12291 9091 12297
rect 9033 12288 9045 12291
rect 8996 12260 9045 12288
rect 8996 12248 9002 12260
rect 9033 12257 9045 12260
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 9122 12248 9128 12300
rect 9180 12248 9186 12300
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 9272 12260 9321 12288
rect 9272 12248 9278 12260
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9309 12251 9367 12257
rect 6585 12223 6643 12229
rect 6585 12189 6597 12223
rect 6631 12189 6643 12223
rect 6585 12183 6643 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 8386 12220 8392 12232
rect 8343 12192 8392 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 4816 12124 4997 12152
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 4985 12115 5043 12121
rect 6178 12112 6184 12164
rect 6236 12112 6242 12164
rect 6932 12152 6960 12183
rect 6380 12124 6960 12152
rect 6380 12096 6408 12124
rect 3476 12056 4752 12084
rect 3476 12044 3482 12056
rect 6362 12044 6368 12096
rect 6420 12044 6426 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 7020 12084 7048 12183
rect 7098 12112 7104 12164
rect 7156 12152 7162 12164
rect 7193 12155 7251 12161
rect 7193 12152 7205 12155
rect 7156 12124 7205 12152
rect 7156 12112 7162 12124
rect 7193 12121 7205 12124
rect 7239 12152 7251 12155
rect 7437 12155 7495 12161
rect 7437 12152 7449 12155
rect 7239 12124 7449 12152
rect 7239 12121 7251 12124
rect 7193 12115 7251 12121
rect 7437 12121 7449 12124
rect 7483 12121 7495 12155
rect 7437 12115 7495 12121
rect 7558 12112 7564 12164
rect 7616 12152 7622 12164
rect 7653 12155 7711 12161
rect 7653 12152 7665 12155
rect 7616 12124 7665 12152
rect 7616 12112 7622 12124
rect 7653 12121 7665 12124
rect 7699 12121 7711 12155
rect 7653 12115 7711 12121
rect 7742 12112 7748 12164
rect 7800 12152 7806 12164
rect 8036 12152 8064 12183
rect 8386 12180 8392 12192
rect 8444 12220 8450 12232
rect 8444 12192 9352 12220
rect 8444 12180 8450 12192
rect 8846 12152 8852 12164
rect 7800 12124 7973 12152
rect 8036 12124 8852 12152
rect 7800 12112 7806 12124
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 6788 12056 7849 12084
rect 6788 12044 6794 12056
rect 7837 12053 7849 12056
rect 7883 12053 7895 12087
rect 7945 12084 7973 12124
rect 8846 12112 8852 12124
rect 8904 12112 8910 12164
rect 8938 12112 8944 12164
rect 8996 12112 9002 12164
rect 9324 12152 9352 12192
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 9513 12223 9571 12229
rect 9513 12220 9525 12223
rect 9508 12189 9525 12220
rect 9559 12189 9571 12223
rect 9508 12183 9571 12189
rect 9508 12152 9536 12183
rect 9324 12124 9536 12152
rect 9600 12084 9628 12328
rect 11054 12248 11060 12300
rect 11112 12296 11118 12300
rect 11440 12297 11468 12328
rect 11977 12359 12035 12365
rect 11977 12325 11989 12359
rect 12023 12356 12035 12359
rect 12158 12356 12164 12368
rect 12023 12328 12164 12356
rect 12023 12325 12035 12328
rect 11977 12319 12035 12325
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 12250 12316 12256 12368
rect 12308 12316 12314 12368
rect 14918 12356 14924 12368
rect 14844 12328 14924 12356
rect 11112 12288 11238 12296
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 11112 12268 11345 12288
rect 11112 12248 11118 12268
rect 11210 12260 11345 12268
rect 11333 12257 11345 12260
rect 11379 12257 11391 12291
rect 11333 12251 11391 12257
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 11425 12251 11483 12257
rect 11624 12260 11805 12288
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 9674 12112 9680 12164
rect 9732 12112 9738 12164
rect 9876 12096 9904 12183
rect 10226 12180 10232 12232
rect 10284 12180 10290 12232
rect 11146 12180 11152 12232
rect 11204 12180 11210 12232
rect 11514 12180 11520 12232
rect 11572 12180 11578 12232
rect 10244 12152 10272 12180
rect 11624 12152 11652 12260
rect 11793 12257 11805 12260
rect 11839 12257 11851 12291
rect 11793 12251 11851 12257
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 11940 12260 12204 12288
rect 11940 12248 11946 12260
rect 12176 12232 12204 12260
rect 11698 12180 11704 12232
rect 11756 12180 11762 12232
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 12069 12223 12127 12229
rect 12069 12220 12081 12223
rect 12032 12192 12081 12220
rect 12032 12180 12038 12192
rect 12069 12189 12081 12192
rect 12115 12189 12127 12223
rect 12069 12183 12127 12189
rect 12158 12180 12164 12232
rect 12216 12180 12222 12232
rect 12268 12220 12296 12316
rect 13170 12288 13176 12300
rect 12912 12260 13176 12288
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 12268 12192 12357 12220
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 12434 12180 12440 12232
rect 12492 12180 12498 12232
rect 12912 12229 12940 12260
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 14844 12288 14872 12328
rect 14918 12316 14924 12328
rect 14976 12316 14982 12368
rect 15028 12356 15056 12396
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 15252 12396 15577 12424
rect 15252 12384 15258 12396
rect 15565 12393 15577 12396
rect 15611 12393 15623 12427
rect 15565 12387 15623 12393
rect 15470 12356 15476 12368
rect 15028 12328 15476 12356
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 14148 12260 14872 12288
rect 14148 12248 14154 12260
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 14369 12223 14427 12229
rect 14369 12220 14381 12223
rect 13127 12192 14381 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 14369 12189 14381 12192
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 14642 12180 14648 12232
rect 14700 12180 14706 12232
rect 14844 12229 14872 12260
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 15068 12260 15976 12288
rect 15068 12248 15074 12260
rect 15948 12232 15976 12260
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 16724 12260 17908 12288
rect 16724 12248 16730 12260
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 14918 12180 14924 12232
rect 14976 12180 14982 12232
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 15160 12192 15301 12220
rect 15160 12180 15166 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 15378 12180 15384 12232
rect 15436 12180 15442 12232
rect 15930 12180 15936 12232
rect 15988 12180 15994 12232
rect 16022 12180 16028 12232
rect 16080 12180 16086 12232
rect 17880 12229 17908 12260
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 10244 12124 11652 12152
rect 11793 12155 11851 12161
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 11882 12152 11888 12164
rect 11839 12124 11888 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 12575 12155 12633 12161
rect 12575 12152 12587 12155
rect 11992 12124 12587 12152
rect 11992 12096 12020 12124
rect 12575 12121 12587 12124
rect 12621 12121 12633 12155
rect 12575 12115 12633 12121
rect 12710 12112 12716 12164
rect 12768 12112 12774 12164
rect 12805 12155 12863 12161
rect 12805 12121 12817 12155
rect 12851 12152 12863 12155
rect 12986 12152 12992 12164
rect 12851 12124 12992 12152
rect 12851 12121 12863 12124
rect 12805 12115 12863 12121
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 15013 12155 15071 12161
rect 15013 12152 15025 12155
rect 14240 12124 15025 12152
rect 14240 12112 14246 12124
rect 15013 12121 15025 12124
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 15838 12112 15844 12164
rect 15896 12152 15902 12164
rect 16301 12155 16359 12161
rect 16301 12152 16313 12155
rect 15896 12124 16313 12152
rect 15896 12112 15902 12124
rect 16301 12121 16313 12124
rect 16347 12121 16359 12155
rect 16301 12115 16359 12121
rect 16758 12112 16764 12164
rect 16816 12112 16822 12164
rect 7945 12056 9628 12084
rect 7837 12047 7895 12053
rect 9858 12044 9864 12096
rect 9916 12044 9922 12096
rect 10045 12087 10103 12093
rect 10045 12053 10057 12087
rect 10091 12084 10103 12087
rect 10226 12084 10232 12096
rect 10091 12056 10232 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 11974 12044 11980 12096
rect 12032 12044 12038 12096
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 14918 12084 14924 12096
rect 12391 12056 14924 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15194 12044 15200 12096
rect 15252 12084 15258 12096
rect 15749 12087 15807 12093
rect 15749 12084 15761 12087
rect 15252 12056 15761 12084
rect 15252 12044 15258 12056
rect 15749 12053 15761 12056
rect 15795 12053 15807 12087
rect 15749 12047 15807 12053
rect 17770 12044 17776 12096
rect 17828 12044 17834 12096
rect 17954 12044 17960 12096
rect 18012 12044 18018 12096
rect 1104 11994 18492 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 18492 11994
rect 1104 11920 18492 11942
rect 1949 11883 2007 11889
rect 1949 11849 1961 11883
rect 1995 11880 2007 11883
rect 2317 11883 2375 11889
rect 2317 11880 2329 11883
rect 1995 11852 2329 11880
rect 1995 11849 2007 11852
rect 1949 11843 2007 11849
rect 2317 11849 2329 11852
rect 2363 11849 2375 11883
rect 2317 11843 2375 11849
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 4065 11883 4123 11889
rect 4065 11880 4077 11883
rect 2464 11852 4077 11880
rect 2464 11840 2470 11852
rect 1854 11704 1860 11756
rect 1912 11704 1918 11756
rect 2516 11753 2544 11852
rect 4065 11849 4077 11852
rect 4111 11849 4123 11883
rect 5537 11883 5595 11889
rect 5537 11880 5549 11883
rect 4065 11843 4123 11849
rect 4172 11852 5549 11880
rect 2682 11772 2688 11824
rect 2740 11772 2746 11824
rect 3326 11772 3332 11824
rect 3384 11812 3390 11824
rect 4172 11812 4200 11852
rect 5537 11849 5549 11852
rect 5583 11849 5595 11883
rect 5902 11880 5908 11892
rect 5537 11843 5595 11849
rect 5644 11852 5908 11880
rect 3384 11784 4200 11812
rect 3384 11772 3390 11784
rect 4338 11772 4344 11824
rect 4396 11812 4402 11824
rect 5644 11812 5672 11852
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6454 11880 6460 11892
rect 6328 11852 6460 11880
rect 6328 11840 6334 11852
rect 6454 11840 6460 11852
rect 6512 11880 6518 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6512 11852 6561 11880
rect 6512 11840 6518 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 7558 11880 7564 11892
rect 6549 11843 6607 11849
rect 6656 11852 7564 11880
rect 6656 11812 6684 11852
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 8110 11880 8116 11892
rect 7708 11852 8116 11880
rect 7708 11840 7714 11852
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9769 11883 9827 11889
rect 9769 11880 9781 11883
rect 9732 11852 9781 11880
rect 9732 11840 9738 11852
rect 9769 11849 9781 11852
rect 9815 11849 9827 11883
rect 9769 11843 9827 11849
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 9916 11852 10180 11880
rect 9916 11840 9922 11852
rect 8386 11812 8392 11824
rect 4396 11784 5395 11812
rect 4396 11772 4402 11784
rect 2496 11747 2554 11753
rect 2496 11713 2508 11747
rect 2542 11713 2554 11747
rect 2496 11707 2554 11713
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11713 2651 11747
rect 2593 11707 2651 11713
rect 1762 11636 1768 11688
rect 1820 11676 1826 11688
rect 2041 11679 2099 11685
rect 2041 11676 2053 11679
rect 1820 11648 2053 11676
rect 1820 11636 1826 11648
rect 2041 11645 2053 11648
rect 2087 11645 2099 11679
rect 2608 11676 2636 11707
rect 2774 11704 2780 11756
rect 2832 11753 2838 11756
rect 2832 11747 2871 11753
rect 2859 11713 2871 11747
rect 2832 11707 2871 11713
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11744 3019 11747
rect 3142 11744 3148 11756
rect 3007 11716 3148 11744
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 2832 11704 2838 11707
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4430 11744 4436 11756
rect 4295 11716 4436 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 4614 11744 4620 11756
rect 4571 11716 4620 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 4980 11747 5038 11753
rect 4980 11713 4992 11747
rect 5026 11713 5038 11747
rect 4980 11707 5038 11713
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 4798 11676 4804 11688
rect 2608 11648 2912 11676
rect 2041 11639 2099 11645
rect 2884 11620 2912 11648
rect 4448 11648 4804 11676
rect 2866 11568 2872 11620
rect 2924 11568 2930 11620
rect 4448 11617 4476 11648
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 4433 11611 4491 11617
rect 4433 11577 4445 11611
rect 4479 11577 4491 11611
rect 4433 11571 4491 11577
rect 1489 11543 1547 11549
rect 1489 11509 1501 11543
rect 1535 11540 1547 11543
rect 1670 11540 1676 11552
rect 1535 11512 1676 11540
rect 1535 11509 1547 11512
rect 1489 11503 1547 11509
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4764 11512 4813 11540
rect 4764 11500 4770 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 4995 11540 5023 11707
rect 5092 11608 5120 11707
rect 5166 11704 5172 11756
rect 5224 11704 5230 11756
rect 5367 11753 5395 11784
rect 5460 11784 5672 11812
rect 5736 11784 6684 11812
rect 6932 11784 8392 11812
rect 5460 11753 5488 11784
rect 5736 11753 5764 11784
rect 6288 11756 6316 11784
rect 5352 11747 5410 11753
rect 5352 11713 5364 11747
rect 5398 11713 5410 11747
rect 5352 11707 5410 11713
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 5367 11676 5395 11707
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 5994 11704 6000 11756
rect 6052 11704 6058 11756
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 6328 11716 6377 11744
rect 6328 11704 6334 11716
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6638 11704 6644 11756
rect 6696 11704 6702 11756
rect 6932 11753 6960 11784
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 7098 11704 7104 11756
rect 7156 11704 7162 11756
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 9858 11744 9864 11756
rect 7377 11707 7435 11713
rect 8266 11716 9864 11744
rect 6546 11676 6552 11688
rect 5367 11648 6552 11676
rect 6546 11636 6552 11648
rect 6604 11636 6610 11688
rect 7392 11676 7420 11707
rect 6932 11648 7420 11676
rect 6932 11620 6960 11648
rect 7558 11636 7564 11688
rect 7616 11676 7622 11688
rect 8266 11676 8294 11716
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 9950 11704 9956 11756
rect 10008 11704 10014 11756
rect 10042 11704 10048 11756
rect 10100 11704 10106 11756
rect 10152 11753 10180 11852
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11422 11880 11428 11892
rect 11296 11852 11428 11880
rect 11296 11840 11302 11852
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11572 11852 11805 11880
rect 11572 11840 11578 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 12710 11840 12716 11892
rect 12768 11840 12774 11892
rect 14182 11880 14188 11892
rect 13004 11852 14188 11880
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 11756 11784 12848 11812
rect 11756 11772 11762 11784
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11744 10195 11747
rect 11517 11747 11575 11753
rect 10183 11716 11376 11744
rect 10183 11713 10195 11716
rect 10137 11707 10195 11713
rect 10229 11679 10287 11685
rect 7616 11648 8294 11676
rect 9646 11648 10088 11676
rect 7616 11636 7622 11648
rect 5810 11608 5816 11620
rect 5092 11580 5816 11608
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 6178 11568 6184 11620
rect 6236 11608 6242 11620
rect 6365 11611 6423 11617
rect 6365 11608 6377 11611
rect 6236 11580 6377 11608
rect 6236 11568 6242 11580
rect 6365 11577 6377 11580
rect 6411 11577 6423 11611
rect 6365 11571 6423 11577
rect 6914 11568 6920 11620
rect 6972 11568 6978 11620
rect 7193 11611 7251 11617
rect 7193 11577 7205 11611
rect 7239 11577 7251 11611
rect 7193 11571 7251 11577
rect 7285 11611 7343 11617
rect 7285 11577 7297 11611
rect 7331 11608 7343 11611
rect 7926 11608 7932 11620
rect 7331 11580 7932 11608
rect 7331 11577 7343 11580
rect 7285 11571 7343 11577
rect 5350 11540 5356 11552
rect 4995 11512 5356 11540
rect 4801 11503 4859 11509
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 7208 11540 7236 11571
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 9646 11608 9674 11648
rect 8266 11580 9674 11608
rect 7466 11540 7472 11552
rect 7208 11512 7472 11540
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 7561 11543 7619 11549
rect 7561 11509 7573 11543
rect 7607 11540 7619 11543
rect 8266 11540 8294 11580
rect 7607 11512 8294 11540
rect 10060 11540 10088 11648
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 11146 11676 11152 11688
rect 10275 11648 11152 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11348 11608 11376 11716
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 11882 11744 11888 11756
rect 11563 11716 11888 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 12820 11753 12848 11784
rect 12805 11748 12863 11753
rect 12805 11747 12880 11748
rect 12805 11713 12817 11747
rect 12851 11744 12880 11747
rect 13004 11744 13032 11852
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 15381 11883 15439 11889
rect 15381 11849 15393 11883
rect 15427 11880 15439 11883
rect 15562 11880 15568 11892
rect 15427 11852 15568 11880
rect 15427 11849 15439 11852
rect 15381 11843 15439 11849
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 15838 11840 15844 11892
rect 15896 11840 15902 11892
rect 13446 11812 13452 11824
rect 13188 11784 13452 11812
rect 13188 11753 13216 11784
rect 13446 11772 13452 11784
rect 13504 11812 13510 11824
rect 15194 11812 15200 11824
rect 13504 11784 15200 11812
rect 13504 11772 13510 11784
rect 15194 11772 15200 11784
rect 15252 11772 15258 11824
rect 15930 11772 15936 11824
rect 15988 11812 15994 11824
rect 15988 11784 16712 11812
rect 15988 11772 15994 11784
rect 12851 11716 13032 11744
rect 13173 11747 13231 11753
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13262 11704 13268 11756
rect 13320 11704 13326 11756
rect 13354 11704 13360 11756
rect 13412 11704 13418 11756
rect 13538 11704 13544 11756
rect 13596 11704 13602 11756
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11744 15531 11747
rect 16114 11744 16120 11756
rect 15519 11716 16120 11744
rect 15519 11713 15531 11716
rect 15473 11707 15531 11713
rect 16114 11704 16120 11716
rect 16172 11744 16178 11756
rect 16684 11753 16712 11784
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 16172 11716 16221 11744
rect 16172 11704 16178 11716
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11744 16727 11747
rect 16715 11716 17540 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11676 11667 11679
rect 11698 11676 11704 11688
rect 11655 11648 11704 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11676 12955 11679
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 12943 11648 13737 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 11808 11608 11836 11639
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 14884 11648 15792 11676
rect 14884 11636 14890 11648
rect 12158 11608 12164 11620
rect 11348 11580 11652 11608
rect 11808 11580 12164 11608
rect 11514 11540 11520 11552
rect 10060 11512 11520 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 11624 11540 11652 11580
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 13354 11608 13360 11620
rect 12268 11580 13360 11608
rect 12268 11540 12296 11580
rect 13354 11568 13360 11580
rect 13412 11568 13418 11620
rect 15102 11568 15108 11620
rect 15160 11608 15166 11620
rect 15197 11611 15255 11617
rect 15197 11608 15209 11611
rect 15160 11580 15209 11608
rect 15160 11568 15166 11580
rect 15197 11577 15209 11580
rect 15243 11577 15255 11611
rect 15764 11608 15792 11648
rect 15838 11636 15844 11688
rect 15896 11636 15902 11688
rect 15930 11636 15936 11688
rect 15988 11636 15994 11688
rect 17512 11685 17540 11716
rect 17770 11704 17776 11756
rect 17828 11704 17834 11756
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 16942 11608 16948 11620
rect 15764 11580 16948 11608
rect 15197 11571 15255 11577
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 17512 11608 17540 11639
rect 17770 11608 17776 11620
rect 17512 11580 17776 11608
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 11624 11512 12296 11540
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 13081 11543 13139 11549
rect 13081 11540 13093 11543
rect 12584 11512 13093 11540
rect 12584 11500 12590 11512
rect 13081 11509 13093 11512
rect 13127 11540 13139 11543
rect 13722 11540 13728 11552
rect 13127 11512 13728 11540
rect 13127 11509 13139 11512
rect 13081 11503 13139 11509
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 16117 11543 16175 11549
rect 16117 11509 16129 11543
rect 16163 11540 16175 11543
rect 16758 11540 16764 11552
rect 16163 11512 16764 11540
rect 16163 11509 16175 11512
rect 16117 11503 16175 11509
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 16850 11500 16856 11552
rect 16908 11500 16914 11552
rect 1104 11450 18492 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 18492 11450
rect 1104 11376 18492 11398
rect 1118 11296 1124 11348
rect 1176 11336 1182 11348
rect 1489 11339 1547 11345
rect 1489 11336 1501 11339
rect 1176 11308 1501 11336
rect 1176 11296 1182 11308
rect 1489 11305 1501 11308
rect 1535 11305 1547 11339
rect 1489 11299 1547 11305
rect 1854 11296 1860 11348
rect 1912 11336 1918 11348
rect 1949 11339 2007 11345
rect 1949 11336 1961 11339
rect 1912 11308 1961 11336
rect 1912 11296 1918 11308
rect 1949 11305 1961 11308
rect 1995 11305 2007 11339
rect 1949 11299 2007 11305
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 3142 11336 3148 11348
rect 2179 11308 3148 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 3936 11308 4261 11336
rect 3936 11296 3942 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 4249 11299 4307 11305
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 4614 11336 4620 11348
rect 4479 11308 4620 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 2777 11271 2835 11277
rect 2777 11268 2789 11271
rect 2056 11240 2789 11268
rect 2056 11209 2084 11240
rect 2777 11237 2789 11240
rect 2823 11237 2835 11271
rect 2777 11231 2835 11237
rect 3786 11228 3792 11280
rect 3844 11268 3850 11280
rect 4065 11271 4123 11277
rect 4065 11268 4077 11271
rect 3844 11240 4077 11268
rect 3844 11228 3850 11240
rect 4065 11237 4077 11240
rect 4111 11237 4123 11271
rect 4264 11268 4292 11299
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 5350 11296 5356 11348
rect 5408 11336 5414 11348
rect 5408 11308 7144 11336
rect 5408 11296 5414 11308
rect 4264 11240 6959 11268
rect 4065 11231 4123 11237
rect 6931 11212 6959 11240
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11169 2099 11203
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 2041 11163 2099 11169
rect 3804 11172 4629 11200
rect 3804 11144 3832 11172
rect 4617 11169 4629 11172
rect 4663 11200 4675 11203
rect 4663 11172 6408 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 1670 11092 1676 11144
rect 1728 11092 1734 11144
rect 2314 11092 2320 11144
rect 2372 11132 2378 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 2372 11104 2513 11132
rect 2372 11092 2378 11104
rect 2501 11101 2513 11104
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 2590 11092 2596 11144
rect 2648 11092 2654 11144
rect 3786 11092 3792 11144
rect 3844 11092 3850 11144
rect 4430 11092 4436 11144
rect 4488 11092 4494 11144
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 6270 11132 6276 11144
rect 4847 11104 6276 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 2406 11024 2412 11076
rect 2464 11024 2470 11076
rect 2682 11024 2688 11076
rect 2740 11064 2746 11076
rect 2777 11067 2835 11073
rect 2777 11064 2789 11067
rect 2740 11036 2789 11064
rect 2740 11024 2746 11036
rect 2777 11033 2789 11036
rect 2823 11033 2835 11067
rect 2777 11027 2835 11033
rect 3234 11024 3240 11076
rect 3292 11064 3298 11076
rect 4709 11067 4767 11073
rect 4709 11064 4721 11067
rect 3292 11036 4721 11064
rect 3292 11024 3298 11036
rect 4709 11033 4721 11036
rect 4755 11064 4767 11067
rect 4982 11064 4988 11076
rect 4755 11036 4988 11064
rect 4755 11033 4767 11036
rect 4709 11027 4767 11033
rect 4982 11024 4988 11036
rect 5040 11024 5046 11076
rect 6380 11064 6408 11172
rect 6914 11160 6920 11212
rect 6972 11160 6978 11212
rect 7116 11200 7144 11308
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7616 11308 7757 11336
rect 7616 11296 7622 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 7926 11296 7932 11348
rect 7984 11296 7990 11348
rect 9306 11336 9312 11348
rect 8864 11308 9312 11336
rect 7374 11228 7380 11280
rect 7432 11228 7438 11280
rect 8386 11228 8392 11280
rect 8444 11268 8450 11280
rect 8444 11240 8800 11268
rect 8444 11228 8450 11240
rect 7116 11172 7696 11200
rect 7116 11141 7144 11172
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 7190 11092 7196 11144
rect 7248 11132 7254 11144
rect 7248 11104 7604 11132
rect 7248 11092 7254 11104
rect 7208 11064 7236 11092
rect 6380 11036 7236 11064
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 7576 11073 7604 11104
rect 7469 11067 7527 11073
rect 7469 11064 7481 11067
rect 7340 11036 7481 11064
rect 7340 11024 7346 11036
rect 7469 11033 7481 11036
rect 7515 11033 7527 11067
rect 7469 11027 7527 11033
rect 7561 11067 7619 11073
rect 7561 11033 7573 11067
rect 7607 11033 7619 11067
rect 7668 11064 7696 11172
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8202 11132 8208 11144
rect 8159 11104 8208 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 8294 11092 8300 11144
rect 8352 11092 8358 11144
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 7668 11036 8156 11064
rect 7561 11027 7619 11033
rect 8128 11008 8156 11036
rect 2317 10999 2375 11005
rect 2317 10965 2329 10999
rect 2363 10996 2375 10999
rect 2866 10996 2872 11008
rect 2363 10968 2872 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 3878 10956 3884 11008
rect 3936 10996 3942 11008
rect 5166 10996 5172 11008
rect 3936 10968 5172 10996
rect 3936 10956 3942 10968
rect 5166 10956 5172 10968
rect 5224 10996 5230 11008
rect 6362 10996 6368 11008
rect 5224 10968 6368 10996
rect 5224 10956 5230 10968
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7761 10999 7819 11005
rect 7761 10996 7773 10999
rect 6972 10968 7773 10996
rect 6972 10956 6978 10968
rect 7761 10965 7773 10968
rect 7807 10965 7819 10999
rect 7761 10959 7819 10965
rect 8110 10956 8116 11008
rect 8168 10956 8174 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8496 10996 8524 11095
rect 8570 11092 8576 11144
rect 8628 11092 8634 11144
rect 8772 11064 8800 11240
rect 8864 11144 8892 11308
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 12066 11336 12072 11348
rect 11756 11308 12072 11336
rect 11756 11296 11762 11308
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 13449 11339 13507 11345
rect 13449 11336 13461 11339
rect 12492 11308 13461 11336
rect 12492 11296 12498 11308
rect 13449 11305 13461 11308
rect 13495 11305 13507 11339
rect 13449 11299 13507 11305
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 15838 11336 15844 11348
rect 14516 11308 15844 11336
rect 14516 11296 14522 11308
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 17218 11336 17224 11348
rect 16540 11308 17224 11336
rect 16540 11296 16546 11308
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 9033 11271 9091 11277
rect 9033 11237 9045 11271
rect 9079 11268 9091 11271
rect 9214 11268 9220 11280
rect 9079 11240 9220 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 14553 11271 14611 11277
rect 14553 11268 14565 11271
rect 11572 11240 14565 11268
rect 11572 11228 11578 11240
rect 14553 11237 14565 11240
rect 14599 11237 14611 11271
rect 14553 11231 14611 11237
rect 15013 11271 15071 11277
rect 15013 11237 15025 11271
rect 15059 11237 15071 11271
rect 16500 11268 16528 11296
rect 15013 11231 15071 11237
rect 15948 11240 16528 11268
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11200 9183 11203
rect 9490 11200 9496 11212
rect 9171 11172 9496 11200
rect 9171 11169 9183 11172
rect 9125 11163 9183 11169
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8904 11104 8953 11132
rect 8904 11092 8910 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 9140 11132 9168 11163
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 11974 11200 11980 11212
rect 10192 11172 11980 11200
rect 10192 11160 10198 11172
rect 8941 11095 8999 11101
rect 9048 11104 9168 11132
rect 9401 11135 9459 11141
rect 9048 11064 9076 11104
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 9582 11132 9588 11144
rect 9447 11104 9588 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10045 11135 10103 11141
rect 10045 11132 10057 11135
rect 9732 11104 10057 11132
rect 9732 11092 9738 11104
rect 10045 11101 10057 11104
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10226 11092 10232 11144
rect 10284 11092 10290 11144
rect 10336 11141 10364 11172
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12802 11200 12808 11212
rect 12492 11172 12808 11200
rect 12492 11160 12498 11172
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 13078 11160 13084 11212
rect 13136 11160 13142 11212
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11200 13231 11203
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 13219 11172 13645 11200
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 14645 11203 14703 11209
rect 13633 11163 13691 11169
rect 13740 11172 14504 11200
rect 13740 11144 13768 11172
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 10502 11092 10508 11144
rect 10560 11092 10566 11144
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 12710 11132 12716 11144
rect 10928 11104 12716 11132
rect 10928 11092 10934 11104
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 13004 11064 13032 11095
rect 8772 11036 9076 11064
rect 9140 11036 13032 11064
rect 13280 11064 13308 11095
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13504 11104 13553 11132
rect 13504 11092 13510 11104
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 13722 11092 13728 11144
rect 13780 11092 13786 11144
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14366 11132 14372 11144
rect 14240 11104 14372 11132
rect 14240 11092 14246 11104
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 14476 11132 14504 11172
rect 14645 11169 14657 11203
rect 14691 11200 14703 11203
rect 15028 11200 15056 11231
rect 14691 11172 15056 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 14476 11104 14749 11132
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11132 15071 11135
rect 15378 11132 15384 11144
rect 15059 11104 15384 11132
rect 15059 11101 15071 11104
rect 15013 11095 15071 11101
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11132 15531 11135
rect 15948 11132 15976 11240
rect 16022 11160 16028 11212
rect 16080 11200 16086 11212
rect 16393 11203 16451 11209
rect 16393 11200 16405 11203
rect 16080 11172 16405 11200
rect 16080 11160 16086 11172
rect 16393 11169 16405 11172
rect 16439 11169 16451 11203
rect 16393 11163 16451 11169
rect 18138 11160 18144 11212
rect 18196 11160 18202 11212
rect 15519 11104 15976 11132
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16298 11132 16304 11144
rect 16172 11104 16304 11132
rect 16172 11092 16178 11104
rect 16298 11092 16304 11104
rect 16356 11092 16362 11144
rect 17954 11132 17960 11144
rect 17802 11104 17960 11132
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 14642 11064 14648 11076
rect 13280 11036 14648 11064
rect 8352 10968 8524 10996
rect 8757 10999 8815 11005
rect 8352 10956 8358 10968
rect 8757 10965 8769 10999
rect 8803 10996 8815 10999
rect 9140 10996 9168 11036
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 15562 11024 15568 11076
rect 15620 11064 15626 11076
rect 15620 11036 16528 11064
rect 15620 11024 15626 11036
rect 8803 10968 9168 10996
rect 8803 10965 8815 10968
rect 8757 10959 8815 10965
rect 9214 10956 9220 11008
rect 9272 10956 9278 11008
rect 9309 10999 9367 11005
rect 9309 10965 9321 10999
rect 9355 10996 9367 10999
rect 9766 10996 9772 11008
rect 9355 10968 9772 10996
rect 9355 10965 9367 10968
rect 9309 10959 9367 10965
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 11790 10996 11796 11008
rect 9916 10968 11796 10996
rect 9916 10956 9922 10968
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 14090 10956 14096 11008
rect 14148 10996 14154 11008
rect 14185 10999 14243 11005
rect 14185 10996 14197 10999
rect 14148 10968 14197 10996
rect 14148 10956 14154 10968
rect 14185 10965 14197 10968
rect 14231 10965 14243 10999
rect 14185 10959 14243 10965
rect 15654 10956 15660 11008
rect 15712 10956 15718 11008
rect 16117 10999 16175 11005
rect 16117 10965 16129 10999
rect 16163 10996 16175 10999
rect 16206 10996 16212 11008
rect 16163 10968 16212 10996
rect 16163 10965 16175 10968
rect 16117 10959 16175 10965
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 16500 10996 16528 11036
rect 16666 11024 16672 11076
rect 16724 11024 16730 11076
rect 17402 10996 17408 11008
rect 16500 10968 17408 10996
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 1104 10906 18492 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 18492 10906
rect 1104 10832 18492 10854
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 2406 10792 2412 10804
rect 2188 10764 2412 10792
rect 2188 10752 2194 10764
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 3694 10752 3700 10804
rect 3752 10752 3758 10804
rect 4062 10752 4068 10804
rect 4120 10752 4126 10804
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 4893 10795 4951 10801
rect 4893 10792 4905 10795
rect 4672 10764 4905 10792
rect 4672 10752 4678 10764
rect 4893 10761 4905 10764
rect 4939 10761 4951 10795
rect 4893 10755 4951 10761
rect 5353 10795 5411 10801
rect 5353 10761 5365 10795
rect 5399 10792 5411 10795
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5399 10764 5641 10792
rect 5399 10761 5411 10764
rect 5353 10755 5411 10761
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 7742 10792 7748 10804
rect 5868 10764 7748 10792
rect 5868 10752 5874 10764
rect 7742 10752 7748 10764
rect 7800 10792 7806 10804
rect 7800 10764 8028 10792
rect 7800 10752 7806 10764
rect 4080 10724 4108 10752
rect 4798 10724 4804 10736
rect 4080 10696 4804 10724
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 5166 10684 5172 10736
rect 5224 10724 5230 10736
rect 5224 10696 5580 10724
rect 5224 10684 5230 10696
rect 3513 10659 3571 10665
rect 3513 10625 3525 10659
rect 3559 10656 3571 10659
rect 3694 10656 3700 10668
rect 3559 10628 3700 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 3844 10628 3893 10656
rect 3844 10616 3850 10628
rect 3881 10625 3893 10628
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 3970 10616 3976 10668
rect 4028 10656 4034 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 4028 10628 4077 10656
rect 4028 10616 4034 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 5258 10656 5264 10668
rect 4295 10628 5264 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4172 10588 4200 10619
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5552 10665 5580 10696
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5718 10656 5724 10668
rect 5675 10628 5724 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 5829 10665 5857 10752
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 7009 10727 7067 10733
rect 7009 10724 7021 10727
rect 6604 10696 7021 10724
rect 6604 10684 6610 10696
rect 7009 10693 7021 10696
rect 7055 10693 7067 10727
rect 7009 10687 7067 10693
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6641 10659 6699 10665
rect 6641 10656 6653 10659
rect 6144 10628 6653 10656
rect 6144 10616 6150 10628
rect 6641 10625 6653 10628
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 7650 10616 7656 10668
rect 7708 10659 7714 10668
rect 8000 10665 8028 10764
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 14182 10792 14188 10804
rect 9916 10764 14188 10792
rect 9916 10752 9922 10764
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 14700 10764 14749 10792
rect 14700 10752 14706 10764
rect 14737 10761 14749 10764
rect 14783 10761 14795 10795
rect 15194 10792 15200 10804
rect 14737 10755 14795 10761
rect 14936 10764 15200 10792
rect 8110 10684 8116 10736
rect 8168 10684 8174 10736
rect 8220 10696 9168 10724
rect 8220 10665 8248 10696
rect 8386 10665 8392 10668
rect 7826 10659 7884 10665
rect 7708 10631 7838 10659
rect 7708 10616 7714 10631
rect 7826 10625 7838 10631
rect 7872 10625 7884 10659
rect 7826 10619 7884 10625
rect 7985 10659 8043 10665
rect 7985 10625 7997 10659
rect 8031 10625 8043 10659
rect 7985 10619 8043 10625
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8343 10659 8392 10665
rect 8343 10625 8355 10659
rect 8389 10625 8392 10659
rect 8343 10619 8392 10625
rect 4172 10560 4752 10588
rect 3329 10455 3387 10461
rect 3329 10421 3341 10455
rect 3375 10452 3387 10455
rect 3970 10452 3976 10464
rect 3375 10424 3976 10452
rect 3375 10421 3387 10424
rect 3329 10415 3387 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 4614 10452 4620 10464
rect 4571 10424 4620 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4724 10452 4752 10560
rect 5074 10548 5080 10600
rect 5132 10548 5138 10600
rect 5169 10591 5227 10597
rect 5169 10557 5181 10591
rect 5215 10557 5227 10591
rect 5169 10551 5227 10557
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 5184 10520 5212 10551
rect 5040 10492 5212 10520
rect 5460 10520 5488 10551
rect 6362 10548 6368 10600
rect 6420 10588 6426 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6420 10560 6561 10588
rect 6420 10548 6426 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 7190 10548 7196 10600
rect 7248 10588 7254 10600
rect 8220 10588 8248 10619
rect 8386 10616 8392 10619
rect 8444 10616 8450 10668
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9140 10656 9168 10696
rect 10226 10684 10232 10736
rect 10284 10724 10290 10736
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 10284 10696 11989 10724
rect 10284 10684 10290 10696
rect 11977 10693 11989 10696
rect 12023 10693 12035 10727
rect 14936 10724 14964 10764
rect 15194 10752 15200 10764
rect 15252 10792 15258 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 15252 10764 15301 10792
rect 15252 10752 15258 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 15289 10755 15347 10761
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15657 10795 15715 10801
rect 15657 10792 15669 10795
rect 15436 10764 15669 10792
rect 15436 10752 15442 10764
rect 15657 10761 15669 10764
rect 15703 10761 15715 10795
rect 15657 10755 15715 10761
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 16669 10795 16727 10801
rect 16669 10792 16681 10795
rect 16632 10764 16681 10792
rect 16632 10752 16638 10764
rect 16669 10761 16681 10764
rect 16715 10761 16727 10795
rect 16669 10755 16727 10761
rect 11977 10687 12035 10693
rect 14476 10696 14964 10724
rect 10870 10656 10876 10668
rect 9140 10628 10876 10656
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 11767 10659 11825 10665
rect 11767 10625 11779 10659
rect 11813 10625 11825 10659
rect 11767 10619 11825 10625
rect 7248 10560 8248 10588
rect 8573 10591 8631 10597
rect 7248 10548 7254 10560
rect 8573 10557 8585 10591
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 9122 10588 9128 10600
rect 8803 10560 9128 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 8110 10520 8116 10532
rect 5460 10492 8116 10520
rect 5040 10480 5046 10492
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 8481 10523 8539 10529
rect 8481 10489 8493 10523
rect 8527 10520 8539 10523
rect 8588 10520 8616 10551
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 10686 10588 10692 10600
rect 9640 10560 10692 10588
rect 9640 10548 9646 10560
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 11609 10591 11667 10597
rect 11609 10557 11621 10591
rect 11655 10557 11667 10591
rect 11782 10588 11810 10619
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 12066 10616 12072 10668
rect 12124 10616 12130 10668
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10656 12311 10659
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 12299 10628 13921 10656
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 11974 10588 11980 10600
rect 11782 10560 11980 10588
rect 11609 10551 11667 10557
rect 8527 10492 8616 10520
rect 8527 10489 8539 10492
rect 8481 10483 8539 10489
rect 9030 10480 9036 10532
rect 9088 10520 9094 10532
rect 11624 10520 11652 10551
rect 11974 10548 11980 10560
rect 12032 10548 12038 10600
rect 13814 10588 13820 10600
rect 12084 10560 13820 10588
rect 9088 10492 11652 10520
rect 9088 10480 9094 10492
rect 5534 10452 5540 10464
rect 4724 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 8665 10455 8723 10461
rect 8665 10452 8677 10455
rect 8444 10424 8677 10452
rect 8444 10412 8450 10424
rect 8665 10421 8677 10424
rect 8711 10421 8723 10455
rect 8665 10415 8723 10421
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10502 10452 10508 10464
rect 10376 10424 10508 10452
rect 10376 10412 10382 10424
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 11624 10452 11652 10492
rect 12084 10452 12112 10560
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 12158 10480 12164 10532
rect 12216 10520 12222 10532
rect 14476 10520 14504 10696
rect 15010 10684 15016 10736
rect 15068 10684 15074 10736
rect 16298 10724 16304 10736
rect 15212 10696 16304 10724
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 15212 10665 15240 10696
rect 16298 10684 16304 10696
rect 16356 10684 16362 10736
rect 16390 10684 16396 10736
rect 16448 10724 16454 10736
rect 16448 10696 17356 10724
rect 16448 10684 16454 10696
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 14608 10628 14749 10656
rect 14608 10616 14614 10628
rect 14737 10625 14749 10628
rect 14783 10625 14795 10659
rect 14737 10619 14795 10625
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10656 14979 10659
rect 15197 10659 15255 10665
rect 15197 10656 15209 10659
rect 14967 10628 15209 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 15197 10625 15209 10628
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10656 15439 10659
rect 15746 10656 15752 10668
rect 15427 10628 15752 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 14752 10588 14780 10619
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 14752 10560 15577 10588
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 12216 10492 14504 10520
rect 12216 10480 12222 10492
rect 15378 10480 15384 10532
rect 15436 10520 15442 10532
rect 15856 10520 15884 10619
rect 15948 10588 15976 10619
rect 16114 10616 16120 10668
rect 16172 10616 16178 10668
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 16264 10628 16957 10656
rect 16264 10616 16270 10628
rect 16945 10625 16957 10628
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 17328 10665 17356 10696
rect 17402 10684 17408 10736
rect 17460 10684 17466 10736
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 17313 10659 17371 10665
rect 17313 10625 17325 10659
rect 17359 10625 17371 10659
rect 17313 10619 17371 10625
rect 16850 10588 16856 10600
rect 15948 10560 16856 10588
rect 15436 10492 15884 10520
rect 15436 10480 15442 10492
rect 11624 10424 12112 10452
rect 14090 10412 14096 10464
rect 14148 10412 14154 10464
rect 14277 10455 14335 10461
rect 14277 10421 14289 10455
rect 14323 10452 14335 10455
rect 15010 10452 15016 10464
rect 14323 10424 15016 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 15102 10412 15108 10464
rect 15160 10452 15166 10464
rect 16206 10452 16212 10464
rect 15160 10424 16212 10452
rect 15160 10412 15166 10424
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16776 10452 16804 10560
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 17144 10520 17172 10619
rect 17678 10616 17684 10668
rect 17736 10616 17742 10668
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 18104 10628 18153 10656
rect 18104 10616 18110 10628
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 18141 10619 18199 10625
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 17276 10560 17509 10588
rect 17276 10548 17282 10560
rect 17497 10557 17509 10560
rect 17543 10588 17555 10591
rect 17543 10560 18000 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 17972 10529 18000 10560
rect 17865 10523 17923 10529
rect 17865 10520 17877 10523
rect 17144 10492 17877 10520
rect 17865 10489 17877 10492
rect 17911 10489 17923 10523
rect 17865 10483 17923 10489
rect 17957 10523 18015 10529
rect 17957 10489 17969 10523
rect 18003 10489 18015 10523
rect 17957 10483 18015 10489
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 16776 10424 17417 10452
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 1104 10362 18492 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 18492 10362
rect 1104 10288 18492 10310
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 9030 10248 9036 10260
rect 3016 10220 5580 10248
rect 3016 10208 3022 10220
rect 4982 10180 4988 10192
rect 4080 10152 4988 10180
rect 4080 10056 4108 10152
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 4614 10112 4620 10124
rect 4264 10084 4620 10112
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 2866 10004 2872 10056
rect 2924 10044 2930 10056
rect 3786 10044 3792 10056
rect 2924 10016 3792 10044
rect 2924 10004 2930 10016
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 3970 10004 3976 10056
rect 4028 10004 4034 10056
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4264 10053 4292 10084
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 5166 10072 5172 10124
rect 5224 10112 5230 10124
rect 5350 10112 5356 10124
rect 5224 10084 5356 10112
rect 5224 10072 5230 10084
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 5552 10112 5580 10220
rect 5828 10220 9036 10248
rect 5718 10112 5724 10124
rect 5552 10084 5724 10112
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 5074 10044 5080 10056
rect 4396 10016 5080 10044
rect 4396 10004 4402 10016
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5552 10053 5580 10084
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 5828 10053 5856 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9398 10208 9404 10260
rect 9456 10208 9462 10260
rect 9858 10208 9864 10260
rect 9916 10208 9922 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 9968 10220 11437 10248
rect 6089 10183 6147 10189
rect 6089 10149 6101 10183
rect 6135 10149 6147 10183
rect 6089 10143 6147 10149
rect 6104 10112 6132 10143
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 7926 10180 7932 10192
rect 7156 10152 7932 10180
rect 7156 10140 7162 10152
rect 7926 10140 7932 10152
rect 7984 10180 7990 10192
rect 9214 10180 9220 10192
rect 7984 10152 9220 10180
rect 7984 10140 7990 10152
rect 9214 10140 9220 10152
rect 9272 10140 9278 10192
rect 9876 10180 9904 10208
rect 9416 10152 9904 10180
rect 9416 10124 9444 10152
rect 6104 10084 8156 10112
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 5538 10047 5596 10053
rect 5538 10013 5550 10047
rect 5584 10013 5596 10047
rect 5538 10007 5596 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 5951 10047 6009 10053
rect 5951 10013 5963 10047
rect 5997 10044 6009 10047
rect 6362 10044 6368 10056
rect 5997 10016 6368 10044
rect 5997 10013 6009 10016
rect 5951 10007 6009 10013
rect 3804 9976 3832 10004
rect 5460 9976 5488 10007
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 7098 10004 7104 10056
rect 7156 10004 7162 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 3804 9948 5488 9976
rect 5718 9936 5724 9988
rect 5776 9936 5782 9988
rect 6273 9979 6331 9985
rect 6273 9945 6285 9979
rect 6319 9976 6331 9979
rect 6546 9976 6552 9988
rect 6319 9948 6552 9976
rect 6319 9945 6331 9948
rect 6273 9939 6331 9945
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 1486 9868 1492 9920
rect 1544 9868 1550 9920
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3108 9880 3801 9908
rect 3108 9868 3114 9880
rect 3789 9877 3801 9880
rect 3835 9877 3847 9911
rect 3789 9871 3847 9877
rect 5626 9868 5632 9920
rect 5684 9908 5690 9920
rect 7208 9908 7236 10007
rect 7466 10004 7472 10056
rect 7524 10004 7530 10056
rect 8128 10053 8156 10084
rect 9398 10072 9404 10124
rect 9456 10072 9462 10124
rect 9858 10112 9864 10124
rect 9692 10084 9864 10112
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 8113 10047 8171 10053
rect 7607 10016 7880 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 7374 9936 7380 9988
rect 7432 9936 7438 9988
rect 5684 9880 7236 9908
rect 5684 9868 5690 9880
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 7852 9908 7880 10016
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 8386 10004 8392 10056
rect 8444 10004 8450 10056
rect 9692 10053 9720 10084
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 9968 10056 9996 10220
rect 11425 10217 11437 10220
rect 11471 10248 11483 10251
rect 11882 10248 11888 10260
rect 11471 10220 11888 10248
rect 11471 10217 11483 10220
rect 11425 10211 11483 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 12066 10208 12072 10260
rect 12124 10208 12130 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15565 10251 15623 10257
rect 15565 10248 15577 10251
rect 15344 10220 15577 10248
rect 15344 10208 15350 10220
rect 15565 10217 15577 10220
rect 15611 10248 15623 10251
rect 16206 10248 16212 10260
rect 15611 10220 16212 10248
rect 15611 10217 15623 10220
rect 15565 10211 15623 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16393 10251 16451 10257
rect 16393 10217 16405 10251
rect 16439 10248 16451 10251
rect 16666 10248 16672 10260
rect 16439 10220 16672 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 17034 10208 17040 10260
rect 17092 10248 17098 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17092 10220 17693 10248
rect 17092 10208 17098 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 17681 10211 17739 10217
rect 15194 10180 15200 10192
rect 10980 10152 15200 10180
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10318 10112 10324 10124
rect 10091 10084 10324 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 10873 10115 10931 10121
rect 10873 10112 10885 10115
rect 10744 10084 10885 10112
rect 10744 10072 10750 10084
rect 10873 10081 10885 10084
rect 10919 10081 10931 10115
rect 10873 10075 10931 10081
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 9769 10047 9827 10053
rect 9769 10013 9781 10047
rect 9815 10044 9827 10047
rect 9950 10044 9956 10056
rect 9815 10016 9956 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 9950 10004 9956 10016
rect 10008 10004 10014 10056
rect 10134 10004 10140 10056
rect 10192 10004 10198 10056
rect 10226 10004 10232 10056
rect 10284 10004 10290 10056
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 10778 10004 10784 10056
rect 10836 10004 10842 10056
rect 10980 10053 11008 10152
rect 15194 10140 15200 10152
rect 15252 10180 15258 10192
rect 16114 10180 16120 10192
rect 15252 10152 16120 10180
rect 15252 10140 15258 10152
rect 16114 10140 16120 10152
rect 16172 10140 16178 10192
rect 15654 10112 15660 10124
rect 11532 10084 15660 10112
rect 10965 10047 11023 10053
rect 10965 10013 10977 10047
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11330 10004 11336 10056
rect 11388 10004 11394 10056
rect 11532 10053 11560 10084
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 11790 10004 11796 10056
rect 11848 10044 11854 10056
rect 15396 10053 15424 10084
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 15764 10084 16620 10112
rect 15562 10053 15568 10056
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 11848 10016 11989 10044
rect 11848 10004 11854 10016
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 15535 10047 15568 10053
rect 15535 10013 15547 10047
rect 15535 10007 15568 10013
rect 7929 9979 7987 9985
rect 7929 9945 7941 9979
rect 7975 9976 7987 9979
rect 8478 9976 8484 9988
rect 7975 9948 8484 9976
rect 7975 9945 7987 9948
rect 7929 9939 7987 9945
rect 8478 9936 8484 9948
rect 8536 9936 8542 9988
rect 8570 9936 8576 9988
rect 8628 9976 8634 9988
rect 9858 9976 9864 9988
rect 8628 9948 9864 9976
rect 8628 9936 8634 9948
rect 9858 9936 9864 9948
rect 9916 9936 9922 9988
rect 10689 9979 10747 9985
rect 10689 9976 10701 9979
rect 10152 9948 10701 9976
rect 10152 9920 10180 9948
rect 10689 9945 10701 9948
rect 10735 9945 10747 9979
rect 10689 9939 10747 9945
rect 11054 9936 11060 9988
rect 11112 9976 11118 9988
rect 12176 9976 12204 10007
rect 15562 10004 15568 10007
rect 15620 10004 15626 10056
rect 13906 9976 13912 9988
rect 11112 9948 13912 9976
rect 11112 9936 11118 9948
rect 13906 9936 13912 9948
rect 13964 9936 13970 9988
rect 14090 9936 14096 9988
rect 14148 9976 14154 9988
rect 15764 9976 15792 10084
rect 16482 10044 16488 10056
rect 14148 9948 15792 9976
rect 15856 10016 16488 10044
rect 14148 9936 14154 9948
rect 8110 9908 8116 9920
rect 7852 9880 8116 9908
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 9398 9908 9404 9920
rect 8343 9880 9404 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 10134 9868 10140 9920
rect 10192 9868 10198 9920
rect 10318 9868 10324 9920
rect 10376 9868 10382 9920
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 10962 9908 10968 9920
rect 10560 9880 10968 9908
rect 10560 9868 10566 9880
rect 10962 9868 10968 9880
rect 11020 9908 11026 9920
rect 12802 9908 12808 9920
rect 11020 9880 12808 9908
rect 11020 9868 11026 9880
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 15856 9908 15884 10016
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16592 10044 16620 10084
rect 16666 10072 16672 10124
rect 16724 10112 16730 10124
rect 16724 10084 18000 10112
rect 16724 10072 16730 10084
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16592 10016 16865 10044
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 17037 10047 17095 10053
rect 17037 10044 17049 10047
rect 17000 10016 17049 10044
rect 17000 10004 17006 10016
rect 17037 10013 17049 10016
rect 17083 10044 17095 10047
rect 17083 10016 17264 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 16022 9936 16028 9988
rect 16080 9936 16086 9988
rect 16114 9936 16120 9988
rect 16172 9976 16178 9988
rect 16209 9979 16267 9985
rect 16209 9976 16221 9979
rect 16172 9948 16221 9976
rect 16172 9936 16178 9948
rect 16209 9945 16221 9948
rect 16255 9945 16267 9979
rect 16209 9939 16267 9945
rect 16298 9936 16304 9988
rect 16356 9976 16362 9988
rect 17129 9979 17187 9985
rect 17129 9976 17141 9979
rect 16356 9948 17141 9976
rect 16356 9936 16362 9948
rect 17129 9945 17141 9948
rect 17175 9945 17187 9979
rect 17236 9976 17264 10016
rect 17310 10004 17316 10056
rect 17368 10004 17374 10056
rect 17402 10004 17408 10056
rect 17460 10004 17466 10056
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10044 17555 10047
rect 17586 10044 17592 10056
rect 17543 10016 17592 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 17862 10004 17868 10056
rect 17920 10004 17926 10056
rect 17972 10053 18000 10084
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 17681 9979 17739 9985
rect 17681 9976 17693 9979
rect 17236 9948 17693 9976
rect 17129 9939 17187 9945
rect 17681 9945 17693 9948
rect 17727 9945 17739 9979
rect 17681 9939 17739 9945
rect 13136 9880 15884 9908
rect 16853 9911 16911 9917
rect 13136 9868 13142 9880
rect 16853 9877 16865 9911
rect 16899 9908 16911 9911
rect 17034 9908 17040 9920
rect 16899 9880 17040 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 1104 9818 18492 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 18492 9818
rect 1104 9744 18492 9766
rect 1489 9707 1547 9713
rect 1489 9673 1501 9707
rect 1535 9704 1547 9707
rect 1670 9704 1676 9716
rect 1535 9676 1676 9704
rect 1535 9673 1547 9676
rect 1489 9667 1547 9673
rect 1670 9664 1676 9676
rect 1728 9664 1734 9716
rect 2516 9676 4016 9704
rect 2314 9596 2320 9648
rect 2372 9596 2378 9648
rect 1854 9528 1860 9580
rect 1912 9528 1918 9580
rect 1946 9528 1952 9580
rect 2004 9568 2010 9580
rect 2406 9568 2412 9580
rect 2004 9540 2412 9568
rect 2004 9528 2010 9540
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 2516 9577 2544 9676
rect 3421 9639 3479 9645
rect 3421 9636 3433 9639
rect 2792 9608 3433 9636
rect 2792 9580 2820 9608
rect 3421 9605 3433 9608
rect 3467 9636 3479 9639
rect 3602 9636 3608 9648
rect 3467 9608 3608 9636
rect 3467 9605 3479 9608
rect 3421 9599 3479 9605
rect 3602 9596 3608 9608
rect 3660 9596 3666 9648
rect 3988 9645 4016 9676
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 5353 9707 5411 9713
rect 5353 9704 5365 9707
rect 5132 9676 5365 9704
rect 5132 9664 5138 9676
rect 5353 9673 5365 9676
rect 5399 9704 5411 9707
rect 5534 9704 5540 9716
rect 5399 9676 5540 9704
rect 5399 9673 5411 9676
rect 5353 9667 5411 9673
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 6365 9707 6423 9713
rect 6365 9704 6377 9707
rect 5776 9676 6377 9704
rect 5776 9664 5782 9676
rect 6365 9673 6377 9676
rect 6411 9673 6423 9707
rect 7006 9704 7012 9716
rect 6365 9667 6423 9673
rect 6472 9676 7012 9704
rect 3973 9639 4031 9645
rect 3743 9605 3801 9611
rect 3743 9590 3755 9605
rect 3712 9580 3755 9590
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2648 9540 2697 9568
rect 2648 9528 2654 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2774 9528 2780 9580
rect 2832 9528 2838 9580
rect 2958 9528 2964 9580
rect 3016 9568 3022 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 3016 9540 3065 9568
rect 3016 9528 3022 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 3142 9528 3148 9580
rect 3200 9528 3206 9580
rect 3694 9528 3700 9580
rect 3752 9571 3755 9580
rect 3789 9602 3801 9605
rect 3973 9605 3985 9639
rect 4019 9636 4031 9639
rect 4062 9636 4068 9648
rect 4019 9608 4068 9636
rect 4019 9605 4031 9608
rect 3789 9571 3816 9602
rect 3973 9599 4031 9605
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 5626 9636 5632 9648
rect 4908 9608 5120 9636
rect 4908 9577 4936 9608
rect 3752 9562 3816 9571
rect 4893 9571 4951 9577
rect 3752 9528 3758 9562
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5092 9568 5120 9608
rect 5368 9608 5632 9636
rect 5368 9568 5396 9608
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 6472 9636 6500 9676
rect 7006 9664 7012 9676
rect 7064 9704 7070 9716
rect 7064 9676 7512 9704
rect 7064 9664 7070 9676
rect 6730 9636 6736 9648
rect 6012 9608 6500 9636
rect 6559 9608 6736 9636
rect 5092 9540 5396 9568
rect 5534 9528 5540 9580
rect 5592 9528 5598 9580
rect 6012 9577 6040 9608
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6193 9571 6251 9577
rect 6193 9537 6205 9571
rect 6239 9568 6251 9571
rect 6362 9568 6368 9580
rect 6239 9540 6368 9568
rect 6239 9537 6251 9540
rect 6193 9531 6251 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6559 9577 6587 9608
rect 6730 9596 6736 9608
rect 6788 9596 6794 9648
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 2130 9460 2136 9512
rect 2188 9460 2194 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9500 5227 9503
rect 5258 9500 5264 9512
rect 5215 9472 5264 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 3528 9432 3556 9463
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 6638 9494 6644 9546
rect 6696 9494 6702 9546
rect 6730 9494 6736 9546
rect 6788 9494 6794 9546
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 7484 9577 7512 9676
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 9309 9707 9367 9713
rect 7800 9676 8294 9704
rect 7800 9664 7806 9676
rect 8266 9636 8294 9676
rect 9309 9673 9321 9707
rect 9355 9704 9367 9707
rect 9490 9704 9496 9716
rect 9355 9676 9496 9704
rect 9355 9673 9367 9676
rect 9309 9667 9367 9673
rect 9490 9664 9496 9676
rect 9548 9704 9554 9716
rect 10226 9704 10232 9716
rect 9548 9676 10232 9704
rect 9548 9664 9554 9676
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 12986 9664 12992 9716
rect 13044 9704 13050 9716
rect 13354 9704 13360 9716
rect 13044 9676 13360 9704
rect 13044 9664 13050 9676
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 8266 9608 9904 9636
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 7558 9528 7564 9580
rect 7616 9528 7622 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7837 9571 7895 9577
rect 7837 9568 7849 9571
rect 7791 9540 7849 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7837 9537 7849 9540
rect 7883 9537 7895 9571
rect 7837 9531 7895 9537
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8202 9568 8208 9580
rect 8067 9540 8208 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9214 9568 9220 9580
rect 9079 9540 9220 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9582 9528 9588 9580
rect 9640 9528 9646 9580
rect 9876 9577 9904 9608
rect 10042 9596 10048 9648
rect 10100 9636 10106 9648
rect 12250 9636 12256 9648
rect 10100 9608 12256 9636
rect 10100 9596 10106 9608
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 12820 9608 14412 9636
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10410 9568 10416 9580
rect 9999 9540 10416 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 11054 9528 11060 9580
rect 11112 9528 11118 9580
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 11882 9568 11888 9580
rect 11287 9540 11888 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12492 9540 12541 9568
rect 12492 9528 12498 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12710 9528 12716 9580
rect 12768 9577 12774 9580
rect 12768 9571 12783 9577
rect 12771 9568 12783 9571
rect 12820 9568 12848 9608
rect 12771 9540 12848 9568
rect 12989 9571 13047 9577
rect 12771 9537 12783 9540
rect 12768 9531 12783 9537
rect 12989 9537 13001 9571
rect 13035 9558 13047 9571
rect 13078 9558 13084 9570
rect 13035 9537 13084 9558
rect 12989 9531 13084 9537
rect 12768 9528 12774 9531
rect 13004 9530 13084 9531
rect 13078 9518 13084 9530
rect 13136 9518 13142 9570
rect 13170 9528 13176 9580
rect 13228 9528 13234 9580
rect 13449 9571 13507 9577
rect 13449 9537 13461 9571
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13906 9571 13964 9577
rect 13906 9537 13918 9571
rect 13952 9558 13964 9571
rect 13998 9558 14004 9580
rect 13952 9537 14004 9558
rect 13906 9531 14004 9537
rect 6825 9503 6883 9509
rect 6641 9469 6653 9494
rect 6687 9469 6699 9494
rect 6641 9463 6699 9469
rect 6733 9469 6745 9494
rect 6779 9469 6791 9494
rect 6733 9463 6791 9469
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 3605 9435 3663 9441
rect 3605 9432 3617 9435
rect 3528 9404 3617 9432
rect 3605 9401 3617 9404
rect 3651 9401 3663 9435
rect 4338 9432 4344 9444
rect 3605 9395 3663 9401
rect 3712 9404 4344 9432
rect 2866 9324 2872 9376
rect 2924 9324 2930 9376
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3712 9364 3740 9404
rect 4338 9392 4344 9404
rect 4396 9392 4402 9444
rect 5997 9435 6055 9441
rect 5997 9401 6009 9435
rect 6043 9432 6055 9435
rect 6086 9432 6092 9444
rect 6043 9404 6092 9432
rect 6043 9401 6055 9404
rect 5997 9395 6055 9401
rect 6086 9392 6092 9404
rect 6144 9432 6150 9444
rect 6840 9432 6868 9463
rect 7282 9460 7288 9512
rect 7340 9460 7346 9512
rect 8570 9460 8576 9512
rect 8628 9500 8634 9512
rect 8938 9500 8944 9512
rect 8628 9472 8944 9500
rect 8628 9460 8634 9472
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9469 10195 9503
rect 13456 9500 13484 9531
rect 10137 9463 10195 9469
rect 13280 9472 13484 9500
rect 6144 9404 6868 9432
rect 6144 9392 6150 9404
rect 8110 9392 8116 9444
rect 8168 9432 8174 9444
rect 8168 9404 9904 9432
rect 8168 9392 8174 9404
rect 3016 9336 3740 9364
rect 3789 9367 3847 9373
rect 3016 9324 3022 9336
rect 3789 9333 3801 9367
rect 3835 9364 3847 9367
rect 5166 9364 5172 9376
rect 3835 9336 5172 9364
rect 3835 9333 3847 9336
rect 3789 9327 3847 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 5902 9364 5908 9376
rect 5776 9336 5908 9364
rect 5776 9324 5782 9336
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 7834 9324 7840 9376
rect 7892 9324 7898 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 9582 9364 9588 9376
rect 8444 9336 9588 9364
rect 8444 9324 8450 9336
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9674 9324 9680 9376
rect 9732 9324 9738 9376
rect 9876 9364 9904 9404
rect 9950 9392 9956 9444
rect 10008 9432 10014 9444
rect 10060 9432 10088 9463
rect 10008 9404 10088 9432
rect 10152 9432 10180 9463
rect 10410 9432 10416 9444
rect 10152 9404 10416 9432
rect 10008 9392 10014 9404
rect 10410 9392 10416 9404
rect 10468 9392 10474 9444
rect 11057 9435 11115 9441
rect 11057 9401 11069 9435
rect 11103 9432 11115 9435
rect 11146 9432 11152 9444
rect 11103 9404 11152 9432
rect 11103 9401 11115 9404
rect 11057 9395 11115 9401
rect 11146 9392 11152 9404
rect 11204 9432 11210 9444
rect 12158 9432 12164 9444
rect 11204 9404 12164 9432
rect 11204 9392 11210 9404
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 13280 9432 13308 9472
rect 13538 9460 13544 9512
rect 13596 9460 13602 9512
rect 13633 9503 13691 9509
rect 13633 9469 13645 9503
rect 13679 9469 13691 9503
rect 13740 9500 13768 9531
rect 13924 9530 14004 9531
rect 13998 9528 14004 9530
rect 14056 9528 14062 9580
rect 14384 9577 14412 9608
rect 16850 9596 16856 9648
rect 16908 9636 16914 9648
rect 17681 9639 17739 9645
rect 17681 9636 17693 9639
rect 16908 9608 17693 9636
rect 16908 9596 16914 9608
rect 17681 9605 17693 9608
rect 17727 9605 17739 9639
rect 17681 9599 17739 9605
rect 17865 9639 17923 9645
rect 17865 9605 17877 9639
rect 17911 9636 17923 9639
rect 18138 9636 18144 9648
rect 17911 9608 18144 9636
rect 17911 9605 17923 9608
rect 17865 9599 17923 9605
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9568 14427 9571
rect 14918 9568 14924 9580
rect 14415 9540 14924 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 17696 9568 17724 9599
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 18046 9568 18052 9580
rect 17696 9540 18052 9568
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 14277 9503 14335 9509
rect 13740 9472 14044 9500
rect 13633 9463 13691 9469
rect 12860 9404 13308 9432
rect 12860 9392 12866 9404
rect 13354 9392 13360 9444
rect 13412 9432 13418 9444
rect 13648 9432 13676 9463
rect 14016 9441 14044 9472
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 14323 9472 15976 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 13412 9404 13676 9432
rect 14001 9435 14059 9441
rect 13412 9392 13418 9404
rect 14001 9401 14013 9435
rect 14047 9401 14059 9435
rect 14001 9395 14059 9401
rect 11514 9364 11520 9376
rect 9876 9336 11520 9364
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 12710 9364 12716 9376
rect 12584 9336 12716 9364
rect 12584 9324 12590 9336
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 12986 9364 12992 9376
rect 12943 9336 12992 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 13265 9367 13323 9373
rect 13265 9333 13277 9367
rect 13311 9364 13323 9367
rect 13630 9364 13636 9376
rect 13311 9336 13636 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 14274 9324 14280 9376
rect 14332 9324 14338 9376
rect 15948 9364 15976 9472
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 17310 9500 17316 9512
rect 16908 9472 17316 9500
rect 16908 9460 16914 9472
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 17494 9460 17500 9512
rect 17552 9460 17558 9512
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 17129 9435 17187 9441
rect 17129 9432 17141 9435
rect 16080 9404 17141 9432
rect 16080 9392 16086 9404
rect 17129 9401 17141 9404
rect 17175 9401 17187 9435
rect 17129 9395 17187 9401
rect 17770 9364 17776 9376
rect 15948 9336 17776 9364
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 1104 9274 18492 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 18492 9274
rect 1104 9200 18492 9222
rect 1673 9163 1731 9169
rect 1673 9129 1685 9163
rect 1719 9160 1731 9163
rect 1854 9160 1860 9172
rect 1719 9132 1860 9160
rect 1719 9129 1731 9132
rect 1673 9123 1731 9129
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 2096 9132 2237 9160
rect 2096 9120 2102 9132
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 2225 9123 2283 9129
rect 3418 9120 3424 9172
rect 3476 9120 3482 9172
rect 3878 9120 3884 9172
rect 3936 9120 3942 9172
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 4982 9160 4988 9172
rect 4672 9132 4988 9160
rect 4672 9120 4678 9132
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 5169 9163 5227 9169
rect 5169 9129 5181 9163
rect 5215 9160 5227 9163
rect 5350 9160 5356 9172
rect 5215 9132 5356 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 5629 9163 5687 9169
rect 5629 9129 5641 9163
rect 5675 9160 5687 9163
rect 5718 9160 5724 9172
rect 5675 9132 5724 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 7466 9160 7472 9172
rect 5828 9132 7472 9160
rect 2056 9024 2084 9120
rect 3283 9095 3341 9101
rect 3283 9061 3295 9095
rect 3329 9092 3341 9095
rect 3896 9092 3924 9120
rect 5828 9092 5856 9132
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 8018 9160 8024 9172
rect 7576 9132 8024 9160
rect 3329 9064 3924 9092
rect 4080 9064 5856 9092
rect 3329 9061 3341 9064
rect 3283 9055 3341 9061
rect 4080 9036 4108 9064
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 6917 9095 6975 9101
rect 6917 9092 6929 9095
rect 6788 9064 6929 9092
rect 6788 9052 6794 9064
rect 6917 9061 6929 9064
rect 6963 9092 6975 9095
rect 6963 9064 7149 9092
rect 6963 9061 6975 9064
rect 6917 9055 6975 9061
rect 2958 9024 2964 9036
rect 1872 8996 2084 9024
rect 2700 8996 2964 9024
rect 1872 8965 1900 8996
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2222 8956 2228 8968
rect 2179 8928 2228 8956
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 1762 8848 1768 8900
rect 1820 8888 1826 8900
rect 1964 8888 1992 8919
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 2314 8916 2320 8968
rect 2372 8916 2378 8968
rect 2406 8916 2412 8968
rect 2464 8916 2470 8968
rect 2700 8965 2728 8996
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3068 8996 3648 9024
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 2424 8888 2452 8916
rect 1820 8860 2452 8888
rect 2792 8888 2820 8919
rect 2866 8916 2872 8968
rect 2924 8916 2930 8968
rect 3068 8965 3096 8996
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8956 3203 8959
rect 3418 8956 3424 8968
rect 3191 8928 3424 8956
rect 3191 8925 3203 8928
rect 3145 8919 3203 8925
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 3620 8965 3648 8996
rect 4062 8984 4068 9036
rect 4120 8984 4126 9036
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 4890 9024 4896 9036
rect 4580 8996 4896 9024
rect 4580 8984 4586 8996
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 3786 8956 3792 8968
rect 3651 8928 3792 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 4338 8916 4344 8968
rect 4396 8916 4402 8968
rect 4816 8965 4844 8996
rect 4890 8984 4896 8996
rect 4948 9024 4954 9036
rect 4948 8996 5304 9024
rect 4948 8984 4954 8996
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 4982 8916 4988 8968
rect 5040 8916 5046 8968
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5166 8956 5172 8968
rect 5123 8928 5172 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 5276 8965 5304 8996
rect 5552 8996 6684 9024
rect 5552 8965 5580 8996
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5684 8928 5733 8956
rect 5684 8916 5690 8928
rect 5721 8925 5733 8928
rect 5767 8956 5779 8959
rect 5994 8956 6000 8968
rect 5767 8928 6000 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 5994 8916 6000 8928
rect 6052 8956 6058 8968
rect 6656 8965 6684 8996
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 6052 8928 6377 8956
rect 6052 8916 6058 8928
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 6822 8956 6828 8968
rect 6687 8928 6828 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 7121 8956 7149 9064
rect 7282 9052 7288 9104
rect 7340 9092 7346 9104
rect 7576 9092 7604 9132
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8662 9120 8668 9172
rect 8720 9160 8726 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8720 9132 9045 9160
rect 8720 9120 8726 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 10686 9160 10692 9172
rect 9364 9132 10692 9160
rect 9364 9120 9370 9132
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11054 9120 11060 9172
rect 11112 9120 11118 9172
rect 12526 9160 12532 9172
rect 11256 9132 12532 9160
rect 9398 9092 9404 9104
rect 7340 9064 7604 9092
rect 7760 9064 9404 9092
rect 7340 9052 7346 9064
rect 7760 8956 7788 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 9585 9095 9643 9101
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 11256 9092 11284 9132
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 14182 9160 14188 9172
rect 13504 9132 14188 9160
rect 13504 9120 13510 9132
rect 14182 9120 14188 9132
rect 14240 9160 14246 9172
rect 15562 9160 15568 9172
rect 14240 9132 15568 9160
rect 14240 9120 14246 9132
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 16298 9120 16304 9172
rect 16356 9120 16362 9172
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16761 9163 16819 9169
rect 16761 9160 16773 9163
rect 16632 9132 16773 9160
rect 16632 9120 16638 9132
rect 16761 9129 16773 9132
rect 16807 9129 16819 9163
rect 16761 9123 16819 9129
rect 16850 9120 16856 9172
rect 16908 9160 16914 9172
rect 17037 9163 17095 9169
rect 17037 9160 17049 9163
rect 16908 9132 17049 9160
rect 16908 9120 16914 9132
rect 17037 9129 17049 9132
rect 17083 9129 17095 9163
rect 17037 9123 17095 9129
rect 9631 9064 11284 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 11330 9052 11336 9104
rect 11388 9092 11394 9104
rect 11425 9095 11483 9101
rect 11425 9092 11437 9095
rect 11388 9064 11437 9092
rect 11388 9052 11394 9064
rect 11425 9061 11437 9064
rect 11471 9092 11483 9095
rect 11701 9095 11759 9101
rect 11701 9092 11713 9095
rect 11471 9064 11713 9092
rect 11471 9061 11483 9064
rect 11425 9055 11483 9061
rect 11701 9061 11713 9064
rect 11747 9061 11759 9095
rect 11701 9055 11759 9061
rect 11793 9095 11851 9101
rect 11793 9061 11805 9095
rect 11839 9092 11851 9095
rect 11974 9092 11980 9104
rect 11839 9064 11980 9092
rect 11839 9061 11851 9064
rect 11793 9055 11851 9061
rect 11974 9052 11980 9064
rect 12032 9052 12038 9104
rect 12158 9052 12164 9104
rect 12216 9092 12222 9104
rect 13354 9092 13360 9104
rect 12216 9064 13360 9092
rect 12216 9052 12222 9064
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 16316 9092 16344 9120
rect 16132 9064 16344 9092
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 11609 9027 11667 9033
rect 7892 8996 10364 9024
rect 7892 8984 7898 8996
rect 7121 8928 7788 8956
rect 7926 8916 7932 8968
rect 7984 8956 7990 8968
rect 7984 8928 8524 8956
rect 7984 8916 7990 8928
rect 4706 8888 4712 8900
rect 2792 8860 4712 8888
rect 1820 8848 1826 8860
rect 4706 8848 4712 8860
rect 4764 8848 4770 8900
rect 4908 8860 6132 8888
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2409 8823 2467 8829
rect 2409 8820 2421 8823
rect 2372 8792 2421 8820
rect 2372 8780 2378 8792
rect 2409 8789 2421 8792
rect 2455 8789 2467 8823
rect 2409 8783 2467 8789
rect 3602 8780 3608 8832
rect 3660 8780 3666 8832
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 4908 8820 4936 8860
rect 3936 8792 4936 8820
rect 4985 8823 5043 8829
rect 3936 8780 3942 8792
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5718 8820 5724 8832
rect 5031 8792 5724 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 5905 8823 5963 8829
rect 5905 8789 5917 8823
rect 5951 8820 5963 8823
rect 5994 8820 6000 8832
rect 5951 8792 6000 8820
rect 5951 8789 5963 8792
rect 5905 8783 5963 8789
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 6104 8820 6132 8860
rect 6178 8848 6184 8900
rect 6236 8848 6242 8900
rect 7193 8891 7251 8897
rect 7193 8857 7205 8891
rect 7239 8888 7251 8891
rect 7466 8888 7472 8900
rect 7239 8860 7472 8888
rect 7239 8857 7251 8860
rect 7193 8851 7251 8857
rect 7466 8848 7472 8860
rect 7524 8848 7530 8900
rect 8205 8891 8263 8897
rect 8205 8857 8217 8891
rect 8251 8857 8263 8891
rect 8496 8888 8524 8928
rect 8570 8916 8576 8968
rect 8628 8916 8634 8968
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8956 9183 8959
rect 9398 8956 9404 8968
rect 9171 8928 9404 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 9582 8888 9588 8900
rect 8496 8860 9588 8888
rect 8205 8851 8263 8857
rect 6362 8820 6368 8832
rect 6104 8792 6368 8820
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 7926 8780 7932 8832
rect 7984 8820 7990 8832
rect 8220 8820 8248 8851
rect 9582 8848 9588 8860
rect 9640 8888 9646 8900
rect 9784 8888 9812 8919
rect 9640 8860 9812 8888
rect 9876 8888 9904 8919
rect 9950 8916 9956 8968
rect 10008 8916 10014 8968
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8956 10103 8959
rect 10134 8956 10140 8968
rect 10091 8928 10140 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10336 8965 10364 8996
rect 11609 8993 11621 9027
rect 11655 9024 11667 9027
rect 12250 9024 12256 9036
rect 11655 8996 12256 9024
rect 11655 8993 11667 8996
rect 11609 8987 11667 8993
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 13449 9027 13507 9033
rect 13449 9024 13461 9027
rect 12584 8996 13461 9024
rect 12584 8984 12590 8996
rect 13449 8993 13461 8996
rect 13495 8993 13507 9027
rect 13449 8987 13507 8993
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 16132 9033 16160 9064
rect 16666 9052 16672 9104
rect 16724 9092 16730 9104
rect 17313 9095 17371 9101
rect 17313 9092 17325 9095
rect 16724 9064 17325 9092
rect 16724 9052 16730 9064
rect 17313 9061 17325 9064
rect 17359 9092 17371 9095
rect 17678 9092 17684 9104
rect 17359 9064 17684 9092
rect 17359 9061 17371 9064
rect 17313 9055 17371 9061
rect 17678 9052 17684 9064
rect 17736 9052 17742 9104
rect 15197 9027 15255 9033
rect 15197 8993 15209 9027
rect 15243 9024 15255 9027
rect 15565 9027 15623 9033
rect 15565 9024 15577 9027
rect 15243 8996 15577 9024
rect 15243 8993 15255 8996
rect 15197 8987 15255 8993
rect 15565 8993 15577 8996
rect 15611 8993 15623 9027
rect 15565 8987 15623 8993
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 8993 16175 9027
rect 16117 8987 16175 8993
rect 16206 8984 16212 9036
rect 16264 8984 16270 9036
rect 17402 9024 17408 9036
rect 16408 8996 17408 9024
rect 16408 8968 16436 8996
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 10244 8888 10272 8919
rect 10520 8888 10548 8919
rect 10594 8916 10600 8968
rect 10652 8916 10658 8968
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8956 11299 8959
rect 11517 8959 11575 8965
rect 11287 8928 11376 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 11054 8888 11060 8900
rect 9876 8860 9996 8888
rect 10244 8860 10364 8888
rect 10520 8860 11060 8888
rect 9640 8848 9646 8860
rect 9968 8832 9996 8860
rect 10336 8832 10364 8860
rect 11054 8848 11060 8860
rect 11112 8848 11118 8900
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 7984 8792 8401 8820
rect 7984 8780 7990 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9950 8820 9956 8832
rect 8812 8792 9956 8820
rect 8812 8780 8818 8792
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10318 8780 10324 8832
rect 10376 8780 10382 8832
rect 10778 8780 10784 8832
rect 10836 8780 10842 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11348 8820 11376 8928
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 13078 8956 13084 8968
rect 11931 8928 13084 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 11532 8888 11560 8919
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8956 13599 8959
rect 14182 8956 14188 8968
rect 13587 8928 14188 8956
rect 13587 8925 13599 8928
rect 13541 8919 13599 8925
rect 13372 8888 13400 8919
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 14550 8956 14556 8968
rect 14424 8928 14556 8956
rect 14424 8916 14430 8928
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 14734 8916 14740 8968
rect 14792 8916 14798 8968
rect 14826 8916 14832 8968
rect 14884 8916 14890 8968
rect 14918 8916 14924 8968
rect 14976 8916 14982 8968
rect 15470 8916 15476 8968
rect 15528 8916 15534 8968
rect 15654 8916 15660 8968
rect 15712 8916 15718 8968
rect 15746 8916 15752 8968
rect 15804 8916 15810 8968
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 15896 8928 16313 8956
rect 15896 8916 15902 8928
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 16301 8919 16359 8925
rect 16390 8916 16396 8968
rect 16448 8916 16454 8968
rect 16776 8965 16804 8996
rect 17402 8984 17408 8996
rect 17460 8984 17466 9036
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8925 16635 8959
rect 16577 8919 16635 8925
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8925 16819 8959
rect 16761 8919 16819 8925
rect 16945 8959 17003 8965
rect 16945 8925 16957 8959
rect 16991 8956 17003 8959
rect 17126 8956 17132 8968
rect 16991 8928 17132 8956
rect 16991 8925 17003 8928
rect 16945 8919 17003 8925
rect 15289 8891 15347 8897
rect 15289 8888 15301 8891
rect 11532 8860 12572 8888
rect 13372 8860 15301 8888
rect 11974 8820 11980 8832
rect 11204 8792 11980 8820
rect 11204 8780 11210 8792
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 12544 8820 12572 8860
rect 15289 8857 15301 8860
rect 15335 8857 15347 8891
rect 15289 8851 15347 8857
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 16592 8888 16620 8919
rect 16264 8860 16620 8888
rect 16264 8848 16270 8860
rect 12894 8820 12900 8832
rect 12544 8792 12900 8820
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13170 8780 13176 8832
rect 13228 8780 13234 8832
rect 14826 8780 14832 8832
rect 14884 8820 14890 8832
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 14884 8792 15945 8820
rect 14884 8780 14890 8792
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 15933 8783 15991 8789
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16960 8820 16988 8919
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 17494 8916 17500 8968
rect 17552 8916 17558 8968
rect 17586 8916 17592 8968
rect 17644 8916 17650 8968
rect 16632 8792 16988 8820
rect 16632 8780 16638 8792
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 17586 8820 17592 8832
rect 17368 8792 17592 8820
rect 17368 8780 17374 8792
rect 17586 8780 17592 8792
rect 17644 8820 17650 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17644 8792 17785 8820
rect 17644 8780 17650 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17773 8783 17831 8789
rect 1104 8730 18492 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 18492 8730
rect 1104 8656 18492 8678
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4982 8616 4988 8628
rect 4212 8588 4988 8616
rect 4212 8576 4218 8588
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 8297 8619 8355 8625
rect 8297 8616 8309 8619
rect 5592 8588 8309 8616
rect 5592 8576 5598 8588
rect 8297 8585 8309 8588
rect 8343 8616 8355 8619
rect 8754 8616 8760 8628
rect 8343 8588 8760 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9364 8588 9505 8616
rect 9364 8576 9370 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 9916 8588 10517 8616
rect 9916 8576 9922 8588
rect 10505 8585 10517 8588
rect 10551 8616 10563 8619
rect 11146 8616 11152 8628
rect 10551 8588 11152 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 12529 8619 12587 8625
rect 12529 8585 12541 8619
rect 12575 8616 12587 8619
rect 12986 8616 12992 8628
rect 12575 8588 12992 8616
rect 12575 8585 12587 8588
rect 12529 8579 12587 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 14182 8576 14188 8628
rect 14240 8616 14246 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14240 8588 14565 8616
rect 14240 8576 14246 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14553 8579 14611 8585
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 15102 8616 15108 8628
rect 14792 8588 15108 8616
rect 14792 8576 14798 8588
rect 15102 8576 15108 8588
rect 15160 8616 15166 8628
rect 15565 8619 15623 8625
rect 15160 8588 15332 8616
rect 15160 8576 15166 8588
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 4264 8520 7021 8548
rect 4264 8492 4292 8520
rect 7009 8517 7021 8520
rect 7055 8548 7067 8551
rect 7098 8548 7104 8560
rect 7055 8520 7104 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 7837 8551 7895 8557
rect 7837 8548 7849 8551
rect 7340 8520 7849 8548
rect 7340 8508 7346 8520
rect 7837 8517 7849 8520
rect 7883 8517 7895 8551
rect 8386 8548 8392 8560
rect 7837 8511 7895 8517
rect 7944 8520 8392 8548
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 2038 8440 2044 8492
rect 2096 8440 2102 8492
rect 4246 8440 4252 8492
rect 4304 8440 4310 8492
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4618 8483 4676 8489
rect 4618 8449 4630 8483
rect 4664 8449 4676 8483
rect 4618 8443 4676 8449
rect 4062 8372 4068 8424
rect 4120 8372 4126 8424
rect 4632 8412 4660 8443
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5258 8480 5264 8492
rect 5031 8452 5264 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6420 8452 6561 8480
rect 6420 8440 6426 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 6914 8480 6920 8492
rect 6871 8452 6920 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 5166 8412 5172 8424
rect 4632 8384 5172 8412
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 6748 8412 6776 8443
rect 6914 8440 6920 8452
rect 6972 8480 6978 8492
rect 6972 8452 7604 8480
rect 6972 8440 6978 8452
rect 7576 8424 7604 8452
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 7944 8489 7972 8520
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 8938 8508 8944 8560
rect 8996 8508 9002 8560
rect 9030 8508 9036 8560
rect 9088 8508 9094 8560
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 9640 8520 9720 8548
rect 9640 8508 9646 8520
rect 8942 8505 9000 8508
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 7800 8452 7941 8480
rect 7800 8440 7806 8452
rect 7929 8449 7941 8452
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 8159 8452 8217 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8942 8471 8954 8505
rect 8988 8471 9000 8505
rect 8942 8465 9000 8471
rect 8205 8443 8263 8449
rect 6748 8384 6868 8412
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 1854 8304 1860 8356
rect 1912 8304 1918 8356
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 4706 8344 4712 8356
rect 4203 8316 4712 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4706 8304 4712 8316
rect 4764 8344 4770 8356
rect 4893 8347 4951 8353
rect 4893 8344 4905 8347
rect 4764 8316 4905 8344
rect 4764 8304 4770 8316
rect 4893 8313 4905 8316
rect 4939 8313 4951 8347
rect 4893 8307 4951 8313
rect 6362 8304 6368 8356
rect 6420 8304 6426 8356
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 4433 8279 4491 8285
rect 4433 8276 4445 8279
rect 3568 8248 4445 8276
rect 3568 8236 3574 8248
rect 4433 8245 4445 8248
rect 4479 8245 4491 8279
rect 4433 8239 4491 8245
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 5534 8276 5540 8288
rect 5040 8248 5540 8276
rect 5040 8236 5046 8248
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 6638 8276 6644 8288
rect 5960 8248 6644 8276
rect 5960 8236 5966 8248
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 6840 8276 6868 8384
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 8128 8412 8156 8443
rect 9122 8440 9128 8492
rect 9180 8440 9186 8492
rect 9692 8489 9720 8520
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 11572 8520 12449 8548
rect 11572 8508 11578 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 14752 8548 14780 8576
rect 12437 8511 12495 8517
rect 12544 8520 14780 8548
rect 14921 8551 14979 8557
rect 12544 8492 12572 8520
rect 14921 8517 14933 8551
rect 14967 8548 14979 8551
rect 15194 8548 15200 8560
rect 14967 8520 15200 8548
rect 14967 8517 14979 8520
rect 14921 8511 14979 8517
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 9243 8483 9301 8489
rect 9243 8449 9255 8483
rect 9289 8449 9301 8483
rect 9243 8443 9301 8449
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 7616 8384 8156 8412
rect 7616 8372 7622 8384
rect 8938 8372 8944 8424
rect 8996 8412 9002 8424
rect 9258 8412 9286 8443
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8480 10011 8483
rect 10042 8480 10048 8492
rect 9999 8452 10048 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 10502 8480 10508 8492
rect 10459 8452 10508 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 8996 8384 9286 8412
rect 9401 8415 9459 8421
rect 8996 8372 9002 8384
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 8110 8304 8116 8356
rect 8168 8304 8174 8356
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8386 8344 8392 8356
rect 8260 8316 8392 8344
rect 8260 8304 8266 8316
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 8628 8316 8769 8344
rect 8628 8304 8634 8316
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 9030 8304 9036 8356
rect 9088 8344 9094 8356
rect 9416 8344 9444 8375
rect 10137 8347 10195 8353
rect 10137 8344 10149 8347
rect 9088 8316 10149 8344
rect 9088 8304 9094 8316
rect 10137 8313 10149 8316
rect 10183 8313 10195 8347
rect 10137 8307 10195 8313
rect 10410 8304 10416 8356
rect 10468 8344 10474 8356
rect 10612 8344 10640 8443
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10744 8452 11069 8480
rect 10744 8440 10750 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11164 8412 11192 8443
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 11422 8440 11428 8492
rect 11480 8480 11486 8492
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11480 8452 11805 8480
rect 11480 8440 11486 8452
rect 11793 8449 11805 8452
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 11974 8440 11980 8492
rect 12032 8440 12038 8492
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8480 12219 8483
rect 12342 8480 12348 8492
rect 12207 8452 12348 8480
rect 12207 8449 12219 8452
rect 12161 8443 12219 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8480 13875 8483
rect 13906 8480 13912 8492
rect 13863 8452 13912 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 13078 8412 13084 8424
rect 11164 8384 13084 8412
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 14016 8412 14044 8443
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 14332 8452 14749 8480
rect 14332 8440 14338 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 14826 8440 14832 8492
rect 14884 8480 14890 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14884 8452 15025 8480
rect 14884 8440 14890 8452
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8480 15163 8483
rect 15304 8480 15332 8588
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15654 8616 15660 8628
rect 15611 8588 15660 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16206 8616 16212 8628
rect 15988 8588 16212 8616
rect 15988 8576 15994 8588
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16316 8588 16528 8616
rect 16025 8551 16083 8557
rect 16025 8517 16037 8551
rect 16071 8548 16083 8551
rect 16316 8548 16344 8588
rect 16071 8520 16344 8548
rect 16500 8548 16528 8588
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 17681 8619 17739 8625
rect 17681 8616 17693 8619
rect 16724 8588 16896 8616
rect 16724 8576 16730 8588
rect 16868 8557 16896 8588
rect 16960 8588 17693 8616
rect 16960 8557 16988 8588
rect 17681 8585 17693 8588
rect 17727 8585 17739 8619
rect 17681 8579 17739 8585
rect 16853 8551 16911 8557
rect 16500 8520 16804 8548
rect 16071 8517 16083 8520
rect 16025 8511 16083 8517
rect 15151 8452 15332 8480
rect 15151 8449 15163 8452
rect 15105 8443 15163 8449
rect 15562 8440 15568 8492
rect 15620 8440 15626 8492
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15804 8452 15945 8480
rect 15804 8440 15810 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 16574 8480 16580 8492
rect 16531 8452 16580 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 13596 8384 14044 8412
rect 13596 8372 13602 8384
rect 14366 8372 14372 8424
rect 14424 8412 14430 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 14424 8384 15393 8412
rect 14424 8372 14430 8384
rect 15381 8381 15393 8384
rect 15427 8412 15439 8415
rect 16022 8412 16028 8424
rect 15427 8384 16028 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 10468 8316 10640 8344
rect 11333 8347 11391 8353
rect 10468 8304 10474 8316
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 11606 8344 11612 8356
rect 11379 8316 11612 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11606 8304 11612 8316
rect 11664 8344 11670 8356
rect 12713 8347 12771 8353
rect 11664 8316 12296 8344
rect 11664 8304 11670 8316
rect 7282 8276 7288 8288
rect 6840 8248 7288 8276
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 8294 8276 8300 8288
rect 7800 8248 8300 8276
rect 7800 8236 7806 8248
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 11514 8236 11520 8288
rect 11572 8236 11578 8288
rect 12268 8276 12296 8316
rect 12713 8313 12725 8347
rect 12759 8313 12771 8347
rect 12713 8307 12771 8313
rect 12728 8276 12756 8307
rect 12894 8304 12900 8356
rect 12952 8304 12958 8356
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 13817 8347 13875 8353
rect 13817 8344 13829 8347
rect 13780 8316 13829 8344
rect 13780 8304 13786 8316
rect 13817 8313 13829 8316
rect 13863 8313 13875 8347
rect 13817 8307 13875 8313
rect 14550 8304 14556 8356
rect 14608 8344 14614 8356
rect 15654 8344 15660 8356
rect 14608 8316 15660 8344
rect 14608 8304 14614 8316
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 16132 8344 16160 8443
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 16776 8489 16804 8520
rect 16853 8517 16865 8551
rect 16899 8517 16911 8551
rect 16853 8511 16911 8517
rect 16945 8551 17003 8557
rect 16945 8517 16957 8551
rect 16991 8517 17003 8551
rect 16945 8511 17003 8517
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 17310 8440 17316 8492
rect 17368 8440 17374 8492
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 16666 8372 16672 8424
rect 16724 8372 16730 8424
rect 16850 8372 16856 8424
rect 16908 8372 16914 8424
rect 16868 8344 16896 8372
rect 16040 8316 16896 8344
rect 17420 8344 17448 8440
rect 17957 8347 18015 8353
rect 17957 8344 17969 8347
rect 17420 8316 17969 8344
rect 16040 8288 16068 8316
rect 17957 8313 17969 8316
rect 18003 8313 18015 8347
rect 17957 8307 18015 8313
rect 12268 8248 12756 8276
rect 15243 8279 15301 8285
rect 15243 8245 15255 8279
rect 15289 8276 15301 8279
rect 15378 8276 15384 8288
rect 15289 8248 15384 8276
rect 15289 8245 15301 8248
rect 15243 8239 15301 8245
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 16022 8236 16028 8288
rect 16080 8236 16086 8288
rect 16298 8236 16304 8288
rect 16356 8236 16362 8288
rect 16850 8236 16856 8288
rect 16908 8276 16914 8288
rect 17313 8279 17371 8285
rect 17313 8276 17325 8279
rect 16908 8248 17325 8276
rect 16908 8236 16914 8248
rect 17313 8245 17325 8248
rect 17359 8245 17371 8279
rect 17313 8239 17371 8245
rect 1104 8186 18492 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 18492 8186
rect 1104 8112 18492 8134
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 1670 8072 1676 8084
rect 1535 8044 1676 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 3694 8032 3700 8084
rect 3752 8072 3758 8084
rect 4982 8072 4988 8084
rect 3752 8044 4988 8072
rect 3752 8032 3758 8044
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5629 8075 5687 8081
rect 5629 8072 5641 8075
rect 5552 8044 5641 8072
rect 5552 8004 5580 8044
rect 5629 8041 5641 8044
rect 5675 8041 5687 8075
rect 5629 8035 5687 8041
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 8938 8072 8944 8084
rect 7147 8044 8944 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9582 8032 9588 8084
rect 9640 8032 9646 8084
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 10226 8072 10232 8084
rect 10183 8044 10232 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 10226 8032 10232 8044
rect 10284 8072 10290 8084
rect 11330 8072 11336 8084
rect 10284 8044 11336 8072
rect 10284 8032 10290 8044
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 11514 8081 11520 8084
rect 11471 8075 11520 8081
rect 11471 8041 11483 8075
rect 11517 8041 11520 8075
rect 11471 8035 11520 8041
rect 11514 8032 11520 8035
rect 11572 8032 11578 8084
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 12158 8072 12164 8084
rect 11756 8044 12164 8072
rect 11756 8032 11762 8044
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12406 8044 12848 8072
rect 7193 8007 7251 8013
rect 2148 7976 5580 8004
rect 5644 7976 7048 8004
rect 1946 7896 1952 7948
rect 2004 7896 2010 7948
rect 2148 7945 2176 7976
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7905 2191 7939
rect 4706 7936 4712 7948
rect 2133 7899 2191 7905
rect 4264 7908 4712 7936
rect 1762 7828 1768 7880
rect 1820 7868 1826 7880
rect 1857 7871 1915 7877
rect 1857 7868 1869 7871
rect 1820 7840 1869 7868
rect 1820 7828 1826 7840
rect 1857 7837 1869 7840
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 4264 7877 4292 7908
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5261 7939 5319 7945
rect 5261 7936 5273 7939
rect 4856 7908 5273 7936
rect 4856 7896 4862 7908
rect 5261 7905 5273 7908
rect 5307 7936 5319 7939
rect 5644 7936 5672 7976
rect 5307 7908 5672 7936
rect 5736 7908 5948 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3936 7840 4077 7868
rect 3936 7828 3942 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4338 7828 4344 7880
rect 4396 7828 4402 7880
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 4890 7868 4896 7880
rect 4479 7840 4896 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5074 7828 5080 7880
rect 5132 7828 5138 7880
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 5534 7828 5540 7880
rect 5592 7828 5598 7880
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 5736 7868 5764 7908
rect 5684 7840 5764 7868
rect 5684 7828 5690 7840
rect 5811 7828 5817 7880
rect 5869 7828 5875 7880
rect 5920 7877 5948 7908
rect 6086 7896 6092 7948
rect 6144 7896 6150 7948
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 6822 7936 6828 7948
rect 6328 7908 6593 7936
rect 6328 7896 6334 7908
rect 5906 7871 5964 7877
rect 5906 7837 5918 7871
rect 5952 7837 5964 7871
rect 5906 7831 5964 7837
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 3602 7760 3608 7812
rect 3660 7800 3666 7812
rect 6196 7800 6224 7831
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6565 7877 6593 7908
rect 6748 7908 6828 7936
rect 6748 7877 6776 7908
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7020 7936 7048 7976
rect 7193 7973 7205 8007
rect 7239 7973 7251 8007
rect 8481 8007 8539 8013
rect 7193 7967 7251 7973
rect 8122 7976 8432 8004
rect 7208 7936 7236 7967
rect 8122 7936 8150 7976
rect 7020 7908 7236 7936
rect 8036 7908 8150 7936
rect 8404 7936 8432 7976
rect 8481 7973 8493 8007
rect 8527 8004 8539 8007
rect 8662 8004 8668 8016
rect 8527 7976 8668 8004
rect 8527 7973 8539 7976
rect 8481 7967 8539 7973
rect 8662 7964 8668 7976
rect 8720 8004 8726 8016
rect 9309 8007 9367 8013
rect 9309 8004 9321 8007
rect 8720 7976 9321 8004
rect 8720 7964 8726 7976
rect 9309 7973 9321 7976
rect 9355 7973 9367 8007
rect 9309 7967 9367 7973
rect 9528 7976 9996 8004
rect 8757 7939 8815 7945
rect 8404 7908 8524 7936
rect 6550 7871 6608 7877
rect 6550 7837 6562 7871
rect 6596 7837 6608 7871
rect 6550 7831 6608 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6963 7871 7021 7877
rect 6963 7837 6975 7871
rect 7009 7868 7021 7871
rect 7098 7868 7104 7880
rect 7009 7840 7104 7868
rect 7009 7837 7021 7840
rect 6963 7831 7021 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 3660 7772 6224 7800
rect 3660 7760 3666 7772
rect 6822 7760 6828 7812
rect 6880 7760 6886 7812
rect 7208 7800 7236 7831
rect 7282 7830 7288 7882
rect 7340 7858 7346 7882
rect 7377 7871 7435 7877
rect 7377 7858 7389 7871
rect 7340 7837 7389 7858
rect 7423 7837 7435 7871
rect 7340 7831 7435 7837
rect 7340 7830 7420 7831
rect 7466 7830 7472 7882
rect 7524 7877 7530 7882
rect 7524 7831 7533 7877
rect 7524 7830 7530 7831
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 8036 7877 8064 7908
rect 8294 7877 8300 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7708 7840 7849 7868
rect 7708 7828 7714 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7837 8079 7871
rect 8275 7871 8300 7877
rect 8021 7831 8079 7837
rect 7742 7800 7748 7812
rect 7208 7772 7748 7800
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 8110 7806 8116 7858
rect 8168 7806 8174 7858
rect 8275 7837 8287 7871
rect 8275 7831 8300 7837
rect 8294 7828 8300 7831
rect 8352 7828 8358 7880
rect 8386 7828 8392 7880
rect 8444 7828 8450 7880
rect 8496 7868 8524 7908
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 9528 7936 9556 7976
rect 8803 7908 9556 7936
rect 9968 7936 9996 7976
rect 10778 7964 10784 8016
rect 10836 8004 10842 8016
rect 12406 8004 12434 8044
rect 10836 7976 12434 8004
rect 10836 7964 10842 7976
rect 12710 7964 12716 8016
rect 12768 7964 12774 8016
rect 12820 8004 12848 8044
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 12952 8044 15577 8072
rect 12952 8032 12958 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 17221 8075 17279 8081
rect 17221 8041 17233 8075
rect 17267 8072 17279 8075
rect 17494 8072 17500 8084
rect 17267 8044 17500 8072
rect 17267 8041 17279 8044
rect 17221 8035 17279 8041
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 14645 8007 14703 8013
rect 12820 7976 13860 8004
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 9968 7908 11621 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 11609 7905 11621 7908
rect 11655 7905 11667 7939
rect 11609 7899 11667 7905
rect 11698 7896 11704 7948
rect 11756 7896 11762 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11808 7908 11897 7936
rect 8573 7871 8631 7877
rect 8573 7868 8585 7871
rect 8496 7840 8585 7868
rect 8573 7837 8585 7840
rect 8619 7868 8631 7871
rect 8846 7868 8852 7880
rect 8619 7840 8852 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 9030 7868 9036 7880
rect 8987 7840 9036 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9490 7868 9496 7880
rect 9447 7840 9496 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9140 7800 9168 7831
rect 8956 7772 9168 7800
rect 9232 7800 9260 7831
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 10100 7840 10149 7868
rect 10100 7828 10106 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11808 7877 11836 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 12728 7936 12756 7964
rect 12897 7939 12955 7945
rect 12897 7936 12909 7939
rect 12728 7908 12909 7936
rect 11885 7899 11943 7905
rect 12897 7905 12909 7908
rect 12943 7905 12955 7939
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 12897 7899 12955 7905
rect 13004 7908 13277 7936
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11296 7840 11345 7868
rect 11296 7828 11302 7840
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 12066 7828 12072 7880
rect 12124 7828 12130 7880
rect 12158 7828 12164 7880
rect 12216 7828 12222 7880
rect 12250 7828 12256 7880
rect 12308 7828 12314 7880
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7837 12403 7871
rect 12345 7831 12403 7837
rect 10318 7800 10324 7812
rect 9232 7772 10324 7800
rect 8956 7744 8984 7772
rect 10318 7760 10324 7772
rect 10376 7800 10382 7812
rect 10686 7800 10692 7812
rect 10376 7772 10692 7800
rect 10376 7760 10382 7772
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 12360 7800 12388 7831
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 12710 7828 12716 7880
rect 12768 7828 12774 7880
rect 12802 7828 12808 7880
rect 12860 7828 12866 7880
rect 10928 7772 12388 7800
rect 10928 7760 10934 7772
rect 12894 7760 12900 7812
rect 12952 7800 12958 7812
rect 13004 7800 13032 7908
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 12952 7772 13032 7800
rect 12952 7760 12958 7772
rect 4706 7692 4712 7744
rect 4764 7692 4770 7744
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 4893 7735 4951 7741
rect 4893 7732 4905 7735
rect 4856 7704 4905 7732
rect 4856 7692 4862 7704
rect 4893 7701 4905 7704
rect 4939 7701 4951 7735
rect 4893 7695 4951 7701
rect 5166 7692 5172 7744
rect 5224 7732 5230 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 5224 7704 7573 7732
rect 5224 7692 5230 7704
rect 7561 7701 7573 7704
rect 7607 7732 7619 7735
rect 7650 7732 7656 7744
rect 7607 7704 7656 7732
rect 7607 7701 7619 7704
rect 7561 7695 7619 7701
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8202 7732 8208 7744
rect 8067 7704 8208 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 10410 7692 10416 7744
rect 10468 7732 10474 7744
rect 12158 7732 12164 7744
rect 10468 7704 12164 7732
rect 10468 7692 10474 7704
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 13096 7732 13124 7831
rect 12308 7704 13124 7732
rect 13464 7732 13492 7831
rect 13722 7828 13728 7880
rect 13780 7828 13786 7880
rect 13832 7868 13860 7976
rect 14645 7973 14657 8007
rect 14691 8004 14703 8007
rect 14691 7976 15148 8004
rect 14691 7973 14703 7976
rect 14645 7967 14703 7973
rect 13909 7939 13967 7945
rect 13909 7905 13921 7939
rect 13955 7936 13967 7939
rect 13955 7908 14504 7936
rect 13955 7905 13967 7908
rect 13909 7899 13967 7905
rect 14476 7877 14504 7908
rect 15010 7896 15016 7948
rect 15068 7896 15074 7948
rect 15120 7945 15148 7976
rect 15378 7964 15384 8016
rect 15436 8004 15442 8016
rect 16114 8004 16120 8016
rect 15436 7976 16120 8004
rect 15436 7964 15442 7976
rect 16114 7964 16120 7976
rect 16172 8004 16178 8016
rect 17405 8007 17463 8013
rect 17405 8004 17417 8007
rect 16172 7976 17417 8004
rect 16172 7964 16178 7976
rect 17405 7973 17417 7976
rect 17451 7973 17463 8007
rect 17405 7967 17463 7973
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7905 15163 7939
rect 15105 7899 15163 7905
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7936 15347 7939
rect 15749 7939 15807 7945
rect 15335 7908 15700 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13832 7840 14105 7868
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14826 7828 14832 7880
rect 14884 7828 14890 7880
rect 14918 7828 14924 7880
rect 14976 7828 14982 7880
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15028 7840 15577 7868
rect 15028 7812 15056 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15672 7868 15700 7908
rect 15749 7905 15761 7939
rect 15795 7936 15807 7939
rect 16666 7936 16672 7948
rect 15795 7908 16672 7936
rect 15795 7905 15807 7908
rect 15749 7899 15807 7905
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 15672 7840 17877 7868
rect 15565 7831 15623 7837
rect 17865 7837 17877 7840
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 13538 7760 13544 7812
rect 13596 7760 13602 7812
rect 13630 7760 13636 7812
rect 13688 7800 13694 7812
rect 14277 7803 14335 7809
rect 14277 7800 14289 7803
rect 13688 7772 14289 7800
rect 13688 7760 13694 7772
rect 14277 7769 14289 7772
rect 14323 7769 14335 7803
rect 14277 7763 14335 7769
rect 14366 7760 14372 7812
rect 14424 7760 14430 7812
rect 15010 7760 15016 7812
rect 15068 7760 15074 7812
rect 15838 7760 15844 7812
rect 15896 7760 15902 7812
rect 16298 7760 16304 7812
rect 16356 7800 16362 7812
rect 16850 7800 16856 7812
rect 16356 7772 16856 7800
rect 16356 7760 16362 7772
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 14734 7732 14740 7744
rect 13464 7704 14740 7732
rect 12308 7692 12314 7704
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 15378 7692 15384 7744
rect 15436 7692 15442 7744
rect 17126 7692 17132 7744
rect 17184 7732 17190 7744
rect 17230 7735 17288 7741
rect 17230 7732 17242 7735
rect 17184 7704 17242 7732
rect 17184 7692 17190 7704
rect 17230 7701 17242 7704
rect 17276 7732 17288 7735
rect 17586 7732 17592 7744
rect 17276 7704 17592 7732
rect 17276 7701 17288 7704
rect 17230 7695 17288 7701
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 18046 7692 18052 7744
rect 18104 7692 18110 7744
rect 1104 7642 18492 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 18492 7642
rect 1104 7568 18492 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 1949 7531 2007 7537
rect 1949 7528 1961 7531
rect 1820 7500 1961 7528
rect 1820 7488 1826 7500
rect 1949 7497 1961 7500
rect 1995 7497 2007 7531
rect 3418 7528 3424 7540
rect 1949 7491 2007 7497
rect 2424 7500 3424 7528
rect 2424 7469 2452 7500
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 4430 7528 4436 7540
rect 3844 7500 4436 7528
rect 3844 7488 3850 7500
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 5261 7531 5319 7537
rect 5261 7528 5273 7531
rect 4632 7500 5273 7528
rect 2409 7463 2467 7469
rect 2409 7429 2421 7463
rect 2455 7429 2467 7463
rect 3881 7463 3939 7469
rect 3881 7460 3893 7463
rect 2409 7423 2467 7429
rect 2976 7432 3893 7460
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 1946 7392 1952 7404
rect 1903 7364 1952 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2590 7352 2596 7404
rect 2648 7352 2654 7404
rect 2694 7398 2752 7401
rect 2866 7398 2872 7404
rect 2694 7395 2872 7398
rect 2694 7361 2706 7395
rect 2740 7370 2872 7395
rect 2740 7364 2774 7370
rect 2740 7361 2752 7364
rect 2694 7355 2752 7361
rect 2866 7352 2872 7370
rect 2924 7352 2930 7404
rect 2976 7401 3004 7432
rect 3881 7429 3893 7432
rect 3927 7429 3939 7463
rect 3881 7423 3939 7429
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3050 7352 3056 7404
rect 3108 7352 3114 7404
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3326 7352 3332 7404
rect 3384 7352 3390 7404
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7293 2191 7327
rect 2133 7287 2191 7293
rect 2148 7256 2176 7287
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 4249 7327 4307 7333
rect 4249 7324 4261 7327
rect 3568 7296 4261 7324
rect 3568 7284 3574 7296
rect 4249 7293 4261 7296
rect 4295 7293 4307 7327
rect 4356 7324 4384 7355
rect 4430 7352 4436 7404
rect 4488 7398 4494 7404
rect 4525 7398 4583 7401
rect 4488 7395 4583 7398
rect 4488 7370 4537 7395
rect 4488 7352 4494 7370
rect 4525 7361 4537 7370
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 4632 7324 4660 7500
rect 5261 7497 5273 7500
rect 5307 7497 5319 7531
rect 5261 7491 5319 7497
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 5994 7528 6000 7540
rect 5500 7500 6000 7528
rect 5500 7488 5506 7500
rect 5994 7488 6000 7500
rect 6052 7528 6058 7540
rect 6822 7528 6828 7540
rect 6052 7500 6828 7528
rect 6052 7488 6058 7500
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 9950 7528 9956 7540
rect 7340 7500 9956 7528
rect 7340 7488 7346 7500
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 11790 7528 11796 7540
rect 10284 7500 11796 7528
rect 10284 7488 10290 7500
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 13630 7488 13636 7540
rect 13688 7488 13694 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 14366 7528 14372 7540
rect 13872 7500 14372 7528
rect 13872 7488 13878 7500
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 14826 7488 14832 7540
rect 14884 7528 14890 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14884 7500 15025 7528
rect 14884 7488 14890 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 15194 7488 15200 7540
rect 15252 7488 15258 7540
rect 15378 7488 15384 7540
rect 15436 7488 15442 7540
rect 4908 7432 5396 7460
rect 4908 7401 4936 7432
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 4356 7296 4660 7324
rect 4816 7324 4844 7355
rect 5074 7352 5080 7404
rect 5132 7352 5138 7404
rect 5166 7352 5172 7404
rect 5224 7352 5230 7404
rect 5258 7324 5264 7336
rect 4816 7296 5264 7324
rect 4249 7287 4307 7293
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 5368 7324 5396 7432
rect 5460 7432 5856 7460
rect 5460 7401 5488 7432
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 5718 7352 5724 7404
rect 5776 7352 5782 7404
rect 5828 7392 5856 7432
rect 6086 7420 6092 7472
rect 6144 7460 6150 7472
rect 10391 7463 10449 7469
rect 10391 7460 10403 7463
rect 6144 7432 10403 7460
rect 6144 7420 6150 7432
rect 10391 7429 10403 7432
rect 10437 7429 10449 7463
rect 10391 7423 10449 7429
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 12526 7460 12532 7472
rect 10560 7432 12532 7460
rect 10560 7420 10566 7432
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 15396 7460 15424 7488
rect 12952 7432 13308 7460
rect 12952 7420 12958 7432
rect 6270 7392 6276 7404
rect 5828 7364 6276 7392
rect 6270 7352 6276 7364
rect 6328 7392 6334 7404
rect 8754 7392 8760 7404
rect 6328 7364 8760 7392
rect 6328 7352 6334 7364
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 10042 7392 10048 7404
rect 9088 7364 10048 7392
rect 9088 7352 9094 7364
rect 10042 7352 10048 7364
rect 10100 7392 10106 7404
rect 10520 7392 10548 7420
rect 10100 7364 10548 7392
rect 10689 7395 10747 7401
rect 10100 7352 10106 7364
rect 10689 7361 10701 7395
rect 10735 7392 10747 7395
rect 11238 7392 11244 7404
rect 10735 7364 11244 7392
rect 10735 7361 10747 7364
rect 10689 7355 10747 7361
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 13280 7401 13308 7432
rect 14384 7432 15424 7460
rect 14384 7401 14412 7432
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 14369 7395 14427 7401
rect 14369 7361 14381 7395
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 7558 7324 7564 7336
rect 5368 7296 7564 7324
rect 7558 7284 7564 7296
rect 7616 7324 7622 7336
rect 7616 7296 8294 7324
rect 7616 7284 7622 7296
rect 2777 7259 2835 7265
rect 2777 7256 2789 7259
rect 2148 7228 2789 7256
rect 2777 7225 2789 7228
rect 2823 7225 2835 7259
rect 2777 7219 2835 7225
rect 4157 7259 4215 7265
rect 4157 7225 4169 7259
rect 4203 7256 4215 7259
rect 6454 7256 6460 7268
rect 4203 7228 6460 7256
rect 4203 7225 4215 7228
rect 4157 7219 4215 7225
rect 6454 7216 6460 7228
rect 6512 7216 6518 7268
rect 8266 7256 8294 7296
rect 10134 7284 10140 7336
rect 10192 7324 10198 7336
rect 10505 7327 10563 7333
rect 10505 7324 10517 7327
rect 10192 7296 10517 7324
rect 10192 7284 10198 7296
rect 10505 7293 10517 7296
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 10226 7256 10232 7268
rect 8266 7228 10232 7256
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 10321 7259 10379 7265
rect 10321 7225 10333 7259
rect 10367 7256 10379 7259
rect 10686 7256 10692 7268
rect 10367 7228 10692 7256
rect 10367 7225 10379 7228
rect 10321 7219 10379 7225
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 13372 7200 13400 7287
rect 13538 7284 13544 7336
rect 13596 7324 13602 7336
rect 14568 7324 14596 7355
rect 13596 7296 14596 7324
rect 13596 7284 13602 7296
rect 14550 7216 14556 7268
rect 14608 7256 14614 7268
rect 14645 7259 14703 7265
rect 14645 7256 14657 7259
rect 14608 7228 14657 7256
rect 14608 7216 14614 7228
rect 14645 7225 14657 7228
rect 14691 7225 14703 7259
rect 14645 7219 14703 7225
rect 14734 7216 14740 7268
rect 14792 7216 14798 7268
rect 14844 7256 14872 7355
rect 15212 7324 15240 7355
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 15381 7395 15439 7401
rect 15381 7392 15393 7395
rect 15344 7364 15393 7392
rect 15344 7352 15350 7364
rect 15381 7361 15393 7364
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15930 7324 15936 7336
rect 15212 7296 15936 7324
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 15562 7256 15568 7268
rect 14844 7228 15568 7256
rect 1489 7191 1547 7197
rect 1489 7157 1501 7191
rect 1535 7188 1547 7191
rect 1670 7188 1676 7200
rect 1535 7160 1676 7188
rect 1535 7157 1547 7160
rect 1489 7151 1547 7157
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 2409 7191 2467 7197
rect 2409 7157 2421 7191
rect 2455 7188 2467 7191
rect 2498 7188 2504 7200
rect 2455 7160 2504 7188
rect 2455 7157 2467 7160
rect 2409 7151 2467 7157
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 3878 7148 3884 7200
rect 3936 7188 3942 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 3936 7160 4629 7188
rect 3936 7148 3942 7160
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 4617 7151 4675 7157
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 5534 7188 5540 7200
rect 4856 7160 5540 7188
rect 4856 7148 4862 7160
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 9030 7188 9036 7200
rect 7708 7160 9036 7188
rect 7708 7148 7714 7160
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10502 7188 10508 7200
rect 10008 7160 10508 7188
rect 10008 7148 10014 7160
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 10962 7188 10968 7200
rect 10643 7160 10968 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 13262 7148 13268 7200
rect 13320 7148 13326 7200
rect 13354 7148 13360 7200
rect 13412 7188 13418 7200
rect 14844 7188 14872 7228
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 13412 7160 14872 7188
rect 13412 7148 13418 7160
rect 1104 7098 18492 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 18492 7098
rect 1104 7024 18492 7046
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 4433 6987 4491 6993
rect 4433 6984 4445 6987
rect 3384 6956 4445 6984
rect 3384 6944 3390 6956
rect 4433 6953 4445 6956
rect 4479 6953 4491 6987
rect 4433 6947 4491 6953
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6178 6984 6184 6996
rect 5592 6956 6184 6984
rect 5592 6944 5598 6956
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 6641 6987 6699 6993
rect 6641 6953 6653 6987
rect 6687 6984 6699 6987
rect 7374 6984 7380 6996
rect 6687 6956 7380 6984
rect 6687 6953 6699 6956
rect 6641 6947 6699 6953
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 9493 6987 9551 6993
rect 9493 6953 9505 6987
rect 9539 6984 9551 6987
rect 9674 6984 9680 6996
rect 9539 6956 9680 6984
rect 9539 6953 9551 6956
rect 9493 6947 9551 6953
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 9953 6987 10011 6993
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10229 6987 10287 6993
rect 10229 6984 10241 6987
rect 9999 6956 10241 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10229 6953 10241 6956
rect 10275 6953 10287 6987
rect 10229 6947 10287 6953
rect 10686 6944 10692 6996
rect 10744 6944 10750 6996
rect 10962 6944 10968 6996
rect 11020 6944 11026 6996
rect 11054 6944 11060 6996
rect 11112 6984 11118 6996
rect 11112 6956 11284 6984
rect 11112 6944 11118 6956
rect 10410 6916 10416 6928
rect 9876 6888 10180 6916
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 3142 6848 3148 6860
rect 2639 6820 3148 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 4522 6808 4528 6860
rect 4580 6848 4586 6860
rect 4709 6851 4767 6857
rect 4709 6848 4721 6851
rect 4580 6820 4721 6848
rect 4580 6808 4586 6820
rect 4709 6817 4721 6820
rect 4755 6817 4767 6851
rect 4709 6811 4767 6817
rect 4893 6851 4951 6857
rect 4893 6817 4905 6851
rect 4939 6848 4951 6851
rect 5169 6851 5227 6857
rect 5169 6848 5181 6851
rect 4939 6820 5181 6848
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 5169 6817 5181 6820
rect 5215 6817 5227 6851
rect 5169 6811 5227 6817
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5718 6848 5724 6860
rect 5399 6820 5724 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 9766 6848 9772 6860
rect 8260 6820 9772 6848
rect 8260 6808 8266 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 1670 6740 1676 6792
rect 1728 6740 1734 6792
rect 2498 6740 2504 6792
rect 2556 6740 2562 6792
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 3786 6780 3792 6792
rect 2731 6752 3792 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4080 6712 4108 6743
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 4338 6740 4344 6792
rect 4396 6740 4402 6792
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 4801 6783 4859 6789
rect 4663 6752 4752 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 4724 6724 4752 6752
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 4430 6712 4436 6724
rect 4080 6684 4436 6712
rect 4430 6672 4436 6684
rect 4488 6672 4494 6724
rect 4706 6672 4712 6724
rect 4764 6672 4770 6724
rect 4816 6712 4844 6743
rect 4982 6740 4988 6792
rect 5040 6780 5046 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 5040 6752 5089 6780
rect 5040 6740 5046 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5258 6740 5264 6792
rect 5316 6780 5322 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5316 6752 5457 6780
rect 5316 6740 5322 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 5626 6740 5632 6792
rect 5684 6740 5690 6792
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6822 6780 6828 6792
rect 6052 6752 6828 6780
rect 6052 6740 6058 6752
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7466 6780 7472 6792
rect 7147 6752 7472 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8294 6780 8300 6792
rect 7984 6752 8300 6780
rect 7984 6740 7990 6752
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9876 6780 9904 6888
rect 10152 6789 10180 6888
rect 10336 6888 10416 6916
rect 10336 6789 10364 6888
rect 10410 6876 10416 6888
rect 10468 6876 10474 6928
rect 11256 6856 11284 6956
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13446 6984 13452 6996
rect 13136 6956 13452 6984
rect 13136 6944 13142 6956
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 11422 6876 11428 6928
rect 11480 6916 11486 6928
rect 13538 6916 13544 6928
rect 11480 6888 13544 6916
rect 11480 6876 11486 6888
rect 13538 6876 13544 6888
rect 13596 6876 13602 6928
rect 13998 6876 14004 6928
rect 14056 6916 14062 6928
rect 14056 6888 15148 6916
rect 14056 6876 14062 6888
rect 11333 6856 11391 6857
rect 11256 6851 11391 6856
rect 11256 6828 11345 6851
rect 11333 6817 11345 6828
rect 11379 6817 11391 6851
rect 11333 6811 11391 6817
rect 14366 6808 14372 6860
rect 14424 6848 14430 6860
rect 15010 6848 15016 6860
rect 14424 6820 15016 6848
rect 14424 6808 14430 6820
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15120 6848 15148 6888
rect 15194 6876 15200 6928
rect 15252 6916 15258 6928
rect 15252 6888 15700 6916
rect 15252 6876 15258 6888
rect 15672 6857 15700 6888
rect 16482 6876 16488 6928
rect 16540 6876 16546 6928
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15120 6820 15577 6848
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6817 15715 6851
rect 16500 6848 16528 6876
rect 17402 6848 17408 6860
rect 15657 6811 15715 6817
rect 15764 6820 17408 6848
rect 9548 6752 9904 6780
rect 10045 6783 10103 6789
rect 9548 6740 9554 6752
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 9582 6712 9588 6724
rect 4816 6684 9588 6712
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 9677 6715 9735 6721
rect 9677 6681 9689 6715
rect 9723 6712 9735 6715
rect 10060 6712 10088 6743
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 11054 6780 11060 6792
rect 10735 6752 11060 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 10226 6712 10232 6724
rect 9723 6684 9996 6712
rect 10060 6684 10232 6712
rect 9723 6681 9735 6684
rect 9677 6675 9735 6681
rect 9968 6656 9996 6684
rect 10226 6672 10232 6684
rect 10284 6672 10290 6724
rect 10962 6672 10968 6724
rect 11020 6712 11026 6724
rect 11164 6712 11192 6743
rect 11238 6740 11244 6792
rect 11296 6740 11302 6792
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11020 6684 11192 6712
rect 11440 6712 11468 6743
rect 11606 6740 11612 6792
rect 11664 6740 11670 6792
rect 14918 6789 14924 6792
rect 14916 6780 14924 6789
rect 14879 6752 14924 6780
rect 14916 6743 14924 6752
rect 14918 6740 14924 6743
rect 14976 6740 14982 6792
rect 15028 6780 15056 6808
rect 15233 6783 15291 6789
rect 15233 6780 15245 6783
rect 15028 6752 15245 6780
rect 15233 6749 15245 6752
rect 15279 6749 15291 6783
rect 15233 6743 15291 6749
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6780 15439 6783
rect 15470 6780 15476 6792
rect 15427 6752 15476 6780
rect 15427 6749 15439 6752
rect 15381 6743 15439 6749
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 15580 6780 15608 6811
rect 15764 6780 15792 6820
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 15580 6752 15792 6780
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 12894 6712 12900 6724
rect 11440 6684 12900 6712
rect 11020 6672 11026 6684
rect 12894 6672 12900 6684
rect 12952 6672 12958 6724
rect 15013 6715 15071 6721
rect 15013 6681 15025 6715
rect 15059 6681 15071 6715
rect 15013 6675 15071 6681
rect 842 6604 848 6656
rect 900 6644 906 6656
rect 1489 6647 1547 6653
rect 1489 6644 1501 6647
rect 900 6616 1501 6644
rect 900 6604 906 6616
rect 1489 6613 1501 6616
rect 1535 6613 1547 6647
rect 1489 6607 1547 6613
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 6914 6644 6920 6656
rect 3108 6616 6920 6644
rect 3108 6604 3114 6616
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7009 6647 7067 6653
rect 7009 6613 7021 6647
rect 7055 6644 7067 6647
rect 7282 6644 7288 6656
rect 7055 6616 7288 6644
rect 7055 6613 7067 6616
rect 7009 6607 7067 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 9306 6604 9312 6656
rect 9364 6604 9370 6656
rect 9477 6647 9535 6653
rect 9477 6613 9489 6647
rect 9523 6644 9535 6647
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 9523 6616 9781 6644
rect 9523 6613 9535 6616
rect 9477 6607 9535 6613
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 9950 6604 9956 6656
rect 10008 6604 10014 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 13354 6644 13360 6656
rect 11664 6616 13360 6644
rect 11664 6604 11670 6616
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14737 6647 14795 6653
rect 14737 6644 14749 6647
rect 14608 6616 14749 6644
rect 14608 6604 14614 6616
rect 14737 6613 14749 6616
rect 14783 6613 14795 6647
rect 15028 6644 15056 6675
rect 15102 6672 15108 6724
rect 15160 6672 15166 6724
rect 15746 6672 15752 6724
rect 15804 6712 15810 6724
rect 15856 6712 15884 6743
rect 15930 6740 15936 6792
rect 15988 6740 15994 6792
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16485 6783 16543 6789
rect 16485 6780 16497 6783
rect 16448 6752 16497 6780
rect 16448 6740 16454 6752
rect 16485 6749 16497 6752
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6780 16911 6783
rect 16942 6780 16948 6792
rect 16899 6752 16948 6780
rect 16899 6749 16911 6752
rect 16853 6743 16911 6749
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17034 6740 17040 6792
rect 17092 6740 17098 6792
rect 15804 6684 15884 6712
rect 15804 6672 15810 6684
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 15028 6616 15485 6644
rect 14737 6607 14795 6613
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15948 6644 15976 6740
rect 16390 6644 16396 6656
rect 15948 6616 16396 6644
rect 15473 6607 15531 6613
rect 16390 6604 16396 6616
rect 16448 6644 16454 6656
rect 16669 6647 16727 6653
rect 16669 6644 16681 6647
rect 16448 6616 16681 6644
rect 16448 6604 16454 6616
rect 16669 6613 16681 6616
rect 16715 6613 16727 6647
rect 16669 6607 16727 6613
rect 17037 6647 17095 6653
rect 17037 6613 17049 6647
rect 17083 6644 17095 6647
rect 17586 6644 17592 6656
rect 17083 6616 17592 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 17586 6604 17592 6616
rect 17644 6604 17650 6656
rect 1104 6554 18492 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 18492 6554
rect 1104 6480 18492 6502
rect 2314 6440 2320 6452
rect 1688 6412 2320 6440
rect 1688 6381 1716 6412
rect 2314 6400 2320 6412
rect 2372 6400 2378 6452
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 3050 6440 3056 6452
rect 2464 6412 3056 6440
rect 2464 6400 2470 6412
rect 1673 6375 1731 6381
rect 1673 6341 1685 6375
rect 1719 6341 1731 6375
rect 1673 6335 1731 6341
rect 1857 6375 1915 6381
rect 1857 6341 1869 6375
rect 1903 6372 1915 6375
rect 1903 6344 2452 6372
rect 1903 6341 1915 6344
rect 1857 6335 1915 6341
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1964 6168 1992 6267
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2424 6313 2452 6344
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6273 2467 6307
rect 2409 6267 2467 6273
rect 2424 6236 2452 6267
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 2700 6313 2728 6412
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 5902 6400 5908 6452
rect 5960 6400 5966 6452
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 6546 6440 6552 6452
rect 6104 6412 6552 6440
rect 2774 6332 2780 6384
rect 2832 6372 2838 6384
rect 3145 6375 3203 6381
rect 3145 6372 3157 6375
rect 2832 6344 3157 6372
rect 2832 6332 2838 6344
rect 3145 6341 3157 6344
rect 3191 6372 3203 6375
rect 3865 6375 3923 6381
rect 3191 6344 3832 6372
rect 3191 6341 3203 6344
rect 3145 6335 3203 6341
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6273 2743 6307
rect 2685 6267 2743 6273
rect 2958 6264 2964 6316
rect 3016 6264 3022 6316
rect 3234 6264 3240 6316
rect 3292 6264 3298 6316
rect 3804 6304 3832 6344
rect 3865 6341 3877 6375
rect 3911 6372 3923 6375
rect 3911 6344 4016 6372
rect 3911 6341 3923 6344
rect 3865 6335 3923 6341
rect 3988 6304 4016 6344
rect 4062 6332 4068 6384
rect 4120 6332 4126 6384
rect 5718 6304 5724 6316
rect 3804 6276 3924 6304
rect 3988 6276 5724 6304
rect 3896 6236 3924 6276
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 5920 6304 6040 6307
rect 6104 6304 6132 6412
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 6972 6412 8708 6440
rect 6972 6400 6978 6412
rect 8110 6372 8116 6384
rect 6196 6344 8116 6372
rect 6196 6313 6224 6344
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 8478 6332 8484 6384
rect 8536 6381 8542 6384
rect 8680 6381 8708 6412
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9122 6440 9128 6452
rect 8812 6412 9128 6440
rect 8812 6400 8818 6412
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 11707 6443 11765 6449
rect 11707 6440 11719 6443
rect 9640 6412 11719 6440
rect 9640 6400 9646 6412
rect 11707 6409 11719 6412
rect 11753 6440 11765 6443
rect 13722 6440 13728 6452
rect 11753 6412 12940 6440
rect 11753 6409 11765 6412
rect 11707 6403 11765 6409
rect 8536 6375 8585 6381
rect 8536 6341 8539 6375
rect 8573 6341 8585 6375
rect 8536 6335 8585 6341
rect 8665 6375 8723 6381
rect 8665 6341 8677 6375
rect 8711 6372 8723 6375
rect 8938 6372 8944 6384
rect 8711 6344 8944 6372
rect 8711 6341 8723 6344
rect 8665 6335 8723 6341
rect 8536 6332 8542 6335
rect 8938 6332 8944 6344
rect 8996 6332 9002 6384
rect 10134 6332 10140 6384
rect 10192 6372 10198 6384
rect 11422 6372 11428 6384
rect 10192 6344 11428 6372
rect 10192 6332 10198 6344
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 11514 6332 11520 6384
rect 11572 6372 11578 6384
rect 11609 6375 11667 6381
rect 11609 6372 11621 6375
rect 11572 6344 11621 6372
rect 11572 6332 11578 6344
rect 11609 6341 11621 6344
rect 11655 6341 11667 6375
rect 12912 6372 12940 6412
rect 13096 6412 13728 6440
rect 12912 6344 13032 6372
rect 11609 6335 11667 6341
rect 5859 6279 6132 6304
rect 5859 6276 5948 6279
rect 6012 6276 6132 6279
rect 6181 6307 6239 6313
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6181 6273 6193 6307
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7098 6304 7104 6316
rect 6972 6276 7104 6304
rect 6972 6264 6978 6276
rect 7098 6264 7104 6276
rect 7156 6304 7162 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7156 6276 7481 6304
rect 7156 6264 7162 6276
rect 7469 6273 7481 6276
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 9030 6304 9036 6316
rect 8895 6276 9036 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 8389 6239 8447 6245
rect 2424 6208 3740 6236
rect 3896 6208 5764 6236
rect 3712 6177 3740 6208
rect 2777 6171 2835 6177
rect 2777 6168 2789 6171
rect 1964 6140 2789 6168
rect 2777 6137 2789 6140
rect 2823 6137 2835 6171
rect 2777 6131 2835 6137
rect 3697 6171 3755 6177
rect 3697 6137 3709 6171
rect 3743 6137 3755 6171
rect 5626 6168 5632 6180
rect 3697 6131 3755 6137
rect 3804 6140 5632 6168
rect 1670 6060 1676 6112
rect 1728 6060 1734 6112
rect 1946 6060 1952 6112
rect 2004 6100 2010 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 2004 6072 2053 6100
rect 2004 6060 2010 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2041 6063 2099 6069
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3804 6100 3832 6140
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 5736 6168 5764 6208
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8938 6236 8944 6248
rect 8435 6208 8944 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 9416 6236 9444 6267
rect 9490 6264 9496 6316
rect 9548 6264 9554 6316
rect 9582 6264 9588 6316
rect 9640 6264 9646 6316
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 9815 6276 11284 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 10778 6236 10784 6248
rect 9180 6208 10784 6236
rect 9180 6196 9186 6208
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 11256 6236 11284 6276
rect 11330 6264 11336 6316
rect 11388 6304 11394 6316
rect 11793 6307 11851 6313
rect 11793 6304 11805 6307
rect 11388 6276 11805 6304
rect 11388 6264 11394 6276
rect 11793 6273 11805 6276
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 12250 6304 12256 6316
rect 11940 6276 12256 6304
rect 11940 6264 11946 6276
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6273 12863 6307
rect 12805 6267 12863 6273
rect 11606 6236 11612 6248
rect 11256 6208 11612 6236
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 5905 6171 5963 6177
rect 5905 6168 5917 6171
rect 5736 6140 5917 6168
rect 5905 6137 5917 6140
rect 5951 6137 5963 6171
rect 5905 6131 5963 6137
rect 7466 6128 7472 6180
rect 7524 6168 7530 6180
rect 7653 6171 7711 6177
rect 7653 6168 7665 6171
rect 7524 6140 7665 6168
rect 7524 6128 7530 6140
rect 7653 6137 7665 6140
rect 7699 6137 7711 6171
rect 7653 6131 7711 6137
rect 7834 6128 7840 6180
rect 7892 6168 7898 6180
rect 12820 6168 12848 6267
rect 12894 6264 12900 6316
rect 12952 6264 12958 6316
rect 13004 6313 13032 6344
rect 13096 6313 13124 6412
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 15102 6400 15108 6452
rect 15160 6440 15166 6452
rect 15657 6443 15715 6449
rect 15657 6440 15669 6443
rect 15160 6412 15669 6440
rect 15160 6400 15166 6412
rect 15657 6409 15669 6412
rect 15703 6409 15715 6443
rect 17034 6440 17040 6452
rect 15657 6403 15715 6409
rect 16316 6412 17040 6440
rect 14090 6372 14096 6384
rect 13556 6344 14096 6372
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13262 6264 13268 6316
rect 13320 6264 13326 6316
rect 13556 6313 13584 6344
rect 14090 6332 14096 6344
rect 14148 6372 14154 6384
rect 16316 6372 16344 6412
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6409 17279 6443
rect 17221 6403 17279 6409
rect 14148 6344 16344 6372
rect 14148 6332 14154 6344
rect 16390 6332 16396 6384
rect 16448 6372 16454 6384
rect 16448 6344 16712 6372
rect 16448 6332 16454 6344
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6273 13599 6307
rect 16206 6304 16212 6316
rect 13541 6267 13599 6273
rect 13832 6276 16212 6304
rect 12912 6236 12940 6264
rect 13357 6239 13415 6245
rect 13357 6236 13369 6239
rect 12912 6208 13369 6236
rect 13357 6205 13369 6208
rect 13403 6205 13415 6239
rect 13357 6199 13415 6205
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13504 6208 13645 6236
rect 13504 6196 13510 6208
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 13633 6199 13691 6205
rect 13722 6196 13728 6248
rect 13780 6196 13786 6248
rect 13832 6245 13860 6276
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 16298 6264 16304 6316
rect 16356 6264 16362 6316
rect 16482 6264 16488 6316
rect 16540 6264 16546 6316
rect 16684 6313 16712 6344
rect 16850 6332 16856 6384
rect 16908 6332 16914 6384
rect 17052 6313 17080 6400
rect 17236 6372 17264 6403
rect 17236 6344 17724 6372
rect 16669 6307 16727 6313
rect 16669 6273 16681 6307
rect 16715 6273 16727 6307
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 16669 6267 16727 6273
rect 16868 6276 16957 6304
rect 16868 6248 16896 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 17310 6264 17316 6316
rect 17368 6264 17374 6316
rect 17402 6264 17408 6316
rect 17460 6264 17466 6316
rect 17586 6264 17592 6316
rect 17644 6264 17650 6316
rect 17696 6313 17724 6344
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 15804 6208 15853 6236
rect 15804 6196 15810 6208
rect 15841 6205 15853 6208
rect 15887 6205 15899 6239
rect 15841 6199 15899 6205
rect 15933 6239 15991 6245
rect 15933 6205 15945 6239
rect 15979 6205 15991 6239
rect 15933 6199 15991 6205
rect 15948 6168 15976 6199
rect 16022 6196 16028 6248
rect 16080 6196 16086 6248
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6236 16175 6239
rect 16393 6239 16451 6245
rect 16393 6236 16405 6239
rect 16163 6208 16405 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 16393 6205 16405 6208
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 16850 6196 16856 6248
rect 16908 6196 16914 6248
rect 16206 6168 16212 6180
rect 7892 6140 9260 6168
rect 12820 6140 13676 6168
rect 15948 6140 16212 6168
rect 7892 6128 7898 6140
rect 3016 6072 3832 6100
rect 3016 6060 3022 6072
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 9030 6060 9036 6112
rect 9088 6060 9094 6112
rect 9122 6060 9128 6112
rect 9180 6060 9186 6112
rect 9232 6100 9260 6140
rect 13648 6112 13676 6140
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 10686 6100 10692 6112
rect 9232 6072 10692 6100
rect 10686 6060 10692 6072
rect 10744 6100 10750 6112
rect 10870 6100 10876 6112
rect 10744 6072 10876 6100
rect 10744 6060 10750 6072
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 17865 6103 17923 6109
rect 17865 6100 17877 6103
rect 13688 6072 17877 6100
rect 13688 6060 13694 6072
rect 17865 6069 17877 6072
rect 17911 6069 17923 6103
rect 17865 6063 17923 6069
rect 1104 6010 18492 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 18492 6010
rect 1104 5936 18492 5958
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 2038 5896 2044 5908
rect 1995 5868 2044 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2498 5896 2504 5908
rect 2455 5868 2504 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 3053 5899 3111 5905
rect 3053 5865 3065 5899
rect 3099 5896 3111 5899
rect 3234 5896 3240 5908
rect 3099 5868 3240 5896
rect 3099 5865 3111 5868
rect 3053 5859 3111 5865
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 4338 5896 4344 5908
rect 3384 5868 4344 5896
rect 3384 5856 3390 5868
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 4672 5868 5212 5896
rect 4672 5856 4678 5868
rect 3510 5788 3516 5840
rect 3568 5828 3574 5840
rect 3568 5800 4108 5828
rect 3568 5788 3574 5800
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 2884 5732 3801 5760
rect 1670 5652 1676 5704
rect 1728 5652 1734 5704
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5692 1823 5695
rect 1854 5692 1860 5704
rect 1811 5664 1860 5692
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 1854 5652 1860 5664
rect 1912 5652 1918 5704
rect 1946 5652 1952 5704
rect 2004 5652 2010 5704
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2682 5692 2688 5704
rect 2639 5664 2688 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2774 5652 2780 5704
rect 2832 5652 2838 5704
rect 2884 5701 2912 5732
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 3789 5723 3847 5729
rect 3878 5720 3884 5772
rect 3936 5760 3942 5772
rect 3973 5763 4031 5769
rect 3973 5760 3985 5763
rect 3936 5732 3985 5760
rect 3936 5720 3942 5732
rect 3973 5729 3985 5732
rect 4019 5729 4031 5763
rect 4080 5760 4108 5800
rect 4798 5788 4804 5840
rect 4856 5788 4862 5840
rect 5184 5828 5212 5868
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 8478 5896 8484 5908
rect 5684 5868 8484 5896
rect 5684 5856 5690 5868
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 8665 5899 8723 5905
rect 8665 5865 8677 5899
rect 8711 5896 8723 5899
rect 8754 5896 8760 5908
rect 8711 5868 8760 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 9582 5896 9588 5908
rect 9048 5868 9588 5896
rect 6914 5828 6920 5840
rect 5184 5800 6920 5828
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 4080 5732 4261 5760
rect 3973 5723 4031 5729
rect 4249 5729 4261 5732
rect 4295 5760 4307 5763
rect 4816 5760 4844 5788
rect 5184 5760 5212 5800
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 7101 5831 7159 5837
rect 7101 5797 7113 5831
rect 7147 5828 7159 5831
rect 9048 5828 9076 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 10502 5856 10508 5908
rect 10560 5896 10566 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 10560 5868 11069 5896
rect 10560 5856 10566 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 13262 5856 13268 5908
rect 13320 5856 13326 5908
rect 14090 5856 14096 5908
rect 14148 5856 14154 5908
rect 14458 5856 14464 5908
rect 14516 5896 14522 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 14516 5868 14841 5896
rect 14516 5856 14522 5868
rect 14829 5865 14841 5868
rect 14875 5896 14887 5899
rect 15470 5896 15476 5908
rect 14875 5868 15476 5896
rect 14875 5865 14887 5868
rect 14829 5859 14887 5865
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16022 5896 16028 5908
rect 15887 5868 16028 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16022 5856 16028 5868
rect 16080 5856 16086 5908
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 17405 5899 17463 5905
rect 17405 5896 17417 5899
rect 17368 5868 17417 5896
rect 17368 5856 17374 5868
rect 17405 5865 17417 5868
rect 17451 5865 17463 5899
rect 17405 5859 17463 5865
rect 7147 5800 9076 5828
rect 7147 5797 7159 5800
rect 7101 5791 7159 5797
rect 9122 5788 9128 5840
rect 9180 5788 9186 5840
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 13449 5831 13507 5837
rect 9364 5800 9444 5828
rect 9364 5788 9370 5800
rect 4295 5732 4844 5760
rect 5092 5732 5212 5760
rect 5629 5763 5687 5769
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3252 5556 3280 5655
rect 3326 5652 3332 5704
rect 3384 5652 3390 5704
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5661 3479 5695
rect 3421 5655 3479 5661
rect 3436 5624 3464 5655
rect 3510 5652 3516 5704
rect 3568 5652 3574 5704
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3752 5664 4077 5692
rect 3752 5652 3758 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4338 5692 4344 5704
rect 4203 5664 4344 5692
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 5092 5701 5120 5732
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 5902 5760 5908 5772
rect 5675 5732 5908 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 7374 5760 7380 5772
rect 6748 5732 7380 5760
rect 6657 5705 6715 5711
rect 5077 5695 5135 5701
rect 5077 5692 5089 5695
rect 4856 5664 5089 5692
rect 4856 5652 4862 5664
rect 5077 5661 5089 5664
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5442 5692 5448 5704
rect 5215 5664 5448 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 4614 5624 4620 5636
rect 3436 5596 4620 5624
rect 4614 5584 4620 5596
rect 4672 5624 4678 5636
rect 5184 5624 5212 5655
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5810 5652 5816 5704
rect 5868 5652 5874 5704
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 6657 5671 6669 5705
rect 6703 5702 6715 5705
rect 6748 5702 6776 5732
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 7834 5720 7840 5772
rect 7892 5720 7898 5772
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8570 5760 8576 5772
rect 8168 5732 8576 5760
rect 8168 5720 8174 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 8757 5763 8815 5769
rect 8757 5729 8769 5763
rect 8803 5760 8815 5763
rect 9140 5760 9168 5788
rect 9416 5769 9444 5800
rect 13449 5797 13461 5831
rect 13495 5797 13507 5831
rect 13449 5791 13507 5797
rect 8803 5732 9168 5760
rect 9401 5763 9459 5769
rect 8803 5729 8815 5732
rect 8757 5723 8815 5729
rect 9401 5729 9413 5763
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 10318 5760 10324 5772
rect 9640 5732 10324 5760
rect 9640 5720 9646 5732
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10778 5720 10784 5772
rect 10836 5720 10842 5772
rect 12710 5720 12716 5772
rect 12768 5720 12774 5772
rect 13464 5760 13492 5791
rect 15286 5788 15292 5840
rect 15344 5828 15350 5840
rect 15381 5831 15439 5837
rect 15381 5828 15393 5831
rect 15344 5800 15393 5828
rect 15344 5788 15350 5800
rect 15381 5797 15393 5800
rect 15427 5797 15439 5831
rect 15381 5791 15439 5797
rect 12820 5732 13492 5760
rect 6703 5674 6776 5702
rect 6917 5695 6975 5701
rect 6703 5671 6715 5674
rect 6657 5665 6715 5671
rect 5997 5655 6055 5661
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 7852 5692 7880 5720
rect 6963 5664 7880 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 4672 5596 5212 5624
rect 4672 5584 4678 5596
rect 5350 5584 5356 5636
rect 5408 5584 5414 5636
rect 6012 5624 6040 5655
rect 8478 5652 8484 5704
rect 8536 5652 8542 5704
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8904 5664 9137 5692
rect 8904 5652 8910 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10796 5692 10824 5720
rect 10643 5664 10824 5692
rect 10873 5695 10931 5701
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 10873 5661 10885 5695
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 6086 5624 6092 5636
rect 6012 5596 6092 5624
rect 6086 5584 6092 5596
rect 6144 5624 6150 5636
rect 6144 5596 6868 5624
rect 6144 5584 6150 5596
rect 3694 5556 3700 5568
rect 3252 5528 3700 5556
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6604 5528 6745 5556
rect 6604 5516 6610 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6840 5556 6868 5596
rect 7834 5584 7840 5636
rect 7892 5624 7898 5636
rect 9324 5624 9352 5655
rect 7892 5596 9352 5624
rect 7892 5584 7898 5596
rect 9398 5584 9404 5636
rect 9456 5624 9462 5636
rect 10781 5627 10839 5633
rect 10781 5624 10793 5627
rect 9456 5596 10793 5624
rect 9456 5584 9462 5596
rect 10781 5593 10793 5596
rect 10827 5593 10839 5627
rect 10888 5624 10916 5655
rect 10962 5652 10968 5704
rect 11020 5652 11026 5704
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 12618 5692 12624 5704
rect 12575 5664 12624 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 11054 5624 11060 5636
rect 10888 5596 11060 5624
rect 10781 5587 10839 5593
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 12452 5624 12480 5655
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 12820 5701 12848 5732
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 14240 5732 14473 5760
rect 14240 5720 14246 5732
rect 14461 5729 14473 5732
rect 14507 5729 14519 5763
rect 14461 5723 14519 5729
rect 14550 5720 14556 5772
rect 14608 5720 14614 5772
rect 16298 5760 16304 5772
rect 15028 5732 16304 5760
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13170 5692 13176 5704
rect 13127 5664 13176 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13354 5652 13360 5704
rect 13412 5692 13418 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 13412 5664 13461 5692
rect 13412 5652 13418 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13449 5655 13507 5661
rect 13556 5664 13737 5692
rect 12897 5627 12955 5633
rect 12897 5624 12909 5627
rect 12452 5596 12909 5624
rect 12897 5593 12909 5596
rect 12943 5593 12955 5627
rect 12897 5587 12955 5593
rect 9950 5556 9956 5568
rect 6840 5528 9956 5556
rect 6733 5519 6791 5525
rect 9950 5516 9956 5528
rect 10008 5556 10014 5568
rect 10226 5556 10232 5568
rect 10008 5528 10232 5556
rect 10008 5516 10014 5528
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 10413 5559 10471 5565
rect 10413 5556 10425 5559
rect 10376 5528 10425 5556
rect 10376 5516 10382 5528
rect 10413 5525 10425 5528
rect 10459 5525 10471 5559
rect 10413 5519 10471 5525
rect 12066 5516 12072 5568
rect 12124 5556 12130 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 12124 5528 12265 5556
rect 12124 5516 12130 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12253 5519 12311 5525
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 13556 5556 13584 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 14274 5652 14280 5704
rect 14332 5652 14338 5704
rect 14366 5652 14372 5704
rect 14424 5652 14430 5704
rect 15028 5701 15056 5732
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 17221 5763 17279 5769
rect 17221 5760 17233 5763
rect 16500 5732 17233 5760
rect 15013 5695 15071 5701
rect 15013 5661 15025 5695
rect 15059 5661 15071 5695
rect 15013 5655 15071 5661
rect 15102 5652 15108 5704
rect 15160 5652 15166 5704
rect 15746 5652 15752 5704
rect 15804 5652 15810 5704
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 16500 5692 16528 5732
rect 17221 5729 17233 5732
rect 17267 5729 17279 5763
rect 17221 5723 17279 5729
rect 16172 5664 16528 5692
rect 16577 5695 16635 5701
rect 16172 5652 16178 5664
rect 16577 5661 16589 5695
rect 16623 5692 16635 5695
rect 16758 5692 16764 5704
rect 16623 5664 16764 5692
rect 16623 5661 16635 5664
rect 16577 5655 16635 5661
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 16942 5652 16948 5704
rect 17000 5692 17006 5704
rect 17037 5695 17095 5701
rect 17037 5692 17049 5695
rect 17000 5664 17049 5692
rect 17000 5652 17006 5664
rect 17037 5661 17049 5664
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 13630 5584 13636 5636
rect 13688 5584 13694 5636
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 15381 5627 15439 5633
rect 15381 5624 15393 5627
rect 13872 5596 15393 5624
rect 13872 5584 13878 5596
rect 15381 5593 15393 5596
rect 15427 5624 15439 5627
rect 15562 5624 15568 5636
rect 15427 5596 15568 5624
rect 15427 5593 15439 5596
rect 15381 5587 15439 5593
rect 15562 5584 15568 5596
rect 15620 5584 15626 5636
rect 15764 5624 15792 5652
rect 16132 5624 16160 5652
rect 15764 5596 16160 5624
rect 16206 5584 16212 5636
rect 16264 5584 16270 5636
rect 17052 5624 17080 5655
rect 17126 5652 17132 5704
rect 17184 5652 17190 5704
rect 17678 5624 17684 5636
rect 17052 5596 17684 5624
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 12492 5528 13584 5556
rect 12492 5516 12498 5528
rect 13722 5516 13728 5568
rect 13780 5556 13786 5568
rect 15102 5556 15108 5568
rect 13780 5528 15108 5556
rect 13780 5516 13786 5528
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 15194 5516 15200 5568
rect 15252 5516 15258 5568
rect 15930 5516 15936 5568
rect 15988 5556 15994 5568
rect 17126 5556 17132 5568
rect 15988 5528 17132 5556
rect 15988 5516 15994 5528
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 1104 5466 18492 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 18492 5466
rect 1104 5392 18492 5414
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 2924 5324 5028 5352
rect 2924 5312 2930 5324
rect 5000 5296 5028 5324
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 5868 5324 6377 5352
rect 5868 5312 5874 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 6696 5324 7788 5352
rect 6696 5312 6702 5324
rect 4982 5244 4988 5296
rect 5040 5284 5046 5296
rect 7760 5284 7788 5324
rect 7834 5312 7840 5364
rect 7892 5312 7898 5364
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9490 5352 9496 5364
rect 9263 5324 9496 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 9824 5324 10425 5352
rect 9824 5312 9830 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 11388 5324 12756 5352
rect 11388 5312 11394 5324
rect 8938 5284 8944 5296
rect 5040 5256 6592 5284
rect 7760 5256 8248 5284
rect 5040 5244 5046 5256
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3602 5216 3608 5228
rect 3375 5188 3608 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 3970 5216 3976 5228
rect 3835 5188 3976 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 3970 5176 3976 5188
rect 4028 5216 4034 5228
rect 4890 5216 4896 5228
rect 4028 5188 4896 5216
rect 4028 5176 4034 5188
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5592 5188 5641 5216
rect 5592 5176 5598 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 3694 5108 3700 5160
rect 3752 5108 3758 5160
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4249 5151 4307 5157
rect 4249 5148 4261 5151
rect 4120 5120 4261 5148
rect 4120 5108 4126 5120
rect 4249 5117 4261 5120
rect 4295 5117 4307 5151
rect 4249 5111 4307 5117
rect 4264 5080 4292 5111
rect 4338 5108 4344 5160
rect 4396 5108 4402 5160
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 4614 5148 4620 5160
rect 4571 5120 4620 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5353 5151 5411 5157
rect 5353 5117 5365 5151
rect 5399 5148 5411 5151
rect 5644 5148 5672 5179
rect 6086 5176 6092 5228
rect 6144 5176 6150 5228
rect 6564 5225 6592 5256
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 6871 5219 6929 5225
rect 6871 5185 6883 5219
rect 6917 5216 6929 5219
rect 7098 5216 7104 5228
rect 6917 5188 7104 5216
rect 6917 5185 6929 5188
rect 6871 5179 6929 5185
rect 6748 5148 6776 5179
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 7190 5176 7196 5228
rect 7248 5176 7254 5228
rect 7374 5225 7380 5228
rect 7341 5219 7380 5225
rect 7341 5185 7353 5219
rect 7341 5179 7380 5185
rect 7374 5176 7380 5179
rect 7432 5176 7438 5228
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 5399 5120 5580 5148
rect 5644 5120 6776 5148
rect 5399 5117 5411 5120
rect 5353 5111 5411 5117
rect 4801 5083 4859 5089
rect 4801 5080 4813 5083
rect 4264 5052 4813 5080
rect 4801 5049 4813 5052
rect 4847 5080 4859 5083
rect 5442 5080 5448 5092
rect 4847 5052 5448 5080
rect 4847 5049 4859 5052
rect 4801 5043 4859 5049
rect 5442 5040 5448 5052
rect 5500 5040 5506 5092
rect 5552 5080 5580 5120
rect 5994 5080 6000 5092
rect 5552 5052 6000 5080
rect 5994 5040 6000 5052
rect 6052 5040 6058 5092
rect 6748 5080 6776 5120
rect 7006 5108 7012 5160
rect 7064 5108 7070 5160
rect 7484 5148 7512 5179
rect 7558 5176 7564 5228
rect 7616 5176 7622 5228
rect 7650 5176 7656 5228
rect 7708 5225 7714 5228
rect 8220 5225 8248 5256
rect 8496 5256 8944 5284
rect 7708 5179 7716 5225
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 7708 5176 7714 5179
rect 8496 5148 8524 5256
rect 8938 5244 8944 5256
rect 8996 5244 9002 5296
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 10134 5284 10140 5296
rect 9180 5256 10140 5284
rect 9180 5244 9186 5256
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 11790 5284 11796 5296
rect 10612 5256 11796 5284
rect 8570 5176 8576 5228
rect 8628 5176 8634 5228
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8720 5188 8769 5216
rect 8720 5176 8726 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5185 9091 5219
rect 9033 5179 9091 5185
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10042 5216 10048 5228
rect 9999 5188 10048 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 7484 5120 8524 5148
rect 8846 5108 8852 5160
rect 8904 5148 8910 5160
rect 9048 5148 9076 5179
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 10612 5225 10640 5256
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 11900 5284 11928 5324
rect 11900 5256 12020 5284
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10870 5176 10876 5228
rect 10928 5176 10934 5228
rect 11992 5225 12020 5256
rect 12250 5244 12256 5296
rect 12308 5244 12314 5296
rect 12434 5244 12440 5296
rect 12492 5244 12498 5296
rect 12728 5284 12756 5324
rect 12802 5312 12808 5364
rect 12860 5312 12866 5364
rect 14093 5355 14151 5361
rect 14093 5321 14105 5355
rect 14139 5352 14151 5355
rect 14274 5352 14280 5364
rect 14139 5324 14280 5352
rect 14139 5321 14151 5324
rect 14093 5315 14151 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 14734 5312 14740 5364
rect 14792 5352 14798 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14792 5324 14933 5352
rect 14792 5312 14798 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 15562 5312 15568 5364
rect 15620 5312 15626 5364
rect 13725 5287 13783 5293
rect 12728 5256 13308 5284
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 12268 5216 12296 5244
rect 11977 5179 12035 5185
rect 12176 5188 12296 5216
rect 12345 5219 12403 5225
rect 11792 5151 11850 5157
rect 11792 5148 11804 5151
rect 8904 5120 11804 5148
rect 8904 5108 8910 5120
rect 11792 5117 11804 5120
rect 11838 5117 11850 5151
rect 11792 5111 11850 5117
rect 11882 5108 11888 5160
rect 11940 5108 11946 5160
rect 12069 5151 12127 5157
rect 12069 5117 12081 5151
rect 12115 5148 12127 5151
rect 12176 5148 12204 5188
rect 12345 5185 12357 5219
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 12115 5120 12204 5148
rect 12253 5151 12311 5157
rect 12115 5117 12127 5120
rect 12069 5111 12127 5117
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12360 5148 12388 5179
rect 12299 5120 12388 5148
rect 12544 5148 12572 5179
rect 12618 5176 12624 5228
rect 12676 5216 12682 5228
rect 12805 5219 12863 5225
rect 12676 5214 12756 5216
rect 12805 5214 12817 5219
rect 12676 5188 12817 5214
rect 12676 5176 12682 5188
rect 12728 5186 12817 5188
rect 12805 5185 12817 5186
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5216 13047 5219
rect 13170 5216 13176 5228
rect 13035 5188 13176 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 13280 5216 13308 5256
rect 13725 5253 13737 5287
rect 13771 5284 13783 5287
rect 15194 5284 15200 5296
rect 13771 5256 15200 5284
rect 13771 5253 13783 5256
rect 13725 5247 13783 5253
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 17034 5244 17040 5296
rect 17092 5284 17098 5296
rect 17129 5287 17187 5293
rect 17129 5284 17141 5287
rect 17092 5256 17141 5284
rect 17092 5244 17098 5256
rect 17129 5253 17141 5256
rect 17175 5253 17187 5287
rect 17129 5247 17187 5253
rect 13280 5214 13584 5216
rect 13630 5214 13636 5228
rect 13280 5188 13636 5214
rect 13556 5186 13636 5188
rect 13630 5176 13636 5186
rect 13688 5176 13694 5228
rect 13906 5176 13912 5228
rect 13964 5176 13970 5228
rect 14182 5176 14188 5228
rect 14240 5176 14246 5228
rect 14366 5176 14372 5228
rect 14424 5176 14430 5228
rect 14458 5176 14464 5228
rect 14516 5176 14522 5228
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 15010 5176 15016 5228
rect 15068 5216 15074 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 15068 5188 15117 5216
rect 15068 5176 15074 5188
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 15286 5176 15292 5228
rect 15344 5176 15350 5228
rect 15470 5176 15476 5228
rect 15528 5216 15534 5228
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 15528 5188 15761 5216
rect 15528 5176 15534 5188
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 16942 5176 16948 5228
rect 17000 5176 17006 5228
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 17276 5188 17325 5216
rect 17276 5176 17282 5188
rect 17313 5185 17325 5188
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 13998 5148 14004 5160
rect 12544 5120 14004 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 15378 5108 15384 5160
rect 15436 5108 15442 5160
rect 7466 5080 7472 5092
rect 6748 5052 7472 5080
rect 7466 5040 7472 5052
rect 7524 5040 7530 5092
rect 9398 5080 9404 5092
rect 7576 5052 9404 5080
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4764 4984 4997 5012
rect 4764 4972 4770 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 6012 5012 6040 5040
rect 7576 5024 7604 5052
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 9858 5040 9864 5092
rect 9916 5080 9922 5092
rect 10045 5083 10103 5089
rect 10045 5080 10057 5083
rect 9916 5052 10057 5080
rect 9916 5040 9922 5052
rect 10045 5049 10057 5052
rect 10091 5049 10103 5083
rect 10045 5043 10103 5049
rect 10137 5083 10195 5089
rect 10137 5049 10149 5083
rect 10183 5080 10195 5083
rect 10410 5080 10416 5092
rect 10183 5052 10416 5080
rect 10183 5049 10195 5052
rect 10137 5043 10195 5049
rect 10410 5040 10416 5052
rect 10468 5040 10474 5092
rect 10502 5040 10508 5092
rect 10560 5080 10566 5092
rect 10689 5083 10747 5089
rect 10689 5080 10701 5083
rect 10560 5052 10701 5080
rect 10560 5040 10566 5052
rect 10689 5049 10701 5052
rect 10735 5049 10747 5083
rect 10689 5043 10747 5049
rect 10781 5083 10839 5089
rect 10781 5049 10793 5083
rect 10827 5080 10839 5083
rect 13814 5080 13820 5092
rect 10827 5052 13820 5080
rect 10827 5049 10839 5052
rect 10781 5043 10839 5049
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 14829 5083 14887 5089
rect 14829 5049 14841 5083
rect 14875 5080 14887 5083
rect 15838 5080 15844 5092
rect 14875 5052 15844 5080
rect 14875 5049 14887 5052
rect 14829 5043 14887 5049
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 7558 5012 7564 5024
rect 6012 4984 7564 5012
rect 4985 4975 5043 4981
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7984 4984 8033 5012
rect 7984 4972 7990 4984
rect 8021 4981 8033 4984
rect 8067 4981 8079 5015
rect 8021 4975 8079 4981
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 9306 5012 9312 5024
rect 8628 4984 9312 5012
rect 8628 4972 8634 4984
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9732 4984 9781 5012
rect 9732 4972 9738 4984
rect 9769 4981 9781 4984
rect 9815 4981 9827 5015
rect 9769 4975 9827 4981
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 12250 5012 12256 5024
rect 11388 4984 12256 5012
rect 11388 4972 11394 4984
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 15286 4972 15292 5024
rect 15344 5012 15350 5024
rect 16850 5012 16856 5024
rect 15344 4984 16856 5012
rect 15344 4972 15350 4984
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 1104 4922 18492 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 18492 4922
rect 1104 4848 18492 4870
rect 2590 4768 2596 4820
rect 2648 4808 2654 4820
rect 3326 4808 3332 4820
rect 2648 4780 3332 4808
rect 2648 4768 2654 4780
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4614 4808 4620 4820
rect 4212 4780 4620 4808
rect 4212 4768 4218 4780
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5776 4780 5917 4808
rect 5776 4768 5782 4780
rect 5905 4777 5917 4780
rect 5951 4777 5963 4811
rect 5905 4771 5963 4777
rect 7098 4768 7104 4820
rect 7156 4768 7162 4820
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 7650 4808 7656 4820
rect 7423 4780 7656 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7800 4780 7849 4808
rect 7800 4768 7806 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 8757 4811 8815 4817
rect 8757 4777 8769 4811
rect 8803 4808 8815 4811
rect 8846 4808 8852 4820
rect 8803 4780 8852 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 8938 4768 8944 4820
rect 8996 4768 9002 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10045 4811 10103 4817
rect 10045 4808 10057 4811
rect 9824 4780 10057 4808
rect 9824 4768 9830 4780
rect 10045 4777 10057 4780
rect 10091 4777 10103 4811
rect 10045 4771 10103 4777
rect 10686 4768 10692 4820
rect 10744 4768 10750 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 11112 4780 11621 4808
rect 11112 4768 11118 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 11609 4771 11667 4777
rect 11790 4768 11796 4820
rect 11848 4768 11854 4820
rect 12526 4808 12532 4820
rect 12176 4780 12532 4808
rect 3878 4700 3884 4752
rect 3936 4740 3942 4752
rect 6270 4740 6276 4752
rect 3936 4712 6276 4740
rect 3936 4700 3942 4712
rect 6270 4700 6276 4712
rect 6328 4700 6334 4752
rect 7116 4740 7144 4768
rect 7469 4743 7527 4749
rect 7469 4740 7481 4743
rect 7116 4712 7481 4740
rect 7469 4709 7481 4712
rect 7515 4709 7527 4743
rect 7469 4703 7527 4709
rect 7929 4743 7987 4749
rect 7929 4709 7941 4743
rect 7975 4740 7987 4743
rect 11149 4743 11207 4749
rect 11149 4740 11161 4743
rect 7975 4712 11161 4740
rect 7975 4709 7987 4712
rect 7929 4703 7987 4709
rect 11149 4709 11161 4712
rect 11195 4740 11207 4743
rect 12176 4740 12204 4780
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 14185 4811 14243 4817
rect 14185 4777 14197 4811
rect 14231 4808 14243 4811
rect 14366 4808 14372 4820
rect 14231 4780 14372 4808
rect 14231 4777 14243 4780
rect 14185 4771 14243 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 14458 4768 14464 4820
rect 14516 4808 14522 4820
rect 14645 4811 14703 4817
rect 14645 4808 14657 4811
rect 14516 4780 14657 4808
rect 14516 4768 14522 4780
rect 14645 4777 14657 4780
rect 14691 4777 14703 4811
rect 14645 4771 14703 4777
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 15252 4780 15301 4808
rect 15252 4768 15258 4780
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15654 4808 15660 4820
rect 15289 4771 15347 4777
rect 15396 4780 15660 4808
rect 12342 4740 12348 4752
rect 11195 4712 12204 4740
rect 12268 4712 12348 4740
rect 11195 4709 11207 4712
rect 11149 4703 11207 4709
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6236 4644 6281 4672
rect 6236 4632 6242 4644
rect 6362 4632 6368 4684
rect 6420 4632 6426 4684
rect 7944 4672 7972 4703
rect 8662 4672 8668 4684
rect 7116 4644 7972 4672
rect 8220 4644 8668 4672
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3467 4576 4077 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 4065 4573 4077 4576
rect 4111 4604 4123 4607
rect 4154 4604 4160 4616
rect 4111 4576 4160 4604
rect 4111 4573 4123 4576
rect 4065 4567 4123 4573
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 4798 4604 4804 4616
rect 4264 4576 4804 4604
rect 3602 4496 3608 4548
rect 3660 4536 3666 4548
rect 4264 4536 4292 4576
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5350 4604 5356 4616
rect 4948 4576 5356 4604
rect 4948 4564 4954 4576
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5442 4564 5448 4616
rect 5500 4564 5506 4616
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 3660 4508 4292 4536
rect 4341 4539 4399 4545
rect 3660 4496 3666 4508
rect 4341 4505 4353 4539
rect 4387 4536 4399 4539
rect 4982 4536 4988 4548
rect 4387 4508 4988 4536
rect 4387 4505 4399 4508
rect 4341 4499 4399 4505
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 6104 4468 6132 4567
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 6454 4564 6460 4616
rect 6512 4604 6518 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6512 4576 6745 4604
rect 6512 4564 6518 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 6914 4564 6920 4616
rect 6972 4564 6978 4616
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7116 4613 7144 4644
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4604 7251 4607
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7239 4576 7757 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 7745 4573 7757 4576
rect 7791 4604 7803 4607
rect 7926 4604 7932 4616
rect 7791 4576 7932 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8018 4564 8024 4616
rect 8076 4564 8082 4616
rect 8220 4613 8248 4644
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 8772 4644 9904 4672
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 8772 4604 8800 4644
rect 8527 4576 8800 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 6178 4496 6184 4548
rect 6236 4536 6242 4548
rect 6638 4536 6644 4548
rect 6236 4508 6644 4536
rect 6236 4496 6242 4508
rect 6638 4496 6644 4508
rect 6696 4536 6702 4548
rect 8496 4536 8524 4567
rect 9122 4564 9128 4616
rect 9180 4564 9186 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9306 4604 9312 4616
rect 9263 4576 9312 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9306 4564 9312 4576
rect 9364 4604 9370 4616
rect 9876 4613 9904 4644
rect 10134 4632 10140 4684
rect 10192 4632 10198 4684
rect 11330 4632 11336 4684
rect 11388 4632 11394 4684
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 11480 4644 11652 4672
rect 11480 4632 11486 4644
rect 9861 4607 9919 4613
rect 9364 4576 9812 4604
rect 9364 4564 9370 4576
rect 6696 4508 8524 4536
rect 6696 4496 6702 4508
rect 8754 4496 8760 4548
rect 8812 4536 8818 4548
rect 9585 4539 9643 4545
rect 9585 4536 9597 4539
rect 8812 4508 9597 4536
rect 8812 4496 8818 4508
rect 9585 4505 9597 4508
rect 9631 4505 9643 4539
rect 9784 4536 9812 4576
rect 9861 4573 9873 4607
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 10686 4604 10692 4616
rect 10551 4576 10692 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4604 10839 4607
rect 11057 4607 11115 4613
rect 10827 4576 10916 4604
rect 10827 4573 10839 4576
rect 10781 4567 10839 4573
rect 10594 4536 10600 4548
rect 9784 4508 10600 4536
rect 9585 4499 9643 4505
rect 10594 4496 10600 4508
rect 10652 4496 10658 4548
rect 6730 4468 6736 4480
rect 6104 4440 6736 4468
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7742 4468 7748 4480
rect 7064 4440 7748 4468
rect 7064 4428 7070 4440
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 8570 4428 8576 4480
rect 8628 4468 8634 4480
rect 9122 4468 9128 4480
rect 8628 4440 9128 4468
rect 8628 4428 8634 4440
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 9766 4468 9772 4480
rect 9723 4440 9772 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 10226 4428 10232 4480
rect 10284 4428 10290 4480
rect 10888 4477 10916 4576
rect 11057 4573 11069 4607
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 10873 4471 10931 4477
rect 10873 4437 10885 4471
rect 10919 4437 10931 4471
rect 11072 4468 11100 4567
rect 11238 4564 11244 4616
rect 11296 4564 11302 4616
rect 11514 4564 11520 4616
rect 11572 4564 11578 4616
rect 11624 4604 11652 4644
rect 11882 4632 11888 4684
rect 11940 4632 11946 4684
rect 12158 4632 12164 4684
rect 12216 4632 12222 4684
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11624 4576 11989 4604
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 12066 4564 12072 4616
rect 12124 4564 12130 4616
rect 12268 4613 12296 4712
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 12434 4700 12440 4752
rect 12492 4740 12498 4752
rect 15396 4740 15424 4780
rect 15654 4768 15660 4780
rect 15712 4808 15718 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15712 4780 15853 4808
rect 15712 4768 15718 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 15841 4771 15899 4777
rect 12492 4712 15424 4740
rect 12492 4700 12498 4712
rect 15470 4700 15476 4752
rect 15528 4740 15534 4752
rect 17034 4740 17040 4752
rect 15528 4712 17040 4740
rect 15528 4700 15534 4712
rect 17034 4700 17040 4712
rect 17092 4700 17098 4752
rect 13906 4632 13912 4684
rect 13964 4672 13970 4684
rect 13964 4644 14320 4672
rect 13964 4632 13970 4644
rect 12253 4607 12311 4613
rect 12253 4604 12265 4607
rect 12176 4576 12265 4604
rect 12176 4468 12204 4576
rect 12253 4573 12265 4576
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 14292 4613 14320 4644
rect 14844 4644 16436 4672
rect 14844 4613 14872 4644
rect 16408 4616 16436 4644
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 16908 4644 17356 4672
rect 16908 4632 16914 4644
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13872 4576 14105 4604
rect 13872 4564 13878 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14829 4607 14887 4613
rect 14829 4604 14841 4607
rect 14323 4576 14841 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14829 4573 14841 4576
rect 14875 4573 14887 4607
rect 15197 4607 15255 4613
rect 15197 4604 15209 4607
rect 14829 4567 14887 4573
rect 14931 4576 15209 4604
rect 12986 4496 12992 4548
rect 13044 4536 13050 4548
rect 13446 4536 13452 4548
rect 13044 4508 13452 4536
rect 13044 4496 13050 4508
rect 13446 4496 13452 4508
rect 13504 4536 13510 4548
rect 14931 4536 14959 4576
rect 15197 4573 15209 4576
rect 15243 4604 15255 4607
rect 15286 4604 15292 4616
rect 15243 4576 15292 4604
rect 15243 4573 15255 4576
rect 15197 4567 15255 4573
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15470 4604 15476 4616
rect 15427 4576 15476 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 15562 4564 15568 4616
rect 15620 4564 15626 4616
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 16577 4607 16635 4613
rect 16577 4604 16589 4607
rect 16448 4576 16589 4604
rect 16448 4564 16454 4576
rect 16577 4573 16589 4576
rect 16623 4573 16635 4607
rect 16577 4567 16635 4573
rect 16942 4564 16948 4616
rect 17000 4564 17006 4616
rect 17328 4613 17356 4644
rect 17313 4607 17371 4613
rect 17313 4573 17325 4607
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 13504 4508 14959 4536
rect 15105 4539 15163 4545
rect 13504 4496 13510 4508
rect 15105 4505 15117 4539
rect 15151 4536 15163 4539
rect 15746 4536 15752 4548
rect 15151 4508 15752 4536
rect 15151 4505 15163 4508
rect 15105 4499 15163 4505
rect 15746 4496 15752 4508
rect 15804 4496 15810 4548
rect 11072 4440 12204 4468
rect 10873 4431 10931 4437
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 14458 4468 14464 4480
rect 12308 4440 14464 4468
rect 12308 4428 12314 4440
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14608 4440 15025 4468
rect 14608 4428 14614 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15013 4431 15071 4437
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 16853 4471 16911 4477
rect 16853 4468 16865 4471
rect 15252 4440 16865 4468
rect 15252 4428 15258 4440
rect 16853 4437 16865 4440
rect 16899 4437 16911 4471
rect 16853 4431 16911 4437
rect 1104 4378 18492 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 18492 4378
rect 1104 4304 18492 4326
rect 5350 4264 5356 4276
rect 4540 4236 5356 4264
rect 3602 4088 3608 4140
rect 3660 4088 3666 4140
rect 4540 4137 4568 4236
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 6178 4224 6184 4276
rect 6236 4224 6242 4276
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 10134 4264 10140 4276
rect 6328 4236 10140 4264
rect 6328 4224 6334 4236
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10226 4224 10232 4276
rect 10284 4224 10290 4276
rect 11238 4224 11244 4276
rect 11296 4264 11302 4276
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 11296 4236 11529 4264
rect 11296 4224 11302 4236
rect 11517 4233 11529 4236
rect 11563 4264 11575 4267
rect 11790 4264 11796 4276
rect 11563 4236 11796 4264
rect 11563 4233 11575 4236
rect 11517 4227 11575 4233
rect 11790 4224 11796 4236
rect 11848 4264 11854 4276
rect 12066 4264 12072 4276
rect 11848 4236 12072 4264
rect 11848 4224 11854 4236
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 12526 4224 12532 4276
rect 12584 4224 12590 4276
rect 13357 4267 13415 4273
rect 13357 4233 13369 4267
rect 13403 4264 13415 4267
rect 13814 4264 13820 4276
rect 13403 4236 13820 4264
rect 13403 4233 13415 4236
rect 13357 4227 13415 4233
rect 13814 4224 13820 4236
rect 13872 4224 13878 4276
rect 14550 4224 14556 4276
rect 14608 4264 14614 4276
rect 15930 4264 15936 4276
rect 14608 4236 15936 4264
rect 14608 4224 14614 4236
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 4614 4156 4620 4208
rect 4672 4196 4678 4208
rect 5997 4199 6055 4205
rect 5997 4196 6009 4199
rect 4672 4168 6009 4196
rect 4672 4156 4678 4168
rect 5997 4165 6009 4168
rect 6043 4165 6055 4199
rect 5997 4159 6055 4165
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 8297 4199 8355 4205
rect 8297 4196 8309 4199
rect 6972 4168 8309 4196
rect 6972 4156 6978 4168
rect 8297 4165 8309 4168
rect 8343 4196 8355 4199
rect 8386 4196 8392 4208
rect 8343 4168 8392 4196
rect 8343 4165 8355 4168
rect 8297 4159 8355 4165
rect 8386 4156 8392 4168
rect 8444 4196 8450 4208
rect 8754 4196 8760 4208
rect 8444 4168 8760 4196
rect 8444 4156 8450 4168
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 8864 4168 9352 4196
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 5350 4088 5356 4140
rect 5408 4128 5414 4140
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5408 4100 5825 4128
rect 5408 4088 5414 4100
rect 5813 4097 5825 4100
rect 5859 4128 5871 4131
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 5859 4100 6469 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6822 4088 6828 4140
rect 6880 4088 6886 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 8864 4128 8892 4168
rect 7524 4100 8892 4128
rect 8941 4131 8999 4137
rect 7524 4088 7530 4100
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 9214 4128 9220 4140
rect 8987 4100 9220 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9324 4128 9352 4168
rect 10686 4156 10692 4208
rect 10744 4196 10750 4208
rect 15194 4196 15200 4208
rect 10744 4168 15200 4196
rect 10744 4156 10750 4168
rect 15194 4156 15200 4168
rect 15252 4156 15258 4208
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9324 4100 9413 4128
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 9401 4091 9459 4097
rect 9600 4100 10149 4128
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 6270 4060 6276 4072
rect 5491 4032 6276 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 9490 4060 9496 4072
rect 8352 4032 9496 4060
rect 8352 4020 8358 4032
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 8570 3992 8576 4004
rect 8527 3964 8576 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 8680 4001 8708 4032
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 9600 4001 9628 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10502 4088 10508 4140
rect 10560 4088 10566 4140
rect 12986 4128 12992 4140
rect 11716 4100 12992 4128
rect 9674 4020 9680 4072
rect 9732 4020 9738 4072
rect 10318 4020 10324 4072
rect 10376 4020 10382 4072
rect 11716 4001 11744 4100
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13136 4100 13829 4128
rect 13136 4088 13142 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 11977 4063 12035 4069
rect 11977 4029 11989 4063
rect 12023 4060 12035 4063
rect 13832 4060 13860 4091
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 13964 4100 14381 4128
rect 13964 4088 13970 4100
rect 14369 4097 14381 4100
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14516 4100 14565 4128
rect 14516 4088 14522 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16448 4100 16681 4128
rect 16448 4088 16454 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16762 4131 16820 4137
rect 16762 4097 16774 4131
rect 16808 4128 16820 4131
rect 16942 4128 16948 4140
rect 16808 4100 16948 4128
rect 16808 4097 16820 4100
rect 16762 4091 16820 4097
rect 14274 4060 14280 4072
rect 12023 4032 13492 4060
rect 13832 4032 14280 4060
rect 12023 4029 12035 4032
rect 11977 4023 12035 4029
rect 8665 3995 8723 4001
rect 8665 3961 8677 3995
rect 8711 3961 8723 3995
rect 8665 3955 8723 3961
rect 9585 3995 9643 4001
rect 9585 3961 9597 3995
rect 9631 3961 9643 3995
rect 9585 3955 9643 3961
rect 11701 3995 11759 4001
rect 11701 3961 11713 3995
rect 11747 3961 11759 3995
rect 11701 3955 11759 3961
rect 12713 3995 12771 4001
rect 12713 3961 12725 3995
rect 12759 3992 12771 3995
rect 12894 3992 12900 4004
rect 12759 3964 12900 3992
rect 12759 3961 12771 3964
rect 12713 3955 12771 3961
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 13464 4001 13492 4032
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 15562 4060 15568 4072
rect 14476 4032 15568 4060
rect 13449 3995 13507 4001
rect 13449 3961 13461 3995
rect 13495 3992 13507 3995
rect 14476 3992 14504 4032
rect 15562 4020 15568 4032
rect 15620 4060 15626 4072
rect 16776 4060 16804 4091
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 15620 4032 16804 4060
rect 15620 4020 15626 4032
rect 13495 3964 14504 3992
rect 14553 3995 14611 4001
rect 13495 3961 13507 3964
rect 13449 3955 13507 3961
rect 14553 3961 14565 3995
rect 14599 3992 14611 3995
rect 15378 3992 15384 4004
rect 14599 3964 15384 3992
rect 14599 3961 14611 3964
rect 14553 3955 14611 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 9493 3927 9551 3933
rect 9493 3893 9505 3927
rect 9539 3924 9551 3927
rect 9766 3924 9772 3936
rect 9539 3896 9772 3924
rect 9539 3893 9551 3896
rect 9493 3887 9551 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10502 3884 10508 3936
rect 10560 3884 10566 3936
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 16853 3927 16911 3933
rect 16853 3924 16865 3927
rect 16816 3896 16865 3924
rect 16816 3884 16822 3896
rect 16853 3893 16865 3896
rect 16899 3893 16911 3927
rect 16853 3887 16911 3893
rect 1104 3834 18492 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 18492 3834
rect 1104 3760 18492 3782
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7285 3723 7343 3729
rect 7285 3720 7297 3723
rect 7064 3692 7297 3720
rect 7064 3680 7070 3692
rect 7285 3689 7297 3692
rect 7331 3689 7343 3723
rect 7285 3683 7343 3689
rect 6822 3612 6828 3664
rect 6880 3652 6886 3664
rect 7377 3655 7435 3661
rect 7377 3652 7389 3655
rect 6880 3624 7389 3652
rect 6880 3612 6886 3624
rect 7377 3621 7389 3624
rect 7423 3621 7435 3655
rect 7377 3615 7435 3621
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3584 7803 3587
rect 8018 3584 8024 3596
rect 7791 3556 8024 3584
rect 7791 3553 7803 3556
rect 7745 3547 7803 3553
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 1104 3290 18492 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 18492 3290
rect 1104 3216 18492 3238
rect 1104 2746 18492 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 18492 2746
rect 1104 2672 18492 2694
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 1104 2202 18492 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 18492 2202
rect 1104 2128 18492 2150
<< via1 >>
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 7748 18912 7800 18964
rect 9680 18912 9732 18964
rect 11612 18912 11664 18964
rect 8944 18844 8996 18896
rect 12624 18844 12676 18896
rect 7932 18776 7984 18828
rect 10324 18776 10376 18828
rect 8024 18708 8076 18760
rect 9404 18708 9456 18760
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 13912 18708 13964 18760
rect 16580 18708 16632 18760
rect 7288 18640 7340 18692
rect 9588 18683 9640 18692
rect 9588 18649 9597 18683
rect 9597 18649 9631 18683
rect 9631 18649 9640 18683
rect 9588 18640 9640 18649
rect 16672 18640 16724 18692
rect 11888 18572 11940 18624
rect 15384 18572 15436 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 1952 18368 2004 18420
rect 2320 18275 2372 18284
rect 2320 18241 2329 18275
rect 2329 18241 2363 18275
rect 2363 18241 2372 18275
rect 2320 18232 2372 18241
rect 2228 18071 2280 18080
rect 2228 18037 2237 18071
rect 2237 18037 2271 18071
rect 2271 18037 2280 18071
rect 2228 18028 2280 18037
rect 3608 18071 3660 18080
rect 3608 18037 3617 18071
rect 3617 18037 3651 18071
rect 3651 18037 3660 18071
rect 3608 18028 3660 18037
rect 7104 18275 7156 18284
rect 7104 18241 7113 18275
rect 7113 18241 7147 18275
rect 7147 18241 7156 18275
rect 7104 18232 7156 18241
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 8024 18411 8076 18420
rect 8024 18377 8033 18411
rect 8033 18377 8067 18411
rect 8067 18377 8076 18411
rect 8024 18368 8076 18377
rect 9404 18411 9456 18420
rect 9404 18377 9413 18411
rect 9413 18377 9447 18411
rect 9447 18377 9456 18411
rect 9404 18368 9456 18377
rect 10324 18368 10376 18420
rect 8024 18232 8076 18284
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 8300 18207 8352 18216
rect 8300 18173 8309 18207
rect 8309 18173 8343 18207
rect 8343 18173 8352 18207
rect 8300 18164 8352 18173
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 8576 18207 8628 18216
rect 8576 18173 8585 18207
rect 8585 18173 8619 18207
rect 8619 18173 8628 18207
rect 8576 18164 8628 18173
rect 10140 18232 10192 18284
rect 11888 18343 11940 18352
rect 11888 18309 11897 18343
rect 11897 18309 11931 18343
rect 11931 18309 11940 18343
rect 13360 18368 13412 18420
rect 11888 18300 11940 18309
rect 13728 18300 13780 18352
rect 12992 18275 13044 18284
rect 9772 18139 9824 18148
rect 9772 18105 9781 18139
rect 9781 18105 9815 18139
rect 9815 18105 9824 18139
rect 9772 18096 9824 18105
rect 10232 18207 10284 18216
rect 10232 18173 10241 18207
rect 10241 18173 10275 18207
rect 10275 18173 10284 18207
rect 10232 18164 10284 18173
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 11980 18164 12032 18216
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 15476 18232 15528 18284
rect 16028 18232 16080 18284
rect 16396 18275 16448 18284
rect 16396 18241 16405 18275
rect 16405 18241 16439 18275
rect 16439 18241 16448 18275
rect 16396 18232 16448 18241
rect 16580 18232 16632 18284
rect 15016 18207 15068 18216
rect 15016 18173 15025 18207
rect 15025 18173 15059 18207
rect 15059 18173 15068 18207
rect 15016 18164 15068 18173
rect 15108 18164 15160 18216
rect 11980 18071 12032 18080
rect 11980 18037 11989 18071
rect 11989 18037 12023 18071
rect 12023 18037 12032 18071
rect 11980 18028 12032 18037
rect 16212 18096 16264 18148
rect 14372 18028 14424 18080
rect 16764 18071 16816 18080
rect 16764 18037 16773 18071
rect 16773 18037 16807 18071
rect 16807 18037 16816 18071
rect 16764 18028 16816 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 7840 17824 7892 17876
rect 2412 17756 2464 17808
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 2596 17552 2648 17604
rect 3608 17688 3660 17740
rect 6736 17756 6788 17808
rect 9036 17824 9088 17876
rect 9772 17824 9824 17876
rect 10232 17824 10284 17876
rect 11704 17824 11756 17876
rect 8300 17756 8352 17808
rect 3884 17663 3936 17672
rect 3884 17629 3893 17663
rect 3893 17629 3927 17663
rect 3927 17629 3936 17663
rect 3884 17620 3936 17629
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 8116 17620 8168 17672
rect 10784 17688 10836 17740
rect 12992 17867 13044 17876
rect 12992 17833 13001 17867
rect 13001 17833 13035 17867
rect 13035 17833 13044 17867
rect 12992 17824 13044 17833
rect 13176 17824 13228 17876
rect 13728 17824 13780 17876
rect 13268 17756 13320 17808
rect 8484 17620 8536 17672
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 9220 17663 9272 17672
rect 9220 17629 9229 17663
rect 9229 17629 9263 17663
rect 9263 17629 9272 17663
rect 9220 17620 9272 17629
rect 9956 17620 10008 17672
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 10416 17663 10468 17672
rect 10416 17629 10425 17663
rect 10425 17629 10459 17663
rect 10459 17629 10468 17663
rect 10416 17620 10468 17629
rect 10600 17620 10652 17672
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 14464 17824 14516 17876
rect 15108 17824 15160 17876
rect 3792 17552 3844 17604
rect 7196 17552 7248 17604
rect 7748 17552 7800 17604
rect 8024 17595 8076 17604
rect 8024 17561 8033 17595
rect 8033 17561 8067 17595
rect 8067 17561 8076 17595
rect 8024 17552 8076 17561
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3240 17484 3292 17493
rect 3700 17484 3752 17536
rect 4068 17527 4120 17536
rect 4068 17493 4077 17527
rect 4077 17493 4111 17527
rect 4111 17493 4120 17527
rect 4068 17484 4120 17493
rect 4804 17484 4856 17536
rect 7656 17484 7708 17536
rect 8760 17552 8812 17604
rect 8852 17484 8904 17536
rect 9312 17527 9364 17536
rect 9312 17493 9321 17527
rect 9321 17493 9355 17527
rect 9355 17493 9364 17527
rect 9312 17484 9364 17493
rect 11704 17595 11756 17604
rect 11704 17561 11713 17595
rect 11713 17561 11747 17595
rect 11747 17561 11756 17595
rect 11704 17552 11756 17561
rect 10508 17484 10560 17536
rect 10600 17484 10652 17536
rect 10968 17484 11020 17536
rect 11336 17484 11388 17536
rect 11980 17552 12032 17604
rect 12716 17620 12768 17672
rect 14372 17731 14424 17740
rect 14372 17697 14381 17731
rect 14381 17697 14415 17731
rect 14415 17697 14424 17731
rect 14372 17688 14424 17697
rect 15016 17688 15068 17740
rect 16212 17731 16264 17740
rect 16212 17697 16221 17731
rect 16221 17697 16255 17731
rect 16255 17697 16264 17731
rect 16212 17688 16264 17697
rect 12624 17595 12676 17604
rect 12624 17561 12633 17595
rect 12633 17561 12667 17595
rect 12667 17561 12676 17595
rect 12624 17552 12676 17561
rect 13912 17663 13964 17672
rect 13912 17629 13921 17663
rect 13921 17629 13955 17663
rect 13955 17629 13964 17663
rect 13912 17620 13964 17629
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 12256 17484 12308 17536
rect 14648 17552 14700 17604
rect 15384 17552 15436 17604
rect 16764 17552 16816 17604
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 15936 17484 15988 17536
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 5816 17280 5868 17332
rect 3240 17212 3292 17264
rect 1952 17144 2004 17196
rect 3332 17187 3384 17196
rect 3332 17153 3341 17187
rect 3341 17153 3375 17187
rect 3375 17153 3384 17187
rect 3332 17144 3384 17153
rect 2688 17076 2740 17128
rect 3792 17144 3844 17196
rect 4620 17187 4672 17196
rect 4620 17153 4629 17187
rect 4629 17153 4663 17187
rect 4663 17153 4672 17187
rect 4620 17144 4672 17153
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 5724 17187 5776 17196
rect 5724 17153 5733 17187
rect 5733 17153 5767 17187
rect 5767 17153 5776 17187
rect 5724 17144 5776 17153
rect 6276 17144 6328 17196
rect 7104 17187 7156 17196
rect 7104 17153 7113 17187
rect 7113 17153 7147 17187
rect 7147 17153 7156 17187
rect 7104 17144 7156 17153
rect 7656 17323 7708 17332
rect 7656 17289 7665 17323
rect 7665 17289 7699 17323
rect 7699 17289 7708 17323
rect 7656 17280 7708 17289
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 9220 17280 9272 17332
rect 9312 17280 9364 17332
rect 9772 17280 9824 17332
rect 7380 17144 7432 17196
rect 2412 17051 2464 17060
rect 2412 17017 2421 17051
rect 2421 17017 2455 17051
rect 2455 17017 2464 17051
rect 2412 17008 2464 17017
rect 6736 17076 6788 17128
rect 7472 17119 7524 17128
rect 7472 17085 7481 17119
rect 7481 17085 7515 17119
rect 7515 17085 7524 17119
rect 7472 17076 7524 17085
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 7196 17008 7248 17060
rect 8576 17076 8628 17128
rect 8852 17187 8904 17196
rect 8852 17153 8861 17187
rect 8861 17153 8895 17187
rect 8895 17153 8904 17187
rect 8852 17144 8904 17153
rect 8944 17187 8996 17196
rect 8944 17153 8953 17187
rect 8953 17153 8987 17187
rect 8987 17153 8996 17187
rect 8944 17144 8996 17153
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9036 17144 9088 17153
rect 9220 17187 9272 17196
rect 9220 17153 9227 17187
rect 9227 17153 9272 17187
rect 9220 17144 9272 17153
rect 9312 17187 9364 17196
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 9772 17144 9824 17196
rect 9680 17076 9732 17128
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 12256 17323 12308 17332
rect 12256 17289 12265 17323
rect 12265 17289 12299 17323
rect 12299 17289 12308 17323
rect 12256 17280 12308 17289
rect 14096 17280 14148 17332
rect 13268 17212 13320 17264
rect 15016 17280 15068 17332
rect 16396 17280 16448 17332
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 9128 17008 9180 17060
rect 1860 16940 1912 16992
rect 2044 16983 2096 16992
rect 2044 16949 2053 16983
rect 2053 16949 2087 16983
rect 2087 16949 2096 16983
rect 2044 16940 2096 16949
rect 3056 16983 3108 16992
rect 3056 16949 3065 16983
rect 3065 16949 3099 16983
rect 3099 16949 3108 16983
rect 3056 16940 3108 16949
rect 5080 16940 5132 16992
rect 5448 16940 5500 16992
rect 6184 16940 6236 16992
rect 7012 16940 7064 16992
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 7288 16940 7340 16949
rect 7564 16940 7616 16992
rect 8392 16940 8444 16992
rect 9588 16940 9640 16992
rect 9680 16940 9732 16992
rect 9864 16940 9916 16992
rect 10324 17076 10376 17128
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 12072 17187 12124 17196
rect 12072 17153 12081 17187
rect 12081 17153 12115 17187
rect 12115 17153 12124 17187
rect 12072 17144 12124 17153
rect 14188 17144 14240 17196
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 16488 17187 16540 17196
rect 16488 17153 16497 17187
rect 16497 17153 16531 17187
rect 16531 17153 16540 17187
rect 16488 17144 16540 17153
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 16672 17144 16724 17153
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 12808 17076 12860 17128
rect 16304 17076 16356 17128
rect 11612 17008 11664 17060
rect 11980 17008 12032 17060
rect 10232 16940 10284 16992
rect 10692 16940 10744 16992
rect 13544 16940 13596 16992
rect 14924 16940 14976 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 1676 16736 1728 16788
rect 3424 16779 3476 16788
rect 3424 16745 3433 16779
rect 3433 16745 3467 16779
rect 3467 16745 3476 16779
rect 3424 16736 3476 16745
rect 3516 16736 3568 16788
rect 3884 16736 3936 16788
rect 5724 16736 5776 16788
rect 3148 16668 3200 16720
rect 3332 16668 3384 16720
rect 3608 16668 3660 16720
rect 2504 16600 2556 16652
rect 1860 16575 1912 16584
rect 1860 16541 1869 16575
rect 1869 16541 1903 16575
rect 1903 16541 1912 16575
rect 1860 16532 1912 16541
rect 2320 16532 2372 16584
rect 2688 16575 2740 16584
rect 2688 16541 2697 16575
rect 2697 16541 2731 16575
rect 2731 16541 2740 16575
rect 2688 16532 2740 16541
rect 4804 16668 4856 16720
rect 7104 16736 7156 16788
rect 7380 16779 7432 16788
rect 7380 16745 7389 16779
rect 7389 16745 7423 16779
rect 7423 16745 7432 16779
rect 7380 16736 7432 16745
rect 9128 16736 9180 16788
rect 9312 16736 9364 16788
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 10508 16736 10560 16788
rect 12072 16736 12124 16788
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 16764 16736 16816 16788
rect 3240 16532 3292 16584
rect 3516 16575 3568 16584
rect 3516 16541 3524 16575
rect 3524 16541 3558 16575
rect 3558 16541 3568 16575
rect 3516 16532 3568 16541
rect 3608 16575 3660 16584
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 3700 16532 3752 16584
rect 2136 16396 2188 16448
rect 3884 16464 3936 16516
rect 7012 16711 7064 16720
rect 7012 16677 7021 16711
rect 7021 16677 7055 16711
rect 7055 16677 7064 16711
rect 7012 16668 7064 16677
rect 8944 16668 8996 16720
rect 12348 16668 12400 16720
rect 4160 16507 4212 16516
rect 4160 16473 4169 16507
rect 4169 16473 4203 16507
rect 4203 16473 4212 16507
rect 4160 16464 4212 16473
rect 4896 16507 4948 16516
rect 4896 16473 4905 16507
rect 4905 16473 4939 16507
rect 4939 16473 4948 16507
rect 4896 16464 4948 16473
rect 5080 16575 5132 16584
rect 5080 16541 5125 16575
rect 5125 16541 5132 16575
rect 5080 16532 5132 16541
rect 5632 16532 5684 16584
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 6368 16532 6420 16584
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 6460 16507 6512 16516
rect 6460 16473 6469 16507
rect 6469 16473 6503 16507
rect 6503 16473 6512 16507
rect 6460 16464 6512 16473
rect 7012 16532 7064 16584
rect 7564 16532 7616 16584
rect 8576 16600 8628 16652
rect 7840 16507 7892 16516
rect 7840 16473 7849 16507
rect 7849 16473 7883 16507
rect 7883 16473 7892 16507
rect 7840 16464 7892 16473
rect 8852 16464 8904 16516
rect 9220 16532 9272 16584
rect 9496 16575 9548 16584
rect 9496 16541 9505 16575
rect 9505 16541 9539 16575
rect 9539 16541 9548 16575
rect 9496 16532 9548 16541
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 11244 16600 11296 16652
rect 9772 16507 9824 16516
rect 9772 16473 9781 16507
rect 9781 16473 9815 16507
rect 9815 16473 9824 16507
rect 9772 16464 9824 16473
rect 10232 16532 10284 16584
rect 10692 16532 10744 16584
rect 11796 16643 11848 16652
rect 11796 16609 11805 16643
rect 11805 16609 11839 16643
rect 11839 16609 11848 16643
rect 11796 16600 11848 16609
rect 11980 16600 12032 16652
rect 12440 16600 12492 16652
rect 12256 16532 12308 16584
rect 13176 16575 13228 16584
rect 13176 16541 13185 16575
rect 13185 16541 13219 16575
rect 13219 16541 13228 16575
rect 13176 16532 13228 16541
rect 13268 16575 13320 16584
rect 13268 16541 13277 16575
rect 13277 16541 13311 16575
rect 13311 16541 13320 16575
rect 13268 16532 13320 16541
rect 13912 16600 13964 16652
rect 14464 16600 14516 16652
rect 15844 16600 15896 16652
rect 16764 16600 16816 16652
rect 14924 16532 14976 16584
rect 15384 16575 15436 16584
rect 15384 16541 15393 16575
rect 15393 16541 15427 16575
rect 15427 16541 15436 16575
rect 15384 16532 15436 16541
rect 14188 16464 14240 16516
rect 7196 16396 7248 16448
rect 9864 16439 9916 16448
rect 9864 16405 9879 16439
rect 9879 16405 9913 16439
rect 9913 16405 9916 16439
rect 9864 16396 9916 16405
rect 10048 16396 10100 16448
rect 10324 16396 10376 16448
rect 10508 16396 10560 16448
rect 11704 16396 11756 16448
rect 14004 16396 14056 16448
rect 14556 16396 14608 16448
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 1860 16192 1912 16244
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 1768 16056 1820 16108
rect 2320 16056 2372 16108
rect 4160 16192 4212 16244
rect 2872 16124 2924 16176
rect 3424 16124 3476 16176
rect 3056 16056 3108 16108
rect 2136 16031 2188 16040
rect 2136 15997 2145 16031
rect 2145 15997 2179 16031
rect 2179 15997 2188 16031
rect 2136 15988 2188 15997
rect 1860 15920 1912 15972
rect 2044 15920 2096 15972
rect 4068 15988 4120 16040
rect 3700 15920 3752 15972
rect 4804 16056 4856 16108
rect 5080 16056 5132 16108
rect 5356 16124 5408 16176
rect 5264 16056 5316 16108
rect 5540 16056 5592 16108
rect 5816 16056 5868 16108
rect 6184 16056 6236 16108
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 6920 16056 6972 16065
rect 6276 15988 6328 16040
rect 8760 16124 8812 16176
rect 9312 16124 9364 16176
rect 1676 15852 1728 15904
rect 3148 15852 3200 15904
rect 5724 15963 5776 15972
rect 5724 15929 5733 15963
rect 5733 15929 5767 15963
rect 5767 15929 5776 15963
rect 5724 15920 5776 15929
rect 6000 15920 6052 15972
rect 6828 15963 6880 15972
rect 6828 15929 6837 15963
rect 6837 15929 6871 15963
rect 6871 15929 6880 15963
rect 6828 15920 6880 15929
rect 7012 15920 7064 15972
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 10324 16124 10376 16176
rect 9956 16056 10008 16108
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 11336 16235 11388 16244
rect 11336 16201 11345 16235
rect 11345 16201 11379 16235
rect 11379 16201 11388 16235
rect 11336 16192 11388 16201
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 10876 16167 10928 16176
rect 10876 16133 10885 16167
rect 10885 16133 10919 16167
rect 10919 16133 10928 16167
rect 10876 16124 10928 16133
rect 11428 16124 11480 16176
rect 11152 16099 11204 16108
rect 10048 15988 10100 16040
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 11336 16056 11388 16108
rect 12072 16124 12124 16176
rect 13268 16192 13320 16244
rect 13912 16192 13964 16244
rect 14556 16192 14608 16244
rect 12348 16124 12400 16176
rect 14004 16124 14056 16176
rect 10784 15988 10836 16040
rect 10968 15988 11020 16040
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 12072 15988 12124 16040
rect 13452 16099 13504 16108
rect 13452 16065 13461 16099
rect 13461 16065 13495 16099
rect 13495 16065 13504 16099
rect 13452 16056 13504 16065
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 13912 16056 13964 16108
rect 14464 16167 14516 16176
rect 14464 16133 14473 16167
rect 14473 16133 14507 16167
rect 14507 16133 14516 16167
rect 14464 16124 14516 16133
rect 15384 16124 15436 16176
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 16764 16124 16816 16176
rect 15476 15988 15528 16040
rect 16948 15988 17000 16040
rect 10416 15920 10468 15972
rect 5264 15852 5316 15904
rect 6092 15852 6144 15904
rect 6460 15852 6512 15904
rect 8024 15852 8076 15904
rect 9772 15852 9824 15904
rect 9864 15895 9916 15904
rect 9864 15861 9873 15895
rect 9873 15861 9907 15895
rect 9907 15861 9916 15895
rect 9864 15852 9916 15861
rect 10692 15852 10744 15904
rect 13544 15920 13596 15972
rect 12164 15852 12216 15904
rect 14004 15895 14056 15904
rect 14004 15861 14013 15895
rect 14013 15861 14047 15895
rect 14047 15861 14056 15895
rect 14004 15852 14056 15861
rect 15292 15920 15344 15972
rect 15936 15920 15988 15972
rect 15200 15852 15252 15904
rect 15568 15852 15620 15904
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 1308 15648 1360 15700
rect 3884 15648 3936 15700
rect 2964 15580 3016 15632
rect 4712 15648 4764 15700
rect 5172 15648 5224 15700
rect 5632 15648 5684 15700
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 2780 15487 2832 15496
rect 2780 15453 2789 15487
rect 2789 15453 2823 15487
rect 2823 15453 2832 15487
rect 2780 15444 2832 15453
rect 3240 15512 3292 15564
rect 3884 15512 3936 15564
rect 6092 15580 6144 15632
rect 6552 15623 6604 15632
rect 6552 15589 6561 15623
rect 6561 15589 6595 15623
rect 6595 15589 6604 15623
rect 6552 15580 6604 15589
rect 6828 15648 6880 15700
rect 7380 15648 7432 15700
rect 7932 15648 7984 15700
rect 8392 15648 8444 15700
rect 8760 15648 8812 15700
rect 9496 15648 9548 15700
rect 10048 15648 10100 15700
rect 10876 15648 10928 15700
rect 12164 15691 12216 15700
rect 12164 15657 12173 15691
rect 12173 15657 12207 15691
rect 12207 15657 12216 15691
rect 12164 15648 12216 15657
rect 12256 15648 12308 15700
rect 7840 15580 7892 15632
rect 5080 15555 5132 15564
rect 5080 15521 5089 15555
rect 5089 15521 5123 15555
rect 5123 15521 5132 15555
rect 5080 15512 5132 15521
rect 6184 15555 6236 15564
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 3332 15487 3384 15496
rect 3332 15453 3341 15487
rect 3341 15453 3375 15487
rect 3375 15453 3384 15487
rect 3332 15444 3384 15453
rect 3424 15487 3476 15496
rect 3424 15453 3433 15487
rect 3433 15453 3467 15487
rect 3467 15453 3476 15487
rect 3424 15444 3476 15453
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 3608 15376 3660 15428
rect 4712 15376 4764 15428
rect 5356 15444 5408 15496
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 6276 15555 6328 15564
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 6276 15512 6328 15521
rect 6920 15512 6972 15564
rect 5632 15487 5684 15496
rect 5632 15453 5641 15487
rect 5641 15453 5675 15487
rect 5675 15453 5684 15487
rect 5632 15444 5684 15453
rect 6736 15444 6788 15496
rect 7472 15487 7524 15496
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 7656 15444 7708 15496
rect 9128 15512 9180 15564
rect 9496 15555 9548 15564
rect 9496 15521 9505 15555
rect 9505 15521 9539 15555
rect 9539 15521 9548 15555
rect 9496 15512 9548 15521
rect 9680 15580 9732 15632
rect 9864 15580 9916 15632
rect 13084 15648 13136 15700
rect 15936 15648 15988 15700
rect 11428 15512 11480 15564
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 8392 15444 8444 15496
rect 8944 15444 8996 15496
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 9680 15444 9732 15496
rect 6368 15376 6420 15428
rect 1952 15308 2004 15360
rect 2136 15308 2188 15360
rect 5172 15308 5224 15360
rect 6000 15308 6052 15360
rect 6920 15308 6972 15360
rect 7104 15376 7156 15428
rect 10324 15444 10376 15496
rect 10876 15444 10928 15496
rect 11060 15444 11112 15496
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 11520 15444 11572 15453
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 8116 15308 8168 15360
rect 9036 15308 9088 15360
rect 9588 15308 9640 15360
rect 9956 15308 10008 15360
rect 10232 15351 10284 15360
rect 10232 15317 10257 15351
rect 10257 15317 10284 15351
rect 10416 15376 10468 15428
rect 11244 15376 11296 15428
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 12164 15444 12216 15496
rect 13360 15444 13412 15496
rect 15108 15512 15160 15564
rect 15660 15512 15712 15564
rect 16856 15512 16908 15564
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 15844 15444 15896 15496
rect 12532 15376 12584 15428
rect 15384 15376 15436 15428
rect 16212 15419 16264 15428
rect 16212 15385 16221 15419
rect 16221 15385 16255 15419
rect 16255 15385 16264 15419
rect 16212 15376 16264 15385
rect 17868 15376 17920 15428
rect 10232 15308 10284 15317
rect 12256 15308 12308 15360
rect 12900 15308 12952 15360
rect 13452 15308 13504 15360
rect 14740 15308 14792 15360
rect 17684 15351 17736 15360
rect 17684 15317 17693 15351
rect 17693 15317 17727 15351
rect 17727 15317 17736 15351
rect 17684 15308 17736 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 4068 15104 4120 15156
rect 5172 15147 5224 15156
rect 5172 15113 5181 15147
rect 5181 15113 5215 15147
rect 5215 15113 5224 15147
rect 5172 15104 5224 15113
rect 5356 15147 5408 15156
rect 5356 15113 5365 15147
rect 5365 15113 5399 15147
rect 5399 15113 5408 15147
rect 5356 15104 5408 15113
rect 6000 15104 6052 15156
rect 6828 15104 6880 15156
rect 7564 15104 7616 15156
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 9680 15147 9732 15156
rect 9680 15113 9689 15147
rect 9689 15113 9723 15147
rect 9723 15113 9732 15147
rect 9680 15104 9732 15113
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 4712 15079 4764 15088
rect 4712 15045 4721 15079
rect 4721 15045 4755 15079
rect 4755 15045 4764 15079
rect 4712 15036 4764 15045
rect 1584 14968 1636 15020
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 2412 14900 2464 14952
rect 5264 14968 5316 15020
rect 7012 15011 7064 15020
rect 7012 14977 7021 15011
rect 7021 14977 7055 15011
rect 7055 14977 7064 15011
rect 7012 14968 7064 14977
rect 7288 14968 7340 15020
rect 8116 15011 8168 15020
rect 8116 14977 8125 15011
rect 8125 14977 8159 15011
rect 8159 14977 8168 15011
rect 8116 14968 8168 14977
rect 9128 15036 9180 15088
rect 10876 15104 10928 15156
rect 14188 15104 14240 15156
rect 14648 15147 14700 15156
rect 14648 15113 14657 15147
rect 14657 15113 14691 15147
rect 14691 15113 14700 15147
rect 14648 15104 14700 15113
rect 16856 15104 16908 15156
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 4160 14900 4212 14952
rect 4804 14900 4856 14952
rect 6828 14900 6880 14952
rect 6920 14900 6972 14952
rect 7748 14900 7800 14952
rect 8208 14900 8260 14952
rect 9128 14900 9180 14952
rect 9496 15011 9548 15020
rect 9496 14977 9505 15011
rect 9505 14977 9539 15011
rect 9539 14977 9548 15011
rect 9496 14968 9548 14977
rect 9680 14968 9732 15020
rect 9864 14968 9916 15020
rect 12532 15036 12584 15088
rect 848 14764 900 14816
rect 2872 14807 2924 14816
rect 2872 14773 2881 14807
rect 2881 14773 2915 14807
rect 2915 14773 2924 14807
rect 2872 14764 2924 14773
rect 3424 14764 3476 14816
rect 3608 14764 3660 14816
rect 5356 14832 5408 14884
rect 5724 14832 5776 14884
rect 6552 14832 6604 14884
rect 6736 14764 6788 14816
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 7380 14832 7432 14884
rect 7748 14764 7800 14816
rect 9312 14832 9364 14884
rect 10324 15011 10376 15020
rect 10324 14977 10333 15011
rect 10333 14977 10367 15011
rect 10367 14977 10376 15011
rect 10324 14968 10376 14977
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 12164 14968 12216 15020
rect 12808 14968 12860 15020
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 10692 14900 10744 14952
rect 11704 14900 11756 14952
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 10416 14764 10468 14816
rect 11060 14764 11112 14816
rect 12164 14832 12216 14884
rect 13452 14900 13504 14952
rect 14372 14968 14424 15020
rect 14464 14943 14516 14952
rect 14464 14909 14473 14943
rect 14473 14909 14507 14943
rect 14507 14909 14516 14943
rect 14464 14900 14516 14909
rect 14924 14968 14976 15020
rect 16028 14968 16080 15020
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 17000 15011
rect 16948 14968 17000 14977
rect 16764 14900 16816 14952
rect 12348 14764 12400 14816
rect 12624 14764 12676 14816
rect 15568 14832 15620 14884
rect 16672 14875 16724 14884
rect 16672 14841 16681 14875
rect 16681 14841 16715 14875
rect 16715 14841 16724 14875
rect 16672 14832 16724 14841
rect 14464 14764 14516 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 3332 14560 3384 14612
rect 1952 14492 2004 14544
rect 2504 14424 2556 14476
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 1860 14356 1912 14408
rect 2412 14399 2464 14408
rect 2136 14331 2188 14340
rect 2136 14297 2145 14331
rect 2145 14297 2179 14331
rect 2179 14297 2188 14331
rect 2136 14288 2188 14297
rect 2044 14220 2096 14272
rect 2412 14365 2421 14399
rect 2421 14365 2455 14399
rect 2455 14365 2464 14399
rect 2412 14356 2464 14365
rect 2872 14424 2924 14476
rect 3976 14492 4028 14544
rect 4436 14492 4488 14544
rect 4712 14603 4764 14612
rect 4712 14569 4721 14603
rect 4721 14569 4755 14603
rect 4755 14569 4764 14603
rect 4712 14560 4764 14569
rect 7288 14560 7340 14612
rect 4804 14492 4856 14544
rect 5356 14492 5408 14544
rect 3608 14467 3660 14476
rect 3608 14433 3617 14467
rect 3617 14433 3651 14467
rect 3651 14433 3660 14467
rect 3608 14424 3660 14433
rect 3792 14424 3844 14476
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 3056 14356 3108 14408
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 2872 14331 2924 14340
rect 2872 14297 2881 14331
rect 2881 14297 2915 14331
rect 2915 14297 2924 14331
rect 2872 14288 2924 14297
rect 3884 14288 3936 14340
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 2320 14263 2372 14272
rect 2320 14229 2329 14263
rect 2329 14229 2363 14263
rect 2363 14229 2372 14263
rect 2320 14220 2372 14229
rect 2596 14263 2648 14272
rect 2596 14229 2605 14263
rect 2605 14229 2639 14263
rect 2639 14229 2648 14263
rect 2596 14220 2648 14229
rect 7012 14424 7064 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 7472 14560 7524 14612
rect 10140 14560 10192 14612
rect 10968 14603 11020 14612
rect 10968 14569 10977 14603
rect 10977 14569 11011 14603
rect 11011 14569 11020 14603
rect 10968 14560 11020 14569
rect 12072 14603 12124 14612
rect 12072 14569 12081 14603
rect 12081 14569 12115 14603
rect 12115 14569 12124 14603
rect 12072 14560 12124 14569
rect 15384 14560 15436 14612
rect 16488 14560 16540 14612
rect 17868 14603 17920 14612
rect 17868 14569 17877 14603
rect 17877 14569 17911 14603
rect 17911 14569 17920 14603
rect 17868 14560 17920 14569
rect 8484 14535 8536 14544
rect 8484 14501 8493 14535
rect 8493 14501 8527 14535
rect 8527 14501 8536 14535
rect 8484 14492 8536 14501
rect 11612 14492 11664 14544
rect 12808 14492 12860 14544
rect 14832 14535 14884 14544
rect 14832 14501 14841 14535
rect 14841 14501 14875 14535
rect 14875 14501 14884 14535
rect 14832 14492 14884 14501
rect 4436 14399 4488 14408
rect 4436 14365 4445 14399
rect 4445 14365 4479 14399
rect 4479 14365 4488 14399
rect 4436 14356 4488 14365
rect 4804 14356 4856 14408
rect 5632 14288 5684 14340
rect 6000 14399 6052 14408
rect 6000 14365 6009 14399
rect 6009 14365 6043 14399
rect 6043 14365 6052 14399
rect 6000 14356 6052 14365
rect 7472 14356 7524 14408
rect 4528 14263 4580 14272
rect 4528 14229 4537 14263
rect 4537 14229 4571 14263
rect 4571 14229 4580 14263
rect 4528 14220 4580 14229
rect 5264 14220 5316 14272
rect 6092 14263 6144 14272
rect 6092 14229 6101 14263
rect 6101 14229 6135 14263
rect 6135 14229 6144 14263
rect 6092 14220 6144 14229
rect 6460 14220 6512 14272
rect 6736 14220 6788 14272
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 8484 14356 8536 14408
rect 12992 14424 13044 14476
rect 8760 14356 8812 14408
rect 9496 14356 9548 14408
rect 9036 14331 9088 14340
rect 9036 14297 9045 14331
rect 9045 14297 9079 14331
rect 9079 14297 9088 14331
rect 9036 14288 9088 14297
rect 9956 14288 10008 14340
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 10508 14399 10560 14408
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 11336 14356 11388 14408
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 12348 14356 12400 14408
rect 12624 14399 12676 14408
rect 12624 14365 12633 14399
rect 12633 14365 12667 14399
rect 12667 14365 12676 14399
rect 12624 14356 12676 14365
rect 12808 14356 12860 14408
rect 16580 14424 16632 14476
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 10968 14331 11020 14340
rect 10968 14297 10977 14331
rect 10977 14297 11011 14331
rect 11011 14297 11020 14331
rect 10968 14288 11020 14297
rect 11152 14288 11204 14340
rect 14096 14288 14148 14340
rect 15016 14331 15068 14340
rect 15016 14297 15025 14331
rect 15025 14297 15059 14331
rect 15059 14297 15068 14331
rect 15016 14288 15068 14297
rect 16580 14288 16632 14340
rect 17960 14288 18012 14340
rect 8484 14220 8536 14272
rect 8852 14220 8904 14272
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 9220 14220 9272 14272
rect 11428 14220 11480 14272
rect 11520 14220 11572 14272
rect 13176 14220 13228 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 3148 14016 3200 14068
rect 2136 13948 2188 14000
rect 2412 13991 2464 14000
rect 2412 13957 2421 13991
rect 2421 13957 2455 13991
rect 2455 13957 2464 13991
rect 2412 13948 2464 13957
rect 2964 13948 3016 14000
rect 2320 13880 2372 13932
rect 3240 13948 3292 14000
rect 1860 13812 1912 13864
rect 2044 13812 2096 13864
rect 2596 13812 2648 13864
rect 3332 13923 3384 13932
rect 3332 13889 3341 13923
rect 3341 13889 3375 13923
rect 3375 13889 3384 13923
rect 3332 13880 3384 13889
rect 3516 13880 3568 13932
rect 3884 13923 3936 13932
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 4068 13923 4120 13932
rect 4068 13889 4077 13923
rect 4077 13889 4111 13923
rect 4111 13889 4120 13923
rect 4068 13880 4120 13889
rect 4712 13948 4764 14000
rect 6276 14016 6328 14068
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 6828 14016 6880 14068
rect 7196 14016 7248 14068
rect 8116 14016 8168 14068
rect 8300 14016 8352 14068
rect 9864 14016 9916 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 10508 14016 10560 14068
rect 11612 14059 11664 14068
rect 11612 14025 11621 14059
rect 11621 14025 11655 14059
rect 11655 14025 11664 14059
rect 11612 14016 11664 14025
rect 12072 14016 12124 14068
rect 12348 14016 12400 14068
rect 12900 14059 12952 14068
rect 12900 14025 12909 14059
rect 12909 14025 12943 14059
rect 12943 14025 12952 14059
rect 12900 14016 12952 14025
rect 13912 14016 13964 14068
rect 14280 14059 14332 14068
rect 14280 14025 14289 14059
rect 14289 14025 14323 14059
rect 14323 14025 14332 14059
rect 14280 14016 14332 14025
rect 16212 14016 16264 14068
rect 17776 14059 17828 14068
rect 17776 14025 17785 14059
rect 17785 14025 17819 14059
rect 17819 14025 17828 14059
rect 17776 14016 17828 14025
rect 1676 13676 1728 13728
rect 3608 13812 3660 13864
rect 4528 13880 4580 13932
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 6000 13880 6052 13932
rect 6736 13991 6788 14000
rect 6736 13957 6745 13991
rect 6745 13957 6779 13991
rect 6779 13957 6788 13991
rect 6736 13948 6788 13957
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 8484 13948 8536 14000
rect 4712 13812 4764 13864
rect 4804 13744 4856 13796
rect 5632 13812 5684 13864
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 6092 13812 6144 13864
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 7748 13880 7800 13932
rect 8116 13880 8168 13932
rect 12256 13948 12308 14000
rect 13176 13948 13228 14000
rect 16396 13948 16448 14000
rect 18052 13991 18104 14000
rect 18052 13957 18061 13991
rect 18061 13957 18095 13991
rect 18095 13957 18104 13991
rect 18052 13948 18104 13957
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 9128 13880 9180 13932
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 9956 13880 10008 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10784 13880 10836 13932
rect 11060 13923 11112 13932
rect 11060 13889 11069 13923
rect 11069 13889 11103 13923
rect 11103 13889 11112 13923
rect 11060 13880 11112 13889
rect 11520 13923 11572 13932
rect 7564 13812 7616 13864
rect 5816 13676 5868 13728
rect 6368 13676 6420 13728
rect 6920 13744 6972 13796
rect 6828 13676 6880 13728
rect 8024 13744 8076 13796
rect 9864 13744 9916 13796
rect 10232 13744 10284 13796
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 12624 13880 12676 13932
rect 12348 13855 12400 13864
rect 12348 13821 12357 13855
rect 12357 13821 12391 13855
rect 12391 13821 12400 13855
rect 12348 13812 12400 13821
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 14004 13923 14056 13932
rect 14004 13889 14013 13923
rect 14013 13889 14047 13923
rect 14047 13889 14056 13923
rect 14004 13880 14056 13889
rect 14464 13880 14516 13932
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 14924 13812 14976 13864
rect 15016 13812 15068 13864
rect 16764 13923 16816 13932
rect 16764 13889 16773 13923
rect 16773 13889 16807 13923
rect 16807 13889 16816 13923
rect 16764 13880 16816 13889
rect 16856 13812 16908 13864
rect 12440 13744 12492 13796
rect 13084 13744 13136 13796
rect 13820 13744 13872 13796
rect 13912 13744 13964 13796
rect 14556 13744 14608 13796
rect 15568 13744 15620 13796
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 7288 13676 7340 13685
rect 8300 13676 8352 13728
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 12164 13676 12216 13728
rect 12348 13676 12400 13728
rect 12624 13676 12676 13728
rect 13636 13676 13688 13728
rect 14464 13676 14516 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 1308 13472 1360 13524
rect 2412 13515 2464 13524
rect 2412 13481 2421 13515
rect 2421 13481 2455 13515
rect 2455 13481 2464 13515
rect 2412 13472 2464 13481
rect 3148 13472 3200 13524
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 3792 13336 3844 13388
rect 3976 13336 4028 13388
rect 4712 13404 4764 13456
rect 3148 13268 3200 13320
rect 3240 13268 3292 13320
rect 4804 13336 4856 13388
rect 5448 13336 5500 13388
rect 6000 13515 6052 13524
rect 6000 13481 6009 13515
rect 6009 13481 6043 13515
rect 6043 13481 6052 13515
rect 6000 13472 6052 13481
rect 6920 13472 6972 13524
rect 8760 13515 8812 13524
rect 8760 13481 8769 13515
rect 8769 13481 8803 13515
rect 8803 13481 8812 13515
rect 8760 13472 8812 13481
rect 9036 13472 9088 13524
rect 9772 13472 9824 13524
rect 10324 13472 10376 13524
rect 6276 13404 6328 13456
rect 8208 13404 8260 13456
rect 6460 13336 6512 13388
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 2780 13243 2832 13252
rect 2780 13209 2789 13243
rect 2789 13209 2823 13243
rect 2823 13209 2832 13243
rect 2780 13200 2832 13209
rect 3516 13200 3568 13252
rect 3700 13200 3752 13252
rect 3976 13200 4028 13252
rect 6092 13268 6144 13320
rect 4712 13200 4764 13252
rect 6368 13268 6420 13320
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 9220 13336 9272 13388
rect 9588 13268 9640 13320
rect 10416 13404 10468 13456
rect 10048 13268 10100 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 12440 13336 12492 13388
rect 9772 13243 9824 13252
rect 9772 13209 9781 13243
rect 9781 13209 9815 13243
rect 9815 13209 9824 13243
rect 9772 13200 9824 13209
rect 5080 13132 5132 13184
rect 5908 13132 5960 13184
rect 8300 13132 8352 13184
rect 9128 13132 9180 13184
rect 9220 13132 9272 13184
rect 10876 13132 10928 13184
rect 11796 13132 11848 13184
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12256 13268 12308 13320
rect 13452 13336 13504 13388
rect 13268 13268 13320 13320
rect 13820 13404 13872 13456
rect 15660 13404 15712 13456
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 16948 13336 17000 13388
rect 16488 13268 16540 13320
rect 12164 13132 12216 13184
rect 15016 13200 15068 13252
rect 12716 13132 12768 13184
rect 13544 13132 13596 13184
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 14004 13132 14056 13184
rect 15292 13132 15344 13184
rect 15844 13132 15896 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 4620 12928 4672 12980
rect 5172 12928 5224 12980
rect 6460 12928 6512 12980
rect 8024 12928 8076 12980
rect 8576 12971 8628 12980
rect 8576 12937 8585 12971
rect 8585 12937 8619 12971
rect 8619 12937 8628 12971
rect 8576 12928 8628 12937
rect 2872 12860 2924 12912
rect 4712 12860 4764 12912
rect 3148 12792 3200 12844
rect 3332 12835 3384 12844
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 3608 12792 3660 12844
rect 3792 12792 3844 12844
rect 5816 12860 5868 12912
rect 6000 12792 6052 12844
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 5080 12724 5132 12776
rect 8576 12792 8628 12844
rect 9680 12928 9732 12980
rect 10048 12928 10100 12980
rect 10876 12928 10928 12980
rect 11060 12860 11112 12912
rect 12072 12860 12124 12912
rect 12348 12860 12400 12912
rect 13912 12971 13964 12980
rect 13912 12937 13921 12971
rect 13921 12937 13955 12971
rect 13955 12937 13964 12971
rect 13912 12928 13964 12937
rect 14832 12928 14884 12980
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 2964 12656 3016 12708
rect 3148 12588 3200 12640
rect 4068 12588 4120 12640
rect 4620 12588 4672 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 6092 12588 6144 12640
rect 7196 12588 7248 12640
rect 8300 12699 8352 12708
rect 8300 12665 8309 12699
rect 8309 12665 8343 12699
rect 8343 12665 8352 12699
rect 8300 12656 8352 12665
rect 8392 12656 8444 12708
rect 9404 12724 9456 12776
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 11336 12724 11388 12776
rect 12532 12724 12584 12776
rect 13268 12835 13320 12844
rect 13268 12801 13277 12835
rect 13277 12801 13311 12835
rect 13311 12801 13320 12835
rect 13268 12792 13320 12801
rect 14280 12860 14332 12912
rect 13912 12792 13964 12844
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13820 12724 13872 12776
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 15108 12860 15160 12912
rect 16764 12928 16816 12980
rect 17684 12860 17736 12912
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 16856 12792 16908 12844
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 14832 12724 14884 12776
rect 8760 12656 8812 12708
rect 9864 12656 9916 12708
rect 10416 12699 10468 12708
rect 10416 12665 10425 12699
rect 10425 12665 10459 12699
rect 10459 12665 10468 12699
rect 10416 12656 10468 12665
rect 10784 12656 10836 12708
rect 12072 12656 12124 12708
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 15476 12724 15528 12776
rect 14280 12588 14332 12640
rect 14556 12588 14608 12640
rect 14648 12588 14700 12640
rect 14924 12588 14976 12640
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 1952 12384 2004 12436
rect 2228 12384 2280 12436
rect 3332 12384 3384 12436
rect 3240 12316 3292 12368
rect 5264 12384 5316 12436
rect 7380 12384 7432 12436
rect 9036 12384 9088 12436
rect 10232 12384 10284 12436
rect 10600 12384 10652 12436
rect 4344 12316 4396 12368
rect 4436 12316 4488 12368
rect 4712 12316 4764 12368
rect 4988 12316 5040 12368
rect 2780 12248 2832 12300
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3332 12180 3384 12232
rect 4068 12248 4120 12300
rect 4252 12223 4304 12232
rect 4252 12189 4287 12223
rect 4287 12189 4304 12223
rect 4252 12180 4304 12189
rect 4620 12180 4672 12232
rect 5540 12248 5592 12300
rect 8760 12316 8812 12368
rect 12716 12384 12768 12436
rect 3884 12112 3936 12164
rect 4528 12112 4580 12164
rect 2688 12044 2740 12096
rect 3424 12044 3476 12096
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 5724 12180 5776 12232
rect 6000 12180 6052 12232
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 7196 12248 7248 12300
rect 7932 12248 7984 12300
rect 8944 12248 8996 12300
rect 9128 12291 9180 12300
rect 9128 12257 9137 12291
rect 9137 12257 9171 12291
rect 9171 12257 9180 12291
rect 9128 12248 9180 12257
rect 9220 12248 9272 12300
rect 6184 12155 6236 12164
rect 6184 12121 6193 12155
rect 6193 12121 6227 12155
rect 6227 12121 6236 12155
rect 6184 12112 6236 12121
rect 6368 12044 6420 12096
rect 6736 12044 6788 12096
rect 7104 12112 7156 12164
rect 7564 12112 7616 12164
rect 7748 12112 7800 12164
rect 8392 12180 8444 12232
rect 8852 12112 8904 12164
rect 8944 12155 8996 12164
rect 8944 12121 8953 12155
rect 8953 12121 8987 12155
rect 8987 12121 8996 12155
rect 8944 12112 8996 12121
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 11060 12248 11112 12300
rect 12164 12316 12216 12368
rect 12256 12316 12308 12368
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 9680 12155 9732 12164
rect 9680 12121 9689 12155
rect 9689 12121 9723 12155
rect 9723 12121 9732 12155
rect 9680 12112 9732 12121
rect 10232 12180 10284 12232
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 11888 12248 11940 12300
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 11980 12180 12032 12232
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 12440 12223 12492 12232
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 12440 12180 12492 12189
rect 13176 12248 13228 12300
rect 14096 12248 14148 12300
rect 14924 12316 14976 12368
rect 15200 12384 15252 12436
rect 15476 12316 15528 12368
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 15016 12248 15068 12300
rect 16672 12248 16724 12300
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15108 12180 15160 12232
rect 15384 12223 15436 12232
rect 15384 12189 15393 12223
rect 15393 12189 15427 12223
rect 15427 12189 15436 12223
rect 15384 12180 15436 12189
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 11888 12112 11940 12164
rect 12716 12155 12768 12164
rect 12716 12121 12725 12155
rect 12725 12121 12759 12155
rect 12759 12121 12768 12155
rect 12716 12112 12768 12121
rect 12992 12112 13044 12164
rect 14188 12112 14240 12164
rect 15844 12112 15896 12164
rect 16764 12112 16816 12164
rect 9864 12044 9916 12096
rect 10232 12044 10284 12096
rect 11980 12044 12032 12096
rect 14924 12044 14976 12096
rect 15200 12044 15252 12096
rect 17776 12087 17828 12096
rect 17776 12053 17785 12087
rect 17785 12053 17819 12087
rect 17819 12053 17828 12087
rect 17776 12044 17828 12053
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2412 11840 2464 11892
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 2688 11815 2740 11824
rect 2688 11781 2697 11815
rect 2697 11781 2731 11815
rect 2731 11781 2740 11815
rect 2688 11772 2740 11781
rect 3332 11772 3384 11824
rect 4344 11772 4396 11824
rect 5908 11840 5960 11892
rect 6276 11840 6328 11892
rect 6460 11840 6512 11892
rect 7564 11840 7616 11892
rect 7656 11840 7708 11892
rect 8116 11840 8168 11892
rect 9680 11840 9732 11892
rect 9864 11840 9916 11892
rect 1768 11636 1820 11688
rect 2780 11747 2832 11756
rect 2780 11713 2825 11747
rect 2825 11713 2832 11747
rect 2780 11704 2832 11713
rect 3148 11704 3200 11756
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 4436 11704 4488 11756
rect 4620 11704 4672 11756
rect 2872 11568 2924 11620
rect 4804 11636 4856 11688
rect 1676 11500 1728 11552
rect 4712 11500 4764 11552
rect 5172 11747 5224 11756
rect 5172 11713 5181 11747
rect 5181 11713 5215 11747
rect 5215 11713 5224 11747
rect 5172 11704 5224 11713
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 6276 11704 6328 11756
rect 6644 11747 6696 11756
rect 6644 11713 6653 11747
rect 6653 11713 6687 11747
rect 6687 11713 6696 11747
rect 6644 11704 6696 11713
rect 8392 11772 8444 11824
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 6552 11636 6604 11688
rect 7564 11636 7616 11688
rect 9864 11704 9916 11756
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 11244 11840 11296 11892
rect 11428 11840 11480 11892
rect 11520 11840 11572 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 11704 11772 11756 11824
rect 5816 11568 5868 11620
rect 6184 11568 6236 11620
rect 6920 11568 6972 11620
rect 5356 11500 5408 11552
rect 7932 11568 7984 11620
rect 7472 11500 7524 11552
rect 11152 11636 11204 11688
rect 11888 11704 11940 11756
rect 14188 11840 14240 11892
rect 15568 11840 15620 11892
rect 15844 11883 15896 11892
rect 15844 11849 15853 11883
rect 15853 11849 15887 11883
rect 15887 11849 15896 11883
rect 15844 11840 15896 11849
rect 13452 11772 13504 11824
rect 15200 11815 15252 11824
rect 15200 11781 15209 11815
rect 15209 11781 15243 11815
rect 15243 11781 15252 11815
rect 15200 11772 15252 11781
rect 15936 11772 15988 11824
rect 13268 11747 13320 11756
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 13360 11747 13412 11756
rect 13360 11713 13369 11747
rect 13369 11713 13403 11747
rect 13403 11713 13412 11747
rect 13360 11704 13412 11713
rect 13544 11747 13596 11756
rect 13544 11713 13553 11747
rect 13553 11713 13587 11747
rect 13587 11713 13596 11747
rect 13544 11704 13596 11713
rect 16120 11704 16172 11756
rect 11704 11636 11756 11688
rect 14832 11636 14884 11688
rect 11520 11500 11572 11552
rect 12164 11568 12216 11620
rect 13360 11568 13412 11620
rect 15108 11568 15160 11620
rect 15844 11679 15896 11688
rect 15844 11645 15853 11679
rect 15853 11645 15887 11679
rect 15887 11645 15896 11679
rect 15844 11636 15896 11645
rect 15936 11679 15988 11688
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 17776 11747 17828 11756
rect 17776 11713 17785 11747
rect 17785 11713 17819 11747
rect 17819 11713 17828 11747
rect 17776 11704 17828 11713
rect 16948 11568 17000 11620
rect 17776 11568 17828 11620
rect 12532 11500 12584 11552
rect 13728 11500 13780 11552
rect 16764 11500 16816 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1124 11296 1176 11348
rect 1860 11296 1912 11348
rect 3148 11296 3200 11348
rect 3884 11296 3936 11348
rect 3792 11228 3844 11280
rect 4620 11296 4672 11348
rect 5356 11296 5408 11348
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 2320 11092 2372 11144
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 2596 11092 2648 11101
rect 3792 11135 3844 11144
rect 3792 11101 3801 11135
rect 3801 11101 3835 11135
rect 3835 11101 3844 11135
rect 3792 11092 3844 11101
rect 4436 11135 4488 11144
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 6276 11092 6328 11144
rect 2412 11067 2464 11076
rect 2412 11033 2421 11067
rect 2421 11033 2455 11067
rect 2455 11033 2464 11067
rect 2412 11024 2464 11033
rect 2688 11024 2740 11076
rect 3240 11024 3292 11076
rect 4988 11024 5040 11076
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 7564 11296 7616 11348
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 7380 11271 7432 11280
rect 7380 11237 7389 11271
rect 7389 11237 7423 11271
rect 7423 11237 7432 11271
rect 7380 11228 7432 11237
rect 8392 11271 8444 11280
rect 8392 11237 8401 11271
rect 8401 11237 8435 11271
rect 8435 11237 8444 11271
rect 8392 11228 8444 11237
rect 7196 11092 7248 11144
rect 7288 11024 7340 11076
rect 8208 11092 8260 11144
rect 8300 11135 8352 11144
rect 8300 11101 8310 11135
rect 8310 11101 8344 11135
rect 8344 11101 8352 11135
rect 8300 11092 8352 11101
rect 2872 10956 2924 11008
rect 3884 10956 3936 11008
rect 5172 10956 5224 11008
rect 6368 10956 6420 11008
rect 6920 10956 6972 11008
rect 8116 10956 8168 11008
rect 8300 10956 8352 11008
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 9312 11296 9364 11348
rect 11704 11296 11756 11348
rect 12072 11296 12124 11348
rect 12440 11296 12492 11348
rect 14464 11296 14516 11348
rect 15844 11296 15896 11348
rect 16488 11296 16540 11348
rect 17224 11296 17276 11348
rect 9220 11228 9272 11280
rect 11520 11228 11572 11280
rect 8852 11092 8904 11144
rect 9496 11160 9548 11212
rect 10140 11160 10192 11212
rect 9588 11092 9640 11144
rect 9680 11092 9732 11144
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 11980 11160 12032 11212
rect 12440 11160 12492 11212
rect 12808 11160 12860 11212
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 10876 11092 10928 11144
rect 12716 11092 12768 11144
rect 13452 11092 13504 11144
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 14188 11092 14240 11144
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 15384 11092 15436 11144
rect 16028 11160 16080 11212
rect 18144 11203 18196 11212
rect 18144 11169 18153 11203
rect 18153 11169 18187 11203
rect 18187 11169 18196 11203
rect 18144 11160 18196 11169
rect 16120 11092 16172 11144
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 17960 11092 18012 11144
rect 14648 11024 14700 11076
rect 15568 11024 15620 11076
rect 9220 10999 9272 11008
rect 9220 10965 9229 10999
rect 9229 10965 9263 10999
rect 9263 10965 9272 10999
rect 9220 10956 9272 10965
rect 9772 10956 9824 11008
rect 9864 10956 9916 11008
rect 11796 10956 11848 11008
rect 14096 10956 14148 11008
rect 15660 10999 15712 11008
rect 15660 10965 15669 10999
rect 15669 10965 15703 10999
rect 15703 10965 15712 10999
rect 15660 10956 15712 10965
rect 16212 10956 16264 11008
rect 16672 11067 16724 11076
rect 16672 11033 16681 11067
rect 16681 11033 16715 11067
rect 16715 11033 16724 11067
rect 16672 11024 16724 11033
rect 17408 10956 17460 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 2136 10752 2188 10804
rect 2412 10752 2464 10804
rect 3700 10795 3752 10804
rect 3700 10761 3709 10795
rect 3709 10761 3743 10795
rect 3743 10761 3752 10795
rect 3700 10752 3752 10761
rect 4068 10752 4120 10804
rect 4620 10752 4672 10804
rect 5816 10752 5868 10804
rect 7748 10752 7800 10804
rect 4804 10684 4856 10736
rect 5172 10684 5224 10736
rect 3700 10616 3752 10668
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 3976 10616 4028 10668
rect 5264 10616 5316 10668
rect 5724 10616 5776 10668
rect 6552 10684 6604 10736
rect 6092 10616 6144 10668
rect 7656 10616 7708 10668
rect 9864 10752 9916 10804
rect 14188 10752 14240 10804
rect 14648 10752 14700 10804
rect 8116 10727 8168 10736
rect 8116 10693 8125 10727
rect 8125 10693 8159 10727
rect 8159 10693 8168 10727
rect 8116 10684 8168 10693
rect 3976 10412 4028 10464
rect 4620 10412 4672 10464
rect 5080 10591 5132 10600
rect 5080 10557 5089 10591
rect 5089 10557 5123 10591
rect 5123 10557 5132 10591
rect 5080 10548 5132 10557
rect 4988 10480 5040 10532
rect 6368 10548 6420 10600
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 7196 10548 7248 10600
rect 8392 10616 8444 10668
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 10232 10684 10284 10736
rect 15200 10752 15252 10804
rect 15384 10752 15436 10804
rect 16580 10752 16632 10804
rect 10876 10616 10928 10668
rect 8116 10480 8168 10532
rect 9128 10548 9180 10600
rect 9588 10548 9640 10600
rect 10692 10548 10744 10600
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 9036 10480 9088 10532
rect 11980 10548 12032 10600
rect 5540 10412 5592 10464
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 8392 10412 8444 10464
rect 10324 10412 10376 10464
rect 10508 10412 10560 10464
rect 13820 10548 13872 10600
rect 12164 10480 12216 10532
rect 15016 10727 15068 10736
rect 15016 10693 15025 10727
rect 15025 10693 15059 10727
rect 15059 10693 15068 10727
rect 15016 10684 15068 10693
rect 14556 10616 14608 10668
rect 16304 10684 16356 10736
rect 16396 10684 16448 10736
rect 15752 10616 15804 10668
rect 15384 10480 15436 10532
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 16212 10659 16264 10668
rect 16212 10625 16221 10659
rect 16221 10625 16255 10659
rect 16255 10625 16264 10659
rect 16212 10616 16264 10625
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17408 10727 17460 10736
rect 17408 10693 17417 10727
rect 17417 10693 17451 10727
rect 17451 10693 17460 10727
rect 17408 10684 17460 10693
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 14096 10412 14148 10421
rect 15016 10412 15068 10464
rect 15108 10412 15160 10464
rect 16212 10412 16264 10464
rect 16856 10548 16908 10600
rect 17684 10659 17736 10668
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 18052 10616 18104 10668
rect 17224 10548 17276 10600
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 2964 10208 3016 10260
rect 4988 10140 5040 10192
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2872 10004 2924 10056
rect 3792 10004 3844 10056
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4620 10072 4672 10124
rect 5172 10072 5224 10124
rect 5356 10072 5408 10124
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 5080 10004 5132 10056
rect 5724 10072 5776 10124
rect 9036 10208 9088 10260
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 9864 10208 9916 10260
rect 7104 10140 7156 10192
rect 7932 10140 7984 10192
rect 9220 10140 9272 10192
rect 6368 10004 6420 10056
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 5724 9979 5776 9988
rect 5724 9945 5733 9979
rect 5733 9945 5767 9979
rect 5767 9945 5776 9979
rect 5724 9936 5776 9945
rect 6552 9936 6604 9988
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 3056 9868 3108 9920
rect 5632 9868 5684 9920
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 9404 10072 9456 10124
rect 7380 9979 7432 9988
rect 7380 9945 7389 9979
rect 7389 9945 7423 9979
rect 7423 9945 7432 9979
rect 7380 9936 7432 9945
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 9864 10072 9916 10124
rect 11888 10208 11940 10260
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 15292 10208 15344 10260
rect 16212 10208 16264 10260
rect 16672 10208 16724 10260
rect 17040 10208 17092 10260
rect 10324 10072 10376 10124
rect 10692 10072 10744 10124
rect 9956 10004 10008 10056
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 15200 10140 15252 10192
rect 16120 10140 16172 10192
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 11796 10004 11848 10056
rect 15660 10072 15712 10124
rect 15568 10047 15620 10056
rect 15568 10013 15581 10047
rect 15581 10013 15620 10047
rect 8484 9936 8536 9988
rect 8576 9936 8628 9988
rect 9864 9979 9916 9988
rect 9864 9945 9873 9979
rect 9873 9945 9907 9979
rect 9907 9945 9916 9979
rect 9864 9936 9916 9945
rect 11060 9936 11112 9988
rect 15568 10004 15620 10013
rect 13912 9936 13964 9988
rect 14096 9936 14148 9988
rect 16488 10047 16540 10056
rect 8116 9868 8168 9920
rect 9404 9868 9456 9920
rect 10140 9868 10192 9920
rect 10324 9911 10376 9920
rect 10324 9877 10333 9911
rect 10333 9877 10367 9911
rect 10367 9877 10376 9911
rect 10324 9868 10376 9877
rect 10508 9868 10560 9920
rect 10968 9868 11020 9920
rect 12808 9868 12860 9920
rect 13084 9868 13136 9920
rect 16488 10013 16497 10047
rect 16497 10013 16531 10047
rect 16531 10013 16540 10047
rect 16488 10004 16540 10013
rect 16672 10072 16724 10124
rect 16948 10004 17000 10056
rect 16028 9979 16080 9988
rect 16028 9945 16037 9979
rect 16037 9945 16071 9979
rect 16071 9945 16080 9979
rect 16028 9936 16080 9945
rect 16120 9936 16172 9988
rect 16304 9936 16356 9988
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 17592 10004 17644 10056
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 17040 9868 17092 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1676 9664 1728 9716
rect 2320 9639 2372 9648
rect 2320 9605 2329 9639
rect 2329 9605 2363 9639
rect 2363 9605 2372 9639
rect 2320 9596 2372 9605
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2412 9528 2464 9580
rect 3608 9596 3660 9648
rect 5080 9664 5132 9716
rect 5540 9664 5592 9716
rect 5724 9664 5776 9716
rect 2596 9528 2648 9580
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 2964 9528 3016 9580
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3700 9528 3752 9580
rect 4068 9596 4120 9648
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 5632 9596 5684 9648
rect 7012 9664 7064 9716
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 6368 9528 6420 9580
rect 6736 9596 6788 9648
rect 2136 9503 2188 9512
rect 2136 9469 2145 9503
rect 2145 9469 2179 9503
rect 2179 9469 2188 9503
rect 2136 9460 2188 9469
rect 5264 9460 5316 9512
rect 6644 9503 6696 9546
rect 6644 9494 6653 9503
rect 6653 9494 6687 9503
rect 6687 9494 6696 9503
rect 6736 9503 6788 9546
rect 6736 9494 6745 9503
rect 6745 9494 6779 9503
rect 6779 9494 6788 9503
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7748 9664 7800 9716
rect 9496 9664 9548 9716
rect 10232 9664 10284 9716
rect 12992 9664 13044 9716
rect 13360 9664 13412 9716
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 8208 9528 8260 9580
rect 9220 9528 9272 9580
rect 9588 9571 9640 9580
rect 9588 9537 9597 9571
rect 9597 9537 9631 9571
rect 9631 9537 9640 9571
rect 9588 9528 9640 9537
rect 10048 9596 10100 9648
rect 12256 9596 12308 9648
rect 10416 9528 10468 9580
rect 11060 9571 11112 9580
rect 11060 9537 11069 9571
rect 11069 9537 11103 9571
rect 11103 9537 11112 9571
rect 11060 9528 11112 9537
rect 11888 9528 11940 9580
rect 12440 9528 12492 9580
rect 12716 9571 12768 9580
rect 12716 9537 12737 9571
rect 12737 9537 12768 9571
rect 12716 9528 12768 9537
rect 13084 9518 13136 9570
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 2964 9324 3016 9376
rect 4344 9392 4396 9444
rect 6092 9392 6144 9444
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 8576 9460 8628 9512
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 8116 9392 8168 9444
rect 5172 9324 5224 9376
rect 5724 9324 5776 9376
rect 5908 9324 5960 9376
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8392 9324 8444 9376
rect 9588 9324 9640 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 9956 9392 10008 9444
rect 10416 9392 10468 9444
rect 11152 9392 11204 9444
rect 12164 9392 12216 9444
rect 12808 9392 12860 9444
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 14004 9528 14056 9580
rect 16856 9596 16908 9648
rect 14924 9528 14976 9580
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 18144 9596 18196 9648
rect 18052 9528 18104 9580
rect 13360 9392 13412 9444
rect 11520 9324 11572 9376
rect 12532 9324 12584 9376
rect 12716 9367 12768 9376
rect 12716 9333 12725 9367
rect 12725 9333 12759 9367
rect 12759 9333 12768 9367
rect 12716 9324 12768 9333
rect 12992 9324 13044 9376
rect 13636 9324 13688 9376
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 17316 9460 17368 9512
rect 17500 9503 17552 9512
rect 17500 9469 17509 9503
rect 17509 9469 17543 9503
rect 17543 9469 17552 9503
rect 17500 9460 17552 9469
rect 16028 9392 16080 9444
rect 17776 9324 17828 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 1860 9120 1912 9172
rect 2044 9120 2096 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 3884 9163 3936 9172
rect 3884 9129 3893 9163
rect 3893 9129 3927 9163
rect 3927 9129 3936 9163
rect 3884 9120 3936 9129
rect 4620 9120 4672 9172
rect 4988 9120 5040 9172
rect 5356 9120 5408 9172
rect 5724 9120 5776 9172
rect 7472 9120 7524 9172
rect 6736 9052 6788 9104
rect 1768 8848 1820 8900
rect 2228 8916 2280 8968
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 2412 8916 2464 8968
rect 2964 8984 3016 9036
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3424 8916 3476 8968
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 4068 8984 4120 8993
rect 4528 8984 4580 9036
rect 3792 8916 3844 8968
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 4344 8959 4396 8968
rect 4344 8925 4353 8959
rect 4353 8925 4387 8959
rect 4387 8925 4396 8959
rect 4344 8916 4396 8925
rect 4896 8984 4948 9036
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 5172 8916 5224 8968
rect 5632 8916 5684 8968
rect 6000 8916 6052 8968
rect 6828 8916 6880 8968
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 7288 9052 7340 9104
rect 8024 9120 8076 9172
rect 8668 9120 8720 9172
rect 9312 9120 9364 9172
rect 10692 9120 10744 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 9404 9052 9456 9104
rect 12532 9120 12584 9172
rect 13452 9120 13504 9172
rect 14188 9120 14240 9172
rect 15568 9120 15620 9172
rect 16304 9120 16356 9172
rect 16580 9120 16632 9172
rect 16856 9120 16908 9172
rect 11336 9052 11388 9104
rect 11980 9052 12032 9104
rect 12164 9052 12216 9104
rect 13360 9052 13412 9104
rect 7840 8984 7892 9036
rect 7932 8916 7984 8968
rect 4712 8848 4764 8900
rect 2320 8780 2372 8832
rect 3608 8823 3660 8832
rect 3608 8789 3617 8823
rect 3617 8789 3651 8823
rect 3651 8789 3660 8823
rect 3608 8780 3660 8789
rect 3884 8780 3936 8832
rect 5724 8780 5776 8832
rect 6000 8780 6052 8832
rect 6184 8891 6236 8900
rect 6184 8857 6193 8891
rect 6193 8857 6227 8891
rect 6227 8857 6236 8891
rect 6184 8848 6236 8857
rect 7472 8891 7524 8900
rect 7472 8857 7481 8891
rect 7481 8857 7515 8891
rect 7515 8857 7524 8891
rect 7472 8848 7524 8857
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9404 8916 9456 8968
rect 6368 8780 6420 8832
rect 7932 8780 7984 8832
rect 9588 8848 9640 8900
rect 9956 8959 10008 8968
rect 9956 8925 9965 8959
rect 9965 8925 9999 8959
rect 9999 8925 10008 8959
rect 9956 8916 10008 8925
rect 10140 8916 10192 8968
rect 12256 8984 12308 9036
rect 12532 8984 12584 9036
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 16672 9052 16724 9104
rect 17684 9052 17736 9104
rect 16212 9027 16264 9036
rect 16212 8993 16221 9027
rect 16221 8993 16255 9027
rect 16255 8993 16264 9027
rect 16212 8984 16264 8993
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 11060 8848 11112 8900
rect 8760 8780 8812 8832
rect 9956 8780 10008 8832
rect 10324 8780 10376 8832
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 11152 8780 11204 8832
rect 13084 8916 13136 8968
rect 14188 8916 14240 8968
rect 14372 8916 14424 8968
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 15476 8959 15528 8968
rect 15476 8925 15485 8959
rect 15485 8925 15519 8959
rect 15519 8925 15528 8959
rect 15476 8916 15528 8925
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 15844 8916 15896 8968
rect 16396 8959 16448 8968
rect 16396 8925 16405 8959
rect 16405 8925 16439 8959
rect 16439 8925 16448 8959
rect 16396 8916 16448 8925
rect 17408 8984 17460 9036
rect 11980 8780 12032 8832
rect 16212 8848 16264 8900
rect 12900 8780 12952 8832
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 14832 8780 14884 8832
rect 16580 8780 16632 8832
rect 17132 8916 17184 8968
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 17316 8780 17368 8832
rect 17592 8780 17644 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 4160 8576 4212 8628
rect 4988 8576 5040 8628
rect 5540 8576 5592 8628
rect 8760 8576 8812 8628
rect 9312 8576 9364 8628
rect 9864 8576 9916 8628
rect 11152 8576 11204 8628
rect 12992 8576 13044 8628
rect 14188 8576 14240 8628
rect 14740 8576 14792 8628
rect 15108 8576 15160 8628
rect 7104 8508 7156 8560
rect 7288 8508 7340 8560
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4068 8415 4120 8424
rect 4068 8381 4077 8415
rect 4077 8381 4111 8415
rect 4111 8381 4120 8415
rect 4068 8372 4120 8381
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5264 8440 5316 8492
rect 6368 8440 6420 8492
rect 5172 8372 5224 8424
rect 6920 8440 6972 8492
rect 7748 8440 7800 8492
rect 8392 8508 8444 8560
rect 8944 8508 8996 8560
rect 9036 8551 9088 8560
rect 9036 8517 9045 8551
rect 9045 8517 9079 8551
rect 9079 8517 9088 8551
rect 9036 8508 9088 8517
rect 9588 8508 9640 8560
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 4712 8304 4764 8356
rect 6368 8347 6420 8356
rect 6368 8313 6377 8347
rect 6377 8313 6411 8347
rect 6411 8313 6420 8347
rect 6368 8304 6420 8313
rect 3516 8236 3568 8288
rect 4988 8236 5040 8288
rect 5540 8236 5592 8288
rect 5908 8236 5960 8288
rect 6644 8236 6696 8288
rect 7564 8372 7616 8424
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 11520 8508 11572 8560
rect 15200 8508 15252 8560
rect 8944 8372 8996 8424
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10048 8440 10100 8492
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10508 8440 10560 8492
rect 8116 8347 8168 8356
rect 8116 8313 8125 8347
rect 8125 8313 8159 8347
rect 8159 8313 8168 8347
rect 8116 8304 8168 8313
rect 8208 8304 8260 8356
rect 8392 8304 8444 8356
rect 8576 8304 8628 8356
rect 9036 8304 9088 8356
rect 10416 8304 10468 8356
rect 10692 8440 10744 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 11428 8440 11480 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 12348 8440 12400 8492
rect 12532 8440 12584 8492
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13912 8440 13964 8492
rect 13084 8372 13136 8424
rect 13544 8372 13596 8424
rect 14280 8440 14332 8492
rect 14832 8440 14884 8492
rect 15660 8576 15712 8628
rect 15936 8576 15988 8628
rect 16212 8576 16264 8628
rect 16672 8576 16724 8628
rect 15568 8483 15620 8492
rect 15568 8449 15577 8483
rect 15577 8449 15611 8483
rect 15611 8449 15620 8483
rect 15568 8440 15620 8449
rect 15752 8440 15804 8492
rect 14372 8372 14424 8424
rect 16028 8372 16080 8424
rect 11612 8304 11664 8356
rect 7288 8236 7340 8288
rect 7748 8236 7800 8288
rect 8300 8236 8352 8288
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 12900 8347 12952 8356
rect 12900 8313 12909 8347
rect 12909 8313 12943 8347
rect 12943 8313 12952 8347
rect 12900 8304 12952 8313
rect 13728 8304 13780 8356
rect 14556 8304 14608 8356
rect 15660 8304 15712 8356
rect 16580 8440 16632 8492
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 16856 8372 16908 8424
rect 15384 8236 15436 8288
rect 16028 8236 16080 8288
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 16856 8236 16908 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 1676 8032 1728 8084
rect 3700 8032 3752 8084
rect 4988 8032 5040 8084
rect 8944 8032 8996 8084
rect 9588 8075 9640 8084
rect 9588 8041 9597 8075
rect 9597 8041 9631 8075
rect 9631 8041 9640 8075
rect 9588 8032 9640 8041
rect 10232 8032 10284 8084
rect 11336 8032 11388 8084
rect 11520 8032 11572 8084
rect 11704 8032 11756 8084
rect 12164 8032 12216 8084
rect 1952 7939 2004 7948
rect 1952 7905 1961 7939
rect 1961 7905 1995 7939
rect 1995 7905 2004 7939
rect 1952 7896 2004 7905
rect 1768 7828 1820 7880
rect 3884 7828 3936 7880
rect 4712 7896 4764 7948
rect 4804 7896 4856 7948
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 4896 7828 4948 7880
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 5632 7828 5684 7880
rect 5817 7871 5869 7880
rect 5817 7837 5826 7871
rect 5826 7837 5860 7871
rect 5860 7837 5869 7871
rect 5817 7828 5869 7837
rect 6092 7939 6144 7948
rect 6092 7905 6101 7939
rect 6101 7905 6135 7939
rect 6135 7905 6144 7939
rect 6092 7896 6144 7905
rect 6276 7896 6328 7948
rect 3608 7760 3660 7812
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 6828 7896 6880 7948
rect 8668 7964 8720 8016
rect 7104 7828 7156 7880
rect 6828 7803 6880 7812
rect 6828 7769 6837 7803
rect 6837 7769 6871 7803
rect 6871 7769 6880 7803
rect 6828 7760 6880 7769
rect 7288 7830 7340 7882
rect 7472 7871 7524 7882
rect 7472 7837 7487 7871
rect 7487 7837 7521 7871
rect 7521 7837 7524 7871
rect 7472 7830 7524 7837
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 8300 7871 8352 7880
rect 7748 7760 7800 7812
rect 8116 7849 8168 7858
rect 8116 7815 8125 7849
rect 8125 7815 8159 7849
rect 8159 7815 8168 7849
rect 8116 7806 8168 7815
rect 8300 7837 8321 7871
rect 8321 7837 8352 7871
rect 8300 7828 8352 7837
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 10784 7964 10836 8016
rect 12716 7964 12768 8016
rect 12900 8032 12952 8084
rect 17500 8032 17552 8084
rect 11704 7939 11756 7948
rect 11704 7905 11713 7939
rect 11713 7905 11747 7939
rect 11747 7905 11756 7939
rect 11704 7896 11756 7905
rect 8852 7828 8904 7880
rect 9036 7828 9088 7880
rect 9496 7828 9548 7880
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 10048 7828 10100 7880
rect 11244 7828 11296 7880
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 10324 7760 10376 7812
rect 10692 7760 10744 7812
rect 10876 7760 10928 7812
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 12900 7760 12952 7812
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 4804 7692 4856 7744
rect 5172 7692 5224 7744
rect 7656 7692 7708 7744
rect 8208 7692 8260 7744
rect 8944 7692 8996 7744
rect 10416 7692 10468 7744
rect 12164 7692 12216 7744
rect 12256 7692 12308 7744
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 15016 7939 15068 7948
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 15384 7964 15436 8016
rect 16120 7964 16172 8016
rect 14832 7871 14884 7880
rect 14832 7837 14841 7871
rect 14841 7837 14875 7871
rect 14875 7837 14884 7871
rect 14832 7828 14884 7837
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 16672 7896 16724 7948
rect 13544 7803 13596 7812
rect 13544 7769 13553 7803
rect 13553 7769 13587 7803
rect 13587 7769 13596 7803
rect 13544 7760 13596 7769
rect 13636 7760 13688 7812
rect 14372 7803 14424 7812
rect 14372 7769 14381 7803
rect 14381 7769 14415 7803
rect 14415 7769 14424 7803
rect 14372 7760 14424 7769
rect 15016 7760 15068 7812
rect 15844 7803 15896 7812
rect 15844 7769 15853 7803
rect 15853 7769 15887 7803
rect 15887 7769 15896 7803
rect 15844 7760 15896 7769
rect 16304 7760 16356 7812
rect 16856 7803 16908 7812
rect 16856 7769 16865 7803
rect 16865 7769 16899 7803
rect 16899 7769 16908 7803
rect 16856 7760 16908 7769
rect 14740 7692 14792 7744
rect 15384 7735 15436 7744
rect 15384 7701 15393 7735
rect 15393 7701 15427 7735
rect 15427 7701 15436 7735
rect 15384 7692 15436 7701
rect 17132 7692 17184 7744
rect 17592 7692 17644 7744
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1768 7488 1820 7540
rect 3424 7488 3476 7540
rect 3792 7488 3844 7540
rect 4436 7488 4488 7540
rect 1952 7352 2004 7404
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 2596 7352 2648 7361
rect 2872 7352 2924 7404
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3056 7352 3108 7361
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 3516 7284 3568 7336
rect 4436 7352 4488 7404
rect 5448 7488 5500 7540
rect 6000 7488 6052 7540
rect 6828 7488 6880 7540
rect 7288 7488 7340 7540
rect 9956 7488 10008 7540
rect 10232 7488 10284 7540
rect 11796 7488 11848 7540
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 13820 7488 13872 7540
rect 14372 7488 14424 7540
rect 14832 7488 14884 7540
rect 15200 7531 15252 7540
rect 15200 7497 15209 7531
rect 15209 7497 15243 7531
rect 15243 7497 15252 7531
rect 15200 7488 15252 7497
rect 15384 7488 15436 7540
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5264 7284 5316 7336
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 6092 7420 6144 7472
rect 10508 7420 10560 7472
rect 12532 7420 12584 7472
rect 12900 7420 12952 7472
rect 6276 7352 6328 7404
rect 8760 7352 8812 7404
rect 9036 7352 9088 7404
rect 10048 7352 10100 7404
rect 11244 7352 11296 7404
rect 7564 7284 7616 7336
rect 6460 7216 6512 7268
rect 10140 7284 10192 7336
rect 10232 7216 10284 7268
rect 10692 7216 10744 7268
rect 13544 7284 13596 7336
rect 14556 7216 14608 7268
rect 14740 7259 14792 7268
rect 14740 7225 14749 7259
rect 14749 7225 14783 7259
rect 14783 7225 14792 7259
rect 14740 7216 14792 7225
rect 15292 7352 15344 7404
rect 15936 7284 15988 7336
rect 1676 7148 1728 7200
rect 2504 7148 2556 7200
rect 3884 7148 3936 7200
rect 4804 7148 4856 7200
rect 5540 7148 5592 7200
rect 7656 7148 7708 7200
rect 9036 7148 9088 7200
rect 9956 7148 10008 7200
rect 10508 7148 10560 7200
rect 10968 7148 11020 7200
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 13360 7148 13412 7200
rect 15568 7216 15620 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3332 6944 3384 6996
rect 5540 6944 5592 6996
rect 6184 6944 6236 6996
rect 7380 6944 7432 6996
rect 9680 6944 9732 6996
rect 10692 6987 10744 6996
rect 10692 6953 10701 6987
rect 10701 6953 10735 6987
rect 10735 6953 10744 6987
rect 10692 6944 10744 6953
rect 10968 6987 11020 6996
rect 10968 6953 10977 6987
rect 10977 6953 11011 6987
rect 11011 6953 11020 6987
rect 10968 6944 11020 6953
rect 11060 6944 11112 6996
rect 3148 6808 3200 6860
rect 4528 6808 4580 6860
rect 5724 6808 5776 6860
rect 8208 6808 8260 6860
rect 9772 6851 9824 6860
rect 9772 6817 9781 6851
rect 9781 6817 9815 6851
rect 9815 6817 9824 6851
rect 9772 6808 9824 6817
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2504 6783 2556 6792
rect 2504 6749 2513 6783
rect 2513 6749 2547 6783
rect 2547 6749 2556 6783
rect 2504 6740 2556 6749
rect 3792 6740 3844 6792
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 4436 6672 4488 6724
rect 4712 6672 4764 6724
rect 4988 6740 5040 6792
rect 5264 6740 5316 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 6000 6740 6052 6792
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 8300 6740 8352 6792
rect 9496 6740 9548 6792
rect 10416 6876 10468 6928
rect 13084 6944 13136 6996
rect 13452 6944 13504 6996
rect 11428 6876 11480 6928
rect 13544 6876 13596 6928
rect 14004 6876 14056 6928
rect 14372 6808 14424 6860
rect 15016 6808 15068 6860
rect 15200 6876 15252 6928
rect 16488 6876 16540 6928
rect 9588 6672 9640 6724
rect 10416 6783 10468 6792
rect 10416 6749 10428 6783
rect 10428 6749 10462 6783
rect 10462 6749 10468 6783
rect 10416 6740 10468 6749
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11060 6740 11112 6792
rect 10232 6672 10284 6724
rect 10968 6672 11020 6724
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 14924 6783 14976 6792
rect 14924 6749 14928 6783
rect 14928 6749 14962 6783
rect 14962 6749 14976 6783
rect 14924 6740 14976 6749
rect 15476 6740 15528 6792
rect 17408 6808 17460 6860
rect 12900 6672 12952 6724
rect 848 6604 900 6656
rect 3056 6604 3108 6656
rect 6920 6604 6972 6656
rect 7288 6604 7340 6656
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 9956 6604 10008 6656
rect 11612 6604 11664 6656
rect 13360 6604 13412 6656
rect 14556 6604 14608 6656
rect 15108 6715 15160 6724
rect 15108 6681 15117 6715
rect 15117 6681 15151 6715
rect 15151 6681 15160 6715
rect 15108 6672 15160 6681
rect 15752 6672 15804 6724
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 16396 6740 16448 6792
rect 16948 6740 17000 6792
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 16396 6604 16448 6656
rect 17592 6604 17644 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2320 6400 2372 6452
rect 2412 6400 2464 6452
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 3056 6400 3108 6452
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 2780 6332 2832 6384
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 4068 6375 4120 6384
rect 4068 6341 4077 6375
rect 4077 6341 4111 6375
rect 4111 6341 4120 6375
rect 4068 6332 4120 6341
rect 5724 6264 5776 6316
rect 6552 6400 6604 6452
rect 6920 6400 6972 6452
rect 8116 6332 8168 6384
rect 8484 6332 8536 6384
rect 8760 6400 8812 6452
rect 9128 6400 9180 6452
rect 9588 6400 9640 6452
rect 8944 6332 8996 6384
rect 10140 6332 10192 6384
rect 11428 6332 11480 6384
rect 11520 6332 11572 6384
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 6920 6264 6972 6316
rect 7104 6264 7156 6316
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 9036 6264 9088 6316
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 1952 6060 2004 6112
rect 2964 6060 3016 6112
rect 5632 6128 5684 6180
rect 8944 6196 8996 6248
rect 9128 6196 9180 6248
rect 9496 6307 9548 6316
rect 9496 6273 9505 6307
rect 9505 6273 9539 6307
rect 9539 6273 9548 6307
rect 9496 6264 9548 6273
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 10784 6196 10836 6248
rect 11336 6264 11388 6316
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 12256 6264 12308 6316
rect 11612 6196 11664 6248
rect 7472 6128 7524 6180
rect 7840 6128 7892 6180
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 13728 6400 13780 6452
rect 15108 6400 15160 6452
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 14096 6332 14148 6384
rect 17040 6400 17092 6452
rect 16396 6332 16448 6384
rect 13452 6196 13504 6248
rect 13728 6239 13780 6248
rect 13728 6205 13737 6239
rect 13737 6205 13771 6239
rect 13771 6205 13780 6239
rect 13728 6196 13780 6205
rect 16212 6264 16264 6316
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 16856 6375 16908 6384
rect 16856 6341 16865 6375
rect 16865 6341 16899 6375
rect 16899 6341 16908 6375
rect 16856 6332 16908 6341
rect 17316 6307 17368 6316
rect 17316 6273 17325 6307
rect 17325 6273 17359 6307
rect 17359 6273 17368 6307
rect 17316 6264 17368 6273
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 17592 6307 17644 6316
rect 17592 6273 17601 6307
rect 17601 6273 17635 6307
rect 17635 6273 17644 6307
rect 17592 6264 17644 6273
rect 15752 6196 15804 6248
rect 16028 6239 16080 6248
rect 16028 6205 16037 6239
rect 16037 6205 16071 6239
rect 16071 6205 16080 6239
rect 16028 6196 16080 6205
rect 16856 6196 16908 6248
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 9036 6103 9088 6112
rect 9036 6069 9045 6103
rect 9045 6069 9079 6103
rect 9079 6069 9088 6103
rect 9036 6060 9088 6069
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 16212 6128 16264 6180
rect 10692 6060 10744 6112
rect 10876 6060 10928 6112
rect 13636 6060 13688 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2044 5856 2096 5908
rect 2504 5856 2556 5908
rect 3240 5856 3292 5908
rect 3332 5856 3384 5908
rect 4344 5856 4396 5908
rect 4620 5856 4672 5908
rect 3516 5788 3568 5840
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 1860 5652 1912 5704
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2688 5652 2740 5704
rect 2780 5695 2832 5704
rect 2780 5661 2789 5695
rect 2789 5661 2823 5695
rect 2823 5661 2832 5695
rect 2780 5652 2832 5661
rect 3884 5720 3936 5772
rect 4804 5788 4856 5840
rect 5632 5856 5684 5908
rect 8484 5856 8536 5908
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 8760 5856 8812 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 6920 5788 6972 5840
rect 9588 5856 9640 5908
rect 10508 5856 10560 5908
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 14464 5856 14516 5908
rect 15476 5856 15528 5908
rect 16028 5856 16080 5908
rect 17316 5856 17368 5908
rect 9128 5788 9180 5840
rect 9312 5788 9364 5840
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 3516 5695 3568 5704
rect 3516 5661 3525 5695
rect 3525 5661 3559 5695
rect 3559 5661 3568 5695
rect 3516 5652 3568 5661
rect 3700 5652 3752 5704
rect 4344 5652 4396 5704
rect 4804 5652 4856 5704
rect 5908 5720 5960 5772
rect 4620 5584 4672 5636
rect 5448 5652 5500 5704
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 7380 5720 7432 5772
rect 7840 5720 7892 5772
rect 8116 5720 8168 5772
rect 8576 5720 8628 5772
rect 9588 5720 9640 5772
rect 10324 5720 10376 5772
rect 10784 5720 10836 5772
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 15292 5788 15344 5840
rect 5356 5627 5408 5636
rect 5356 5593 5365 5627
rect 5365 5593 5399 5627
rect 5399 5593 5408 5627
rect 5356 5584 5408 5593
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 8852 5652 8904 5704
rect 6092 5584 6144 5636
rect 3700 5516 3752 5568
rect 6552 5516 6604 5568
rect 7840 5584 7892 5636
rect 9404 5584 9456 5636
rect 10968 5695 11020 5704
rect 10968 5661 10977 5695
rect 10977 5661 11011 5695
rect 11011 5661 11020 5695
rect 10968 5652 11020 5661
rect 11060 5584 11112 5636
rect 12624 5652 12676 5704
rect 14188 5720 14240 5772
rect 14556 5763 14608 5772
rect 14556 5729 14565 5763
rect 14565 5729 14599 5763
rect 14599 5729 14608 5763
rect 14556 5720 14608 5729
rect 13176 5652 13228 5704
rect 13360 5695 13412 5704
rect 13360 5661 13369 5695
rect 13369 5661 13403 5695
rect 13403 5661 13412 5695
rect 13360 5652 13412 5661
rect 9956 5516 10008 5568
rect 10232 5516 10284 5568
rect 10324 5516 10376 5568
rect 12072 5516 12124 5568
rect 12440 5516 12492 5568
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 16304 5720 16356 5772
rect 15108 5695 15160 5704
rect 15108 5661 15117 5695
rect 15117 5661 15151 5695
rect 15151 5661 15160 5695
rect 15108 5652 15160 5661
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16120 5652 16172 5704
rect 16764 5652 16816 5704
rect 16948 5652 17000 5704
rect 13636 5627 13688 5636
rect 13636 5593 13645 5627
rect 13645 5593 13679 5627
rect 13679 5593 13688 5627
rect 13636 5584 13688 5593
rect 13820 5584 13872 5636
rect 15568 5584 15620 5636
rect 16212 5627 16264 5636
rect 16212 5593 16221 5627
rect 16221 5593 16255 5627
rect 16255 5593 16264 5627
rect 16212 5584 16264 5593
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 17684 5584 17736 5636
rect 13728 5516 13780 5568
rect 15108 5516 15160 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 15936 5516 15988 5568
rect 17132 5516 17184 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2872 5312 2924 5364
rect 5816 5312 5868 5364
rect 6644 5312 6696 5364
rect 4988 5244 5040 5296
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 9496 5312 9548 5364
rect 9772 5312 9824 5364
rect 11336 5312 11388 5364
rect 3608 5176 3660 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 4896 5176 4948 5228
rect 5540 5176 5592 5228
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 4068 5108 4120 5160
rect 4344 5151 4396 5160
rect 4344 5117 4353 5151
rect 4353 5117 4387 5151
rect 4387 5117 4396 5151
rect 4344 5108 4396 5117
rect 4620 5108 4672 5160
rect 6092 5219 6144 5228
rect 6092 5185 6101 5219
rect 6101 5185 6135 5219
rect 6135 5185 6144 5219
rect 6092 5176 6144 5185
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 7104 5176 7156 5228
rect 7196 5219 7248 5228
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 7380 5219 7432 5228
rect 7380 5185 7387 5219
rect 7387 5185 7432 5219
rect 7380 5176 7432 5185
rect 5448 5040 5500 5092
rect 6000 5040 6052 5092
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 7656 5219 7708 5228
rect 7656 5185 7670 5219
rect 7670 5185 7704 5219
rect 7704 5185 7708 5219
rect 7656 5176 7708 5185
rect 8944 5244 8996 5296
rect 9128 5244 9180 5296
rect 10140 5244 10192 5296
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 8668 5176 8720 5228
rect 8852 5108 8904 5160
rect 10048 5176 10100 5228
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 11796 5244 11848 5296
rect 10876 5219 10928 5228
rect 10876 5185 10885 5219
rect 10885 5185 10919 5219
rect 10919 5185 10928 5219
rect 10876 5176 10928 5185
rect 12256 5244 12308 5296
rect 12440 5287 12492 5296
rect 12440 5253 12449 5287
rect 12449 5253 12483 5287
rect 12483 5253 12492 5287
rect 12440 5244 12492 5253
rect 12808 5355 12860 5364
rect 12808 5321 12817 5355
rect 12817 5321 12851 5355
rect 12851 5321 12860 5355
rect 12808 5312 12860 5321
rect 14280 5312 14332 5364
rect 14740 5312 14792 5364
rect 15568 5355 15620 5364
rect 15568 5321 15577 5355
rect 15577 5321 15611 5355
rect 15611 5321 15620 5355
rect 15568 5312 15620 5321
rect 11888 5151 11940 5160
rect 11888 5117 11897 5151
rect 11897 5117 11931 5151
rect 11931 5117 11940 5151
rect 11888 5108 11940 5117
rect 12624 5176 12676 5228
rect 13176 5176 13228 5228
rect 15200 5244 15252 5296
rect 17040 5244 17092 5296
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 13912 5219 13964 5228
rect 13912 5185 13921 5219
rect 13921 5185 13955 5219
rect 13955 5185 13964 5219
rect 13912 5176 13964 5185
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 14464 5219 14516 5228
rect 14464 5185 14473 5219
rect 14473 5185 14507 5219
rect 14507 5185 14516 5219
rect 14464 5176 14516 5185
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 15016 5176 15068 5228
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 15476 5176 15528 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 17224 5176 17276 5228
rect 14004 5108 14056 5160
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 7472 5040 7524 5092
rect 4712 4972 4764 5024
rect 9404 5040 9456 5092
rect 9864 5040 9916 5092
rect 10416 5040 10468 5092
rect 10508 5040 10560 5092
rect 13820 5040 13872 5092
rect 15844 5040 15896 5092
rect 7564 4972 7616 5024
rect 7932 4972 7984 5024
rect 8576 4972 8628 5024
rect 9312 4972 9364 5024
rect 9680 4972 9732 5024
rect 11336 4972 11388 5024
rect 12256 4972 12308 5024
rect 15292 4972 15344 5024
rect 16856 4972 16908 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2596 4768 2648 4820
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 4160 4768 4212 4820
rect 4620 4768 4672 4820
rect 5724 4768 5776 4820
rect 7104 4768 7156 4820
rect 7656 4768 7708 4820
rect 7748 4768 7800 4820
rect 8852 4768 8904 4820
rect 8944 4811 8996 4820
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 9772 4768 9824 4820
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 11060 4768 11112 4820
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 3884 4700 3936 4752
rect 6276 4700 6328 4752
rect 12532 4768 12584 4820
rect 14372 4768 14424 4820
rect 14464 4768 14516 4820
rect 15200 4768 15252 4820
rect 6184 4675 6236 4684
rect 6184 4641 6194 4675
rect 6194 4641 6228 4675
rect 6228 4641 6236 4675
rect 6184 4632 6236 4641
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 4160 4564 4212 4616
rect 4804 4607 4856 4616
rect 3608 4539 3660 4548
rect 3608 4505 3617 4539
rect 3617 4505 3651 4539
rect 3651 4505 3660 4539
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 5356 4564 5408 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 3608 4496 3660 4505
rect 4988 4496 5040 4548
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 6460 4564 6512 4616
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 7932 4564 7984 4616
rect 8024 4607 8076 4616
rect 8024 4573 8033 4607
rect 8033 4573 8067 4607
rect 8067 4573 8076 4607
rect 8024 4564 8076 4573
rect 8668 4632 8720 4684
rect 6184 4496 6236 4548
rect 6644 4496 6696 4548
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 9312 4564 9364 4616
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 11428 4632 11480 4684
rect 8760 4539 8812 4548
rect 8760 4505 8769 4539
rect 8769 4505 8803 4539
rect 8803 4505 8812 4539
rect 8760 4496 8812 4505
rect 10692 4564 10744 4616
rect 10600 4496 10652 4548
rect 6736 4428 6788 4480
rect 7012 4428 7064 4480
rect 7748 4428 7800 4480
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 9128 4428 9180 4480
rect 9772 4428 9824 4480
rect 10232 4471 10284 4480
rect 10232 4437 10241 4471
rect 10241 4437 10275 4471
rect 10275 4437 10284 4471
rect 10232 4428 10284 4437
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 11520 4564 11572 4573
rect 11888 4675 11940 4684
rect 11888 4641 11897 4675
rect 11897 4641 11931 4675
rect 11931 4641 11940 4675
rect 11888 4632 11940 4641
rect 12164 4675 12216 4684
rect 12164 4641 12173 4675
rect 12173 4641 12207 4675
rect 12207 4641 12216 4675
rect 12164 4632 12216 4641
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 12348 4700 12400 4752
rect 12440 4700 12492 4752
rect 15660 4768 15712 4820
rect 15476 4700 15528 4752
rect 17040 4700 17092 4752
rect 13912 4632 13964 4684
rect 13820 4564 13872 4616
rect 16856 4632 16908 4684
rect 12992 4496 13044 4548
rect 13452 4496 13504 4548
rect 15292 4564 15344 4616
rect 15476 4564 15528 4616
rect 15568 4607 15620 4616
rect 15568 4573 15577 4607
rect 15577 4573 15611 4607
rect 15611 4573 15620 4607
rect 15568 4564 15620 4573
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 16948 4607 17000 4616
rect 16948 4573 16957 4607
rect 16957 4573 16991 4607
rect 16991 4573 17000 4607
rect 16948 4564 17000 4573
rect 15752 4496 15804 4548
rect 12256 4428 12308 4480
rect 14464 4428 14516 4480
rect 14556 4428 14608 4480
rect 15200 4428 15252 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 3608 4088 3660 4097
rect 5356 4224 5408 4276
rect 6184 4267 6236 4276
rect 6184 4233 6193 4267
rect 6193 4233 6227 4267
rect 6227 4233 6236 4267
rect 6184 4224 6236 4233
rect 6276 4224 6328 4276
rect 10140 4224 10192 4276
rect 10232 4267 10284 4276
rect 10232 4233 10241 4267
rect 10241 4233 10275 4267
rect 10275 4233 10284 4267
rect 10232 4224 10284 4233
rect 11244 4224 11296 4276
rect 11796 4224 11848 4276
rect 12072 4224 12124 4276
rect 12532 4267 12584 4276
rect 12532 4233 12541 4267
rect 12541 4233 12575 4267
rect 12575 4233 12584 4267
rect 12532 4224 12584 4233
rect 13820 4224 13872 4276
rect 14556 4224 14608 4276
rect 15936 4224 15988 4276
rect 4620 4156 4672 4208
rect 6920 4156 6972 4208
rect 8392 4156 8444 4208
rect 8760 4156 8812 4208
rect 5356 4088 5408 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 7472 4088 7524 4140
rect 9220 4088 9272 4140
rect 10692 4156 10744 4208
rect 15200 4156 15252 4208
rect 6276 4020 6328 4072
rect 8300 4020 8352 4072
rect 8576 3952 8628 4004
rect 9496 4020 9548 4072
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 12992 4131 13044 4140
rect 9680 4063 9732 4072
rect 9680 4029 9689 4063
rect 9689 4029 9723 4063
rect 9723 4029 9732 4063
rect 9680 4020 9732 4029
rect 10324 4063 10376 4072
rect 10324 4029 10333 4063
rect 10333 4029 10367 4063
rect 10367 4029 10376 4063
rect 10324 4020 10376 4029
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 13084 4088 13136 4140
rect 13912 4088 13964 4140
rect 14464 4088 14516 4140
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 16396 4131 16448 4140
rect 16396 4097 16405 4131
rect 16405 4097 16439 4131
rect 16439 4097 16448 4131
rect 16396 4088 16448 4097
rect 12900 3952 12952 4004
rect 14280 4020 14332 4072
rect 15568 4020 15620 4072
rect 16948 4088 17000 4140
rect 15384 3952 15436 4004
rect 9772 3884 9824 3936
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 16764 3884 16816 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 7012 3680 7064 3732
rect 6828 3612 6880 3664
rect 8024 3544 8076 3596
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 9036 2388 9088 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 9036 2252 9088 2304
rect 11612 2252 11664 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 7746 20956 7802 21756
rect 9678 20956 9734 21756
rect 11610 20956 11666 21756
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 7760 18970 7788 20956
rect 9692 18970 9720 20956
rect 11624 18970 11652 20956
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 16425 1532 17478
rect 1688 16794 1716 17614
rect 1964 17202 1992 18362
rect 5170 18320 5226 18329
rect 2320 18284 2372 18290
rect 7300 18290 7328 18634
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 5170 18255 5226 18264
rect 7104 18284 7156 18290
rect 2320 18226 2372 18232
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1872 16590 1900 16934
rect 1860 16584 1912 16590
rect 1860 16526 1912 16532
rect 1490 16416 1546 16425
rect 1490 16351 1546 16360
rect 1872 16250 1900 16526
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1306 15736 1362 15745
rect 1306 15671 1308 15680
rect 1360 15671 1362 15680
rect 1308 15642 1360 15648
rect 1688 15502 1716 15846
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 848 14816 900 14822
rect 848 14758 900 14764
rect 860 14521 888 14758
rect 1596 14618 1624 14962
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 846 14512 902 14521
rect 846 14447 902 14456
rect 1780 14414 1808 16050
rect 1860 15972 1912 15978
rect 1860 15914 1912 15920
rect 1872 14414 1900 15914
rect 1964 15366 1992 17138
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2056 15978 2084 16934
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 2148 16046 2176 16390
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2044 15972 2096 15978
rect 2044 15914 2096 15920
rect 2240 15502 2268 18022
rect 2332 16590 2360 18226
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 2412 17808 2464 17814
rect 2412 17750 2464 17756
rect 2424 17066 2452 17750
rect 3620 17746 3648 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 5184 17678 5212 18255
rect 7104 18226 7156 18232
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7116 17882 7144 18226
rect 7852 17882 7880 18362
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 3884 17672 3936 17678
rect 5172 17672 5224 17678
rect 3884 17614 3936 17620
rect 4066 17640 4122 17649
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 3792 17604 3844 17610
rect 3792 17546 3844 17552
rect 2412 17060 2464 17066
rect 2412 17002 2464 17008
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2332 16114 2360 16526
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2424 15722 2452 17002
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2516 16250 2544 16594
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2424 15694 2544 15722
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 1952 14544 2004 14550
rect 1952 14486 2004 14492
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1676 13728 1728 13734
rect 1306 13696 1362 13705
rect 1676 13670 1728 13676
rect 1306 13631 1362 13640
rect 1320 13530 1348 13631
rect 1308 13524 1360 13530
rect 1308 13466 1360 13472
rect 1688 13326 1716 13670
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1780 11694 1808 14350
rect 1872 13870 1900 14350
rect 1964 14074 1992 14486
rect 2148 14346 2176 15302
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2056 13954 2084 14214
rect 2148 14006 2176 14282
rect 1964 13926 2084 13954
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1964 12442 1992 13926
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1768 11688 1820 11694
rect 1122 11656 1178 11665
rect 1768 11630 1820 11636
rect 1122 11591 1178 11600
rect 1136 11354 1164 11591
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1124 11348 1176 11354
rect 1124 11290 1176 11296
rect 1688 11150 1716 11494
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9625 1532 9862
rect 1688 9722 1716 9998
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 1780 8906 1808 11630
rect 1872 11354 1900 11698
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 2056 10418 2084 13806
rect 2148 10810 2176 13942
rect 2240 13433 2268 15438
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2424 14414 2452 14894
rect 2516 14482 2544 15694
rect 2608 15008 2636 17546
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3252 17270 3280 17478
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2700 16590 2728 17070
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2688 15020 2740 15026
rect 2608 14980 2688 15008
rect 2688 14962 2740 14968
rect 2700 14929 2728 14962
rect 2686 14920 2742 14929
rect 2686 14855 2742 14864
rect 2686 14512 2742 14521
rect 2504 14476 2556 14482
rect 2686 14447 2742 14456
rect 2504 14418 2556 14424
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2332 13938 2360 14214
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2424 13530 2452 13942
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2226 13424 2282 13433
rect 2226 13359 2282 13368
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1872 10390 2084 10418
rect 1872 9738 1900 10390
rect 2134 10024 2190 10033
rect 2134 9959 2190 9968
rect 1872 9710 2084 9738
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1872 9178 1900 9522
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1872 8514 1900 9114
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1780 8486 1900 8514
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1688 8090 1716 8434
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1780 7886 1808 8486
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1780 7546 1808 7822
rect 1872 7585 1900 8298
rect 1964 7954 1992 9522
rect 2056 9178 2084 9710
rect 2148 9518 2176 9959
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2240 8974 2268 12378
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2332 9654 2360 11086
rect 2424 11082 2452 11834
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2516 10962 2544 14418
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2608 13870 2636 14214
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2700 12186 2728 14447
rect 2792 13258 2820 15438
rect 2884 15026 2912 16118
rect 3068 16114 3096 16934
rect 3344 16726 3372 17138
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3332 16720 3384 16726
rect 3332 16662 3384 16668
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 3160 15910 3188 16662
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 14482 2912 14758
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2976 14414 3004 15574
rect 3056 15496 3108 15502
rect 3054 15464 3056 15473
rect 3108 15464 3110 15473
rect 3054 15399 3110 15408
rect 3160 15348 3188 15846
rect 3252 15570 3280 16526
rect 3436 16182 3464 16730
rect 3528 16590 3556 16730
rect 3608 16720 3660 16726
rect 3608 16662 3660 16668
rect 3620 16590 3648 16662
rect 3712 16590 3740 17478
rect 3804 17202 3832 17546
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3896 16794 3924 17614
rect 5172 17614 5224 17620
rect 4066 17575 4122 17584
rect 4080 17542 4108 17575
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3068 15320 3188 15348
rect 3068 14414 3096 15320
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 12306 2820 13194
rect 2884 13025 2912 14282
rect 3160 14074 3188 14350
rect 3252 14113 3280 15506
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3344 14618 3372 15438
rect 3436 14822 3464 15438
rect 3620 15434 3648 16526
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3238 14104 3294 14113
rect 3148 14068 3200 14074
rect 3238 14039 3294 14048
rect 3148 14010 3200 14016
rect 2964 14000 3016 14006
rect 2964 13942 3016 13948
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 2870 13016 2926 13025
rect 2870 12951 2926 12960
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2884 12434 2912 12854
rect 2976 12714 3004 13942
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3160 13326 3188 13466
rect 3252 13326 3280 13942
rect 3344 13938 3372 14554
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3146 12880 3202 12889
rect 3146 12815 3148 12824
rect 3200 12815 3202 12824
rect 3332 12844 3384 12850
rect 3148 12786 3200 12792
rect 3332 12786 3384 12792
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 2884 12406 3004 12434
rect 2870 12336 2926 12345
rect 2780 12300 2832 12306
rect 2870 12271 2926 12280
rect 2780 12242 2832 12248
rect 2608 11150 2636 12174
rect 2700 12158 2820 12186
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2700 11830 2728 12038
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2792 11762 2820 12158
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2884 11626 2912 12271
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2700 10962 2728 11018
rect 2884 11014 2912 11562
rect 2516 10934 2728 10962
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2424 9586 2452 10746
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2608 9489 2636 9522
rect 2594 9480 2650 9489
rect 2594 9415 2650 9424
rect 2318 9072 2374 9081
rect 2318 9007 2374 9016
rect 2332 8974 2360 9007
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1858 7576 1914 7585
rect 1768 7540 1820 7546
rect 1858 7511 1914 7520
rect 1768 7482 1820 7488
rect 1964 7410 1992 7890
rect 1952 7404 2004 7410
rect 1872 7364 1952 7392
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6798 1716 7142
rect 1676 6792 1728 6798
rect 846 6760 902 6769
rect 1676 6734 1728 6740
rect 846 6695 902 6704
rect 860 6662 888 6695
rect 848 6656 900 6662
rect 848 6598 900 6604
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5710 1716 6054
rect 1872 5710 1900 7364
rect 1952 7346 2004 7352
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5710 1992 6054
rect 2056 5914 2084 8434
rect 2332 6458 2360 8774
rect 2424 6458 2452 8910
rect 2608 7410 2636 9415
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2516 6798 2544 7142
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2332 6322 2360 6394
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2516 5914 2544 6258
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2608 4826 2636 7346
rect 2700 5710 2728 10934
rect 2884 10062 2912 10950
rect 2976 10266 3004 12406
rect 3160 11762 3188 12582
rect 3344 12442 3372 12786
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 3160 11354 3188 11698
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3252 11234 3280 12310
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 11830 3372 12174
rect 3436 12102 3464 14758
rect 3620 14482 3648 14758
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3528 13258 3556 13874
rect 3608 13864 3660 13870
rect 3712 13852 3740 15914
rect 3896 15706 3924 16458
rect 4080 16046 4108 17478
rect 4816 17202 4844 17478
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4172 16250 4200 16458
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 16040 4120 16046
rect 3988 16000 4068 16028
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3660 13824 3740 13852
rect 3608 13806 3660 13812
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3620 12850 3648 13806
rect 3804 13512 3832 14418
rect 3896 14346 3924 15506
rect 3988 14550 4016 16000
rect 4068 15982 4120 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 3976 14544 4028 14550
rect 3974 14512 3976 14521
rect 4028 14512 4030 14521
rect 3974 14447 4030 14456
rect 4080 14414 4108 15098
rect 4172 14958 4200 15438
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4448 14414 4476 14486
rect 4068 14408 4120 14414
rect 3974 14376 4030 14385
rect 3884 14340 3936 14346
rect 4068 14350 4120 14356
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 3974 14311 4030 14320
rect 3884 14282 3936 14288
rect 3882 13968 3938 13977
rect 3882 13903 3884 13912
rect 3936 13903 3938 13912
rect 3884 13874 3936 13880
rect 3712 13484 3832 13512
rect 3712 13258 3740 13484
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3804 13002 3832 13330
rect 3712 12974 3832 13002
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3332 11824 3384 11830
rect 3332 11766 3384 11772
rect 3160 11206 3280 11234
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2976 9586 3004 10202
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2792 7392 2820 9522
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2884 8974 2912 9318
rect 2976 9042 3004 9318
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2872 7404 2924 7410
rect 2792 7364 2872 7392
rect 2872 7346 2924 7352
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2792 5710 2820 6326
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2884 5370 2912 7346
rect 2976 6322 3004 8978
rect 3068 7410 3096 9862
rect 3160 9586 3188 11206
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 6866 3188 7346
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6458 3096 6598
rect 3056 6452 3108 6458
rect 3252 6440 3280 11018
rect 3436 9178 3464 12038
rect 3712 10810 3740 12974
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 12209 3832 12786
rect 3896 12345 3924 13874
rect 3988 13394 4016 14311
rect 4080 13938 4108 14350
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 13938 4568 14214
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3882 12336 3938 12345
rect 3882 12271 3938 12280
rect 3790 12200 3846 12209
rect 3790 12135 3846 12144
rect 3884 12164 3936 12170
rect 3804 11286 3832 12135
rect 3884 12106 3936 12112
rect 3896 11354 3924 12106
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3698 10704 3754 10713
rect 3804 10674 3832 11086
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3698 10639 3700 10648
rect 3752 10639 3754 10648
rect 3792 10668 3844 10674
rect 3700 10610 3752 10616
rect 3792 10610 3844 10616
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3608 9648 3660 9654
rect 3606 9616 3608 9625
rect 3660 9616 3662 9625
rect 3606 9551 3662 9560
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 7857 3464 8910
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3422 7848 3478 7857
rect 3422 7783 3478 7792
rect 3436 7546 3464 7783
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3344 7002 3372 7346
rect 3528 7342 3556 8230
rect 3620 7818 3648 8774
rect 3712 8090 3740 9522
rect 3804 8974 3832 9998
rect 3896 9178 3924 10950
rect 3988 10674 4016 13194
rect 4080 12646 4108 13874
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 12986 4660 17138
rect 4816 16726 4844 17138
rect 5354 17096 5410 17105
rect 5354 17031 5410 17040
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 5092 16590 5120 16934
rect 5080 16584 5132 16590
rect 4894 16552 4950 16561
rect 5080 16526 5132 16532
rect 4894 16487 4896 16496
rect 4948 16487 4950 16496
rect 4896 16458 4948 16464
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5368 16182 5396 17031
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 5080 16108 5132 16114
rect 5080 16050 5132 16056
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 4710 15736 4766 15745
rect 4710 15671 4712 15680
rect 4764 15671 4766 15680
rect 4712 15642 4764 15648
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4724 15094 4752 15370
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4724 14618 4752 15030
rect 4816 14958 4844 16050
rect 5092 15570 5120 16050
rect 5276 15910 5304 16050
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5460 15722 5488 16934
rect 5736 16794 5764 17138
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5276 15694 5488 15722
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 5184 15366 5212 15642
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 5184 14793 5212 15098
rect 5276 15026 5304 15694
rect 5552 15609 5580 16050
rect 5644 16017 5672 16526
rect 5736 16425 5764 16730
rect 5722 16416 5778 16425
rect 5722 16351 5778 16360
rect 5828 16266 5856 17274
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6196 16590 6224 16934
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 5736 16238 5856 16266
rect 5630 16008 5686 16017
rect 5736 15978 5764 16238
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 5630 15943 5686 15952
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5538 15600 5594 15609
rect 5538 15535 5594 15544
rect 5644 15502 5672 15642
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5368 15162 5396 15438
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5170 14784 5226 14793
rect 5170 14719 5226 14728
rect 5276 14657 5304 14962
rect 5368 14890 5396 15098
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5262 14648 5318 14657
rect 4712 14612 4764 14618
rect 5262 14583 5318 14592
rect 4712 14554 4764 14560
rect 4724 14006 4752 14554
rect 5368 14550 5396 14826
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 4816 14414 4844 14486
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 5644 14346 5672 15438
rect 5736 14890 5764 15914
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4712 14000 4764 14006
rect 4712 13942 4764 13948
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4724 13462 4752 13806
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4816 13394 4844 13738
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12918 4752 13194
rect 5092 13190 5120 13874
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4344 12368 4396 12374
rect 4250 12336 4306 12345
rect 4068 12300 4120 12306
rect 4344 12310 4396 12316
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 4250 12271 4306 12280
rect 4068 12242 4120 12248
rect 4080 10810 4108 12242
rect 4264 12238 4292 12271
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4158 11792 4214 11801
rect 4158 11727 4160 11736
rect 4212 11727 4214 11736
rect 4160 11698 4212 11704
rect 4264 11665 4292 12174
rect 4356 11830 4384 12310
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4448 11762 4476 12310
rect 4632 12238 4660 12582
rect 4724 12374 4752 12854
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4540 12073 4568 12106
rect 5000 12084 5028 12310
rect 5092 12238 5120 12718
rect 5184 12646 5212 12922
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4526 12064 4582 12073
rect 4526 11999 4582 12008
rect 4816 12056 5028 12084
rect 5092 12084 5120 12174
rect 5184 12152 5212 12582
rect 5276 12442 5304 14214
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5184 12124 5396 12152
rect 5092 12056 5304 12084
rect 4816 11778 4844 12056
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4620 11756 4672 11762
rect 4816 11750 4936 11778
rect 4620 11698 4672 11704
rect 4250 11656 4306 11665
rect 4250 11591 4306 11600
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11354 4660 11698
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4724 11200 4752 11494
rect 4540 11172 4752 11200
rect 4436 11144 4488 11150
rect 4540 11132 4568 11172
rect 4488 11104 4568 11132
rect 4436 11086 4488 11092
rect 4816 11064 4844 11630
rect 4632 11036 4844 11064
rect 4632 10810 4660 11036
rect 4908 10996 4936 11750
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5184 11665 5212 11698
rect 5170 11656 5226 11665
rect 5170 11591 5226 11600
rect 4986 11112 5042 11121
rect 4986 11047 4988 11056
rect 5040 11047 5042 11056
rect 4988 11018 5040 11024
rect 5184 11014 5212 11591
rect 4724 10968 4936 10996
rect 5172 11008 5224 11014
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3988 10577 4016 10610
rect 3974 10568 4030 10577
rect 3974 10503 4030 10512
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 3988 10062 4016 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4342 10160 4398 10169
rect 4632 10130 4660 10406
rect 4342 10095 4398 10104
rect 4620 10124 4672 10130
rect 4356 10062 4384 10095
rect 4620 10066 4672 10072
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4080 9654 4108 9998
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3884 9172 3936 9178
rect 4080 9160 4108 9590
rect 4356 9450 4384 9998
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4620 9172 4672 9178
rect 4080 9132 4200 9160
rect 3884 9114 3936 9120
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3252 6412 3372 6440
rect 3056 6394 3108 6400
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 2976 6118 3004 6258
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 3252 5914 3280 6258
rect 3344 5914 3372 6412
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3344 5710 3372 5850
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3528 5710 3556 5782
rect 3712 5710 3740 8026
rect 3804 7546 3832 8910
rect 3896 8838 3924 9114
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3896 7886 3924 8463
rect 4080 8430 4108 8978
rect 4172 8634 4200 9132
rect 4620 9114 4672 9120
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4252 8968 4304 8974
rect 4344 8968 4396 8974
rect 4252 8910 4304 8916
rect 4342 8936 4344 8945
rect 4396 8936 4398 8945
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4264 8498 4292 8910
rect 4342 8871 4398 8880
rect 4356 8498 4384 8871
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4068 8424 4120 8430
rect 3988 8372 4068 8378
rect 3988 8366 4120 8372
rect 3988 8350 4108 8366
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3804 6798 3832 7482
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3896 6118 3924 7142
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3712 5574 3740 5646
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3344 4729 3372 4762
rect 3330 4720 3386 4729
rect 3330 4655 3386 4664
rect 3620 4554 3648 5170
rect 3712 5166 3740 5510
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3896 4758 3924 5714
rect 3988 5234 4016 8350
rect 4356 8294 4384 8434
rect 4080 8266 4384 8294
rect 4540 8276 4568 8978
rect 4632 8537 4660 9114
rect 4724 8906 4752 10968
rect 5172 10950 5224 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 4816 10169 4844 10678
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 10305 5028 10474
rect 4986 10296 5042 10305
rect 4986 10231 5042 10240
rect 5000 10198 5028 10231
rect 4988 10192 5040 10198
rect 4802 10160 4858 10169
rect 4988 10134 5040 10140
rect 4802 10095 4858 10104
rect 5092 10062 5120 10542
rect 5184 10130 5212 10678
rect 5276 10674 5304 12056
rect 5368 11676 5396 12124
rect 5460 11801 5488 13330
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5446 11792 5502 11801
rect 5446 11727 5502 11736
rect 5368 11648 5488 11676
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5368 11354 5396 11494
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5368 10418 5396 11290
rect 5276 10390 5396 10418
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4988 9580 5040 9586
rect 4816 9540 4988 9568
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4816 8616 4844 9540
rect 4988 9522 5040 9528
rect 5092 9330 5120 9658
rect 5276 9518 5304 10390
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5172 9376 5224 9382
rect 4908 9302 5120 9330
rect 5170 9344 5172 9353
rect 5224 9344 5226 9353
rect 4908 9042 4936 9302
rect 5170 9279 5226 9288
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 5000 8974 5028 9114
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5172 8968 5224 8974
rect 5276 8956 5304 9454
rect 5368 9178 5396 10066
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5224 8928 5304 8956
rect 5172 8910 5224 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4988 8628 5040 8634
rect 4816 8588 4936 8616
rect 4618 8528 4674 8537
rect 4724 8498 4839 8514
rect 4618 8463 4674 8472
rect 4712 8492 4839 8498
rect 4764 8486 4839 8492
rect 4712 8434 4764 8440
rect 4811 8412 4839 8486
rect 4811 8384 4844 8412
rect 4712 8356 4764 8362
rect 4618 8290 4674 8299
rect 4712 8298 4764 8304
rect 4080 7528 4108 8266
rect 4540 8248 4618 8276
rect 4618 8225 4674 8234
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4342 7984 4398 7993
rect 4724 7954 4752 8298
rect 4816 7954 4844 8384
rect 4908 8265 4936 8588
rect 5276 8616 5304 8928
rect 4988 8570 5040 8576
rect 5092 8588 5304 8616
rect 5000 8294 5028 8570
rect 4988 8288 5040 8294
rect 4894 8256 4950 8265
rect 4988 8230 5040 8236
rect 4894 8191 4950 8200
rect 4342 7919 4398 7928
rect 4712 7948 4764 7954
rect 4356 7886 4384 7919
rect 4712 7890 4764 7896
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4908 7886 4936 8191
rect 4986 8120 5042 8129
rect 4986 8055 4988 8064
rect 5040 8055 5042 8064
rect 4988 8026 5040 8032
rect 5092 7886 5120 8588
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5172 8424 5224 8430
rect 5276 8401 5304 8434
rect 5172 8366 5224 8372
rect 5262 8392 5318 8401
rect 5184 7886 5212 8366
rect 5262 8327 5318 8336
rect 5368 7886 5396 9114
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5184 7750 5212 7822
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 5172 7744 5224 7750
rect 5460 7732 5488 11648
rect 5552 10849 5580 12242
rect 5538 10840 5594 10849
rect 5538 10775 5594 10784
rect 5552 10470 5580 10775
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 9722 5580 10406
rect 5644 9926 5672 13806
rect 5736 12238 5764 13806
rect 5828 13734 5856 16050
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 6012 15366 6040 15914
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6104 15638 6132 15846
rect 6092 15632 6144 15638
rect 6092 15574 6144 15580
rect 6196 15570 6224 16050
rect 6288 16046 6316 17138
rect 6748 17134 6776 17750
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 6736 17128 6788 17134
rect 7116 17105 7144 17138
rect 6736 17070 6788 17076
rect 7102 17096 7158 17105
rect 6748 16590 6776 17070
rect 7208 17066 7236 17546
rect 7300 17513 7328 17614
rect 7286 17504 7342 17513
rect 7286 17439 7342 17448
rect 7576 17241 7604 17614
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7668 17338 7696 17478
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7562 17232 7618 17241
rect 7380 17196 7432 17202
rect 7562 17167 7618 17176
rect 7380 17138 7432 17144
rect 7102 17031 7158 17040
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7024 16726 7052 16934
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6288 15570 6316 15982
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6000 15360 6052 15366
rect 5920 15320 6000 15348
rect 5920 13818 5948 15320
rect 6000 15302 6052 15308
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6012 14414 6040 15098
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6012 13938 6040 14350
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6104 13977 6132 14214
rect 6182 14104 6238 14113
rect 6288 14074 6316 15506
rect 6380 15434 6408 16526
rect 6460 16516 6512 16522
rect 6460 16458 6512 16464
rect 6472 15910 6500 16458
rect 6748 16232 6776 16526
rect 6656 16204 6776 16232
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6656 15722 6684 16204
rect 6920 16108 6972 16114
rect 7024 16096 7052 16526
rect 6972 16068 7052 16096
rect 6920 16050 6972 16056
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6472 15694 6684 15722
rect 6840 15706 6868 15914
rect 6828 15700 6880 15706
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6472 14278 6500 15694
rect 6828 15642 6880 15648
rect 6552 15632 6604 15638
rect 6550 15600 6552 15609
rect 6604 15600 6606 15609
rect 6550 15535 6606 15544
rect 6734 15600 6790 15609
rect 6734 15535 6790 15544
rect 6748 15502 6776 15535
rect 6736 15496 6788 15502
rect 6656 15456 6736 15484
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6182 14039 6238 14048
rect 6276 14068 6328 14074
rect 6090 13968 6146 13977
rect 6000 13932 6052 13938
rect 6196 13938 6224 14039
rect 6276 14010 6328 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6090 13903 6146 13912
rect 6184 13932 6236 13938
rect 6000 13874 6052 13880
rect 6184 13874 6236 13880
rect 6092 13864 6144 13870
rect 5920 13790 6040 13818
rect 6092 13806 6144 13812
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5828 12918 5856 13670
rect 6012 13530 6040 13790
rect 6104 13705 6132 13806
rect 6090 13696 6146 13705
rect 6090 13631 6146 13640
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5828 11744 5856 12854
rect 5920 11898 5948 13126
rect 6012 12850 6040 13466
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 6012 12434 6040 12786
rect 6104 12646 6132 13262
rect 6092 12640 6144 12646
rect 6090 12608 6092 12617
rect 6144 12608 6146 12617
rect 6090 12543 6146 12552
rect 6012 12406 6132 12434
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 6012 11762 6040 12174
rect 5736 11716 5856 11744
rect 5908 11756 5960 11762
rect 5736 10674 5764 11716
rect 5908 11698 5960 11704
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5828 10810 5856 11562
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5814 10432 5870 10441
rect 5814 10367 5870 10376
rect 5724 10124 5776 10130
rect 5828 10112 5856 10367
rect 5776 10084 5856 10112
rect 5724 10066 5776 10072
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5736 9722 5764 9930
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 8634 5580 9522
rect 5644 8974 5672 9590
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5736 9178 5764 9318
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5736 8673 5764 8774
rect 5722 8664 5778 8673
rect 5540 8628 5592 8634
rect 5722 8599 5778 8608
rect 5540 8570 5592 8576
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5552 7886 5580 8230
rect 5630 7984 5686 7993
rect 5630 7919 5686 7928
rect 5644 7886 5672 7919
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5172 7686 5224 7692
rect 5276 7704 5488 7732
rect 5552 7721 5580 7822
rect 5538 7712 5594 7721
rect 4436 7540 4488 7546
rect 4080 7500 4200 7528
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4080 7313 4108 7346
rect 4066 7304 4122 7313
rect 4066 7239 4122 7248
rect 4172 7188 4200 7500
rect 4436 7482 4488 7488
rect 4448 7410 4476 7482
rect 4724 7449 4752 7686
rect 4710 7440 4766 7449
rect 4436 7404 4488 7410
rect 4710 7375 4766 7384
rect 4436 7346 4488 7352
rect 4816 7290 4844 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5078 7440 5134 7449
rect 5078 7375 5080 7384
rect 5132 7375 5134 7384
rect 5172 7404 5224 7410
rect 5080 7346 5132 7352
rect 5172 7346 5224 7352
rect 5184 7313 5212 7346
rect 5276 7342 5304 7704
rect 5538 7647 5594 7656
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5264 7336 5316 7342
rect 5170 7304 5226 7313
rect 4816 7262 5028 7290
rect 4080 7160 4200 7188
rect 4804 7200 4856 7206
rect 4080 6780 4108 7160
rect 4804 7142 4856 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4160 6792 4212 6798
rect 4080 6752 4160 6780
rect 4344 6792 4396 6798
rect 4160 6734 4212 6740
rect 4342 6760 4344 6769
rect 4396 6760 4398 6769
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 4080 6390 4108 6423
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4172 6100 4200 6734
rect 4342 6695 4398 6704
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4448 6168 4476 6666
rect 4540 6236 4568 6802
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4724 6361 4752 6666
rect 4710 6352 4766 6361
rect 4710 6287 4766 6296
rect 4540 6225 4752 6236
rect 4540 6216 4766 6225
rect 4540 6208 4710 6216
rect 4448 6140 4660 6168
rect 4710 6151 4766 6160
rect 4080 6072 4200 6100
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4080 5166 4108 6072
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5914 4660 6140
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4356 5710 4384 5850
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4356 5166 4384 5646
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4632 5166 4660 5578
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4344 5160 4396 5166
rect 4344 5102 4396 5108
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4826 4660 5102
rect 4724 5030 4752 6151
rect 4816 5846 4844 7142
rect 5000 6798 5028 7262
rect 5264 7278 5316 7284
rect 5170 7239 5226 7248
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5184 6644 5212 7239
rect 5262 6896 5318 6905
rect 5262 6831 5318 6840
rect 5276 6798 5304 6831
rect 5264 6792 5316 6798
rect 5316 6752 5396 6780
rect 5264 6734 5316 6740
rect 5184 6616 5304 6644
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5276 6361 5304 6616
rect 5262 6352 5318 6361
rect 5262 6287 5318 6296
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 4172 4622 4200 4762
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 3620 4146 3648 4490
rect 4632 4214 4660 4762
rect 4816 4622 4844 5646
rect 5368 5642 5396 6752
rect 5460 5710 5488 7482
rect 5552 7206 5580 7647
rect 5736 7410 5764 8599
rect 5828 7970 5856 10084
rect 5920 9382 5948 11698
rect 5998 11656 6054 11665
rect 5998 11591 6054 11600
rect 5908 9376 5960 9382
rect 5906 9344 5908 9353
rect 5960 9344 5962 9353
rect 5906 9279 5962 9288
rect 6012 9194 6040 11591
rect 6104 10674 6132 12406
rect 6196 12288 6224 13874
rect 6288 13462 6316 14010
rect 6380 13841 6408 14010
rect 6366 13832 6422 13841
rect 6366 13767 6422 13776
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6380 13326 6408 13670
rect 6472 13394 6500 14214
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6196 12260 6316 12288
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6196 11626 6224 12106
rect 6288 11898 6316 12260
rect 6472 12238 6500 12922
rect 6564 12617 6592 14826
rect 6550 12608 6606 12617
rect 6550 12543 6606 12552
rect 6550 12472 6606 12481
rect 6550 12407 6606 12416
rect 6460 12232 6512 12238
rect 6366 12200 6422 12209
rect 6460 12174 6512 12180
rect 6366 12135 6422 12144
rect 6380 12102 6408 12135
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6366 11928 6422 11937
rect 6276 11892 6328 11898
rect 6366 11863 6422 11872
rect 6460 11892 6512 11898
rect 6276 11834 6328 11840
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6288 11506 6316 11698
rect 6196 11478 6316 11506
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 6196 10577 6224 11478
rect 6274 11384 6330 11393
rect 6274 11319 6330 11328
rect 6288 11150 6316 11319
rect 6380 11257 6408 11863
rect 6460 11834 6512 11840
rect 6366 11248 6422 11257
rect 6366 11183 6422 11192
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6380 10606 6408 10950
rect 6368 10600 6420 10606
rect 6182 10568 6238 10577
rect 6368 10542 6420 10548
rect 6182 10503 6238 10512
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 10062 6408 10406
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6368 9580 6420 9586
rect 6472 9568 6500 11834
rect 6564 11694 6592 12407
rect 6656 11762 6684 15456
rect 6736 15438 6788 15444
rect 6840 15162 6868 15642
rect 6932 15570 6960 16050
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6920 15360 6972 15366
rect 7024 15348 7052 15914
rect 7116 15434 7144 16730
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7208 15745 7236 16390
rect 7300 16289 7328 16934
rect 7392 16794 7420 17138
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7286 16280 7342 16289
rect 7286 16215 7342 16224
rect 7194 15736 7250 15745
rect 7194 15671 7250 15680
rect 7104 15428 7156 15434
rect 7104 15370 7156 15376
rect 6972 15320 7052 15348
rect 6920 15302 6972 15308
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 7024 15026 7052 15320
rect 7208 15314 7236 15671
rect 7116 15286 7236 15314
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6748 14278 6776 14758
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 14006 6776 14214
rect 6840 14074 6868 14894
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6932 13920 6960 14894
rect 7024 14482 7052 14962
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7012 13932 7064 13938
rect 6932 13892 7012 13920
rect 7012 13874 7064 13880
rect 6920 13796 6972 13802
rect 7116 13784 7144 15286
rect 7300 15026 7328 16215
rect 7484 16153 7512 17070
rect 7576 16998 7604 17070
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 16590 7604 16934
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7654 16552 7710 16561
rect 7654 16487 7710 16496
rect 7470 16144 7526 16153
rect 7470 16079 7526 16088
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14482 7236 14758
rect 7300 14618 7328 14962
rect 7392 14890 7420 15642
rect 7668 15502 7696 16487
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7484 14618 7512 15438
rect 7576 15162 7604 15438
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7760 14958 7788 17546
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7852 15638 7880 16458
rect 7944 15706 7972 18770
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 8036 18426 8064 18702
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 8956 18290 8984 18838
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9416 18426 9444 18702
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9600 18329 9628 18634
rect 10336 18426 10364 18770
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 9586 18320 9642 18329
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8944 18284 8996 18290
rect 9586 18255 9642 18264
rect 10140 18284 10192 18290
rect 8944 18226 8996 18232
rect 8036 17610 8064 18226
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8312 17814 8340 18158
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8116 17672 8168 17678
rect 8168 17632 8248 17660
rect 8116 17614 8168 17620
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 8220 17218 8248 17632
rect 8312 17338 8340 17750
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8404 17218 8432 18158
rect 8484 17672 8536 17678
rect 8588 17660 8616 18158
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8536 17632 8616 17660
rect 8668 17672 8720 17678
rect 8484 17614 8536 17620
rect 8668 17614 8720 17620
rect 8220 17190 8432 17218
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7840 15632 7892 15638
rect 7892 15580 7972 15586
rect 7840 15574 7972 15580
rect 7852 15558 7972 15574
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 6920 13738 6972 13744
rect 7024 13756 7144 13784
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12102 6776 13262
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6564 10742 6592 11630
rect 6734 11112 6790 11121
rect 6734 11047 6790 11056
rect 6552 10736 6604 10742
rect 6604 10696 6684 10724
rect 6552 10678 6604 10684
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6420 9540 6500 9568
rect 6368 9522 6420 9528
rect 6092 9444 6144 9450
rect 6564 9432 6592 9930
rect 6656 9761 6684 10696
rect 6748 10033 6776 11047
rect 6734 10024 6790 10033
rect 6734 9959 6790 9968
rect 6734 9888 6790 9897
rect 6734 9823 6790 9832
rect 6642 9752 6698 9761
rect 6642 9687 6698 9696
rect 6656 9552 6684 9687
rect 6748 9654 6776 9823
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6644 9546 6696 9552
rect 6644 9488 6696 9494
rect 6736 9546 6788 9552
rect 6736 9488 6788 9494
rect 6748 9432 6776 9488
rect 6564 9404 6776 9432
rect 6092 9386 6144 9392
rect 5920 9166 6040 9194
rect 5920 8294 5948 9166
rect 6104 9024 6132 9386
rect 6550 9208 6606 9217
rect 6748 9194 6776 9404
rect 6550 9143 6606 9152
rect 6656 9166 6776 9194
rect 6104 8996 6500 9024
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6012 8838 6040 8910
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6090 8800 6146 8809
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5828 7942 5948 7970
rect 5817 7880 5869 7886
rect 5817 7822 5869 7828
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5644 7041 5672 7346
rect 5630 7032 5686 7041
rect 5540 6996 5592 7002
rect 5630 6967 5686 6976
rect 5540 6938 5592 6944
rect 5552 6798 5580 6938
rect 5736 6866 5764 7346
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5446 5400 5502 5409
rect 5446 5335 5502 5344
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 4622 4936 5170
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5000 4554 5028 5238
rect 5460 5098 5488 5335
rect 5552 5234 5580 6734
rect 5644 6186 5672 6734
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5644 5914 5672 6122
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5460 4622 5488 5034
rect 5736 4826 5764 6258
rect 5828 5794 5856 7822
rect 5920 7426 5948 7942
rect 6012 7546 6040 8774
rect 6090 8735 6146 8744
rect 6104 8294 6132 8735
rect 6196 8537 6224 8842
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6182 8528 6238 8537
rect 6380 8498 6408 8774
rect 6182 8463 6238 8472
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6104 8266 6224 8294
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6104 7478 6132 7890
rect 6092 7472 6144 7478
rect 5920 7398 6040 7426
rect 6092 7414 6144 7420
rect 6012 6882 6040 7398
rect 6196 7002 6224 8266
rect 6274 7984 6330 7993
rect 6274 7919 6276 7928
rect 6328 7919 6330 7928
rect 6276 7890 6328 7896
rect 6288 7732 6316 7890
rect 6380 7857 6408 8298
rect 6472 7886 6500 8996
rect 6460 7880 6512 7886
rect 6366 7848 6422 7857
rect 6460 7822 6512 7828
rect 6366 7783 6422 7792
rect 6288 7704 6408 7732
rect 6274 7576 6330 7585
rect 6274 7511 6330 7520
rect 6288 7410 6316 7511
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6012 6854 6132 6882
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5906 6488 5962 6497
rect 6012 6458 6040 6734
rect 5906 6423 5908 6432
rect 5960 6423 5962 6432
rect 6000 6452 6052 6458
rect 5908 6394 5960 6400
rect 6000 6394 6052 6400
rect 6104 6338 6132 6854
rect 6012 6310 6132 6338
rect 5828 5778 5948 5794
rect 5828 5772 5960 5778
rect 5828 5766 5908 5772
rect 5908 5714 5960 5720
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5828 5370 5856 5646
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 6012 5098 6040 6310
rect 6288 6100 6316 7346
rect 6380 6225 6408 7704
rect 6472 7274 6500 7822
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6564 6458 6592 9143
rect 6656 8945 6684 9166
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6642 8936 6698 8945
rect 6642 8871 6698 8880
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6366 6216 6422 6225
rect 6366 6151 6422 6160
rect 6288 6072 6408 6100
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6104 5234 6132 5578
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5368 4282 5396 4558
rect 6196 4554 6224 4626
rect 6288 4622 6316 4694
rect 6380 4690 6408 6072
rect 6564 5574 6592 6394
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6656 5370 6684 8230
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6458 4720 6514 4729
rect 6368 4684 6420 4690
rect 6458 4655 6514 4664
rect 6368 4626 6420 4632
rect 6472 4622 6500 4655
rect 6276 4616 6328 4622
rect 6274 4584 6276 4593
rect 6460 4616 6512 4622
rect 6328 4584 6330 4593
rect 6184 4548 6236 4554
rect 6460 4558 6512 4564
rect 6656 4554 6684 5170
rect 6274 4519 6330 4528
rect 6644 4548 6696 4554
rect 6184 4490 6236 4496
rect 6644 4490 6696 4496
rect 6196 4282 6224 4490
rect 6748 4486 6776 9046
rect 6840 8974 6868 13670
rect 6932 13530 6960 13738
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6932 11218 6960 11562
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10606 6960 10950
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 9500 6960 10542
rect 7024 9722 7052 13756
rect 7208 12646 7236 14010
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7208 12306 7236 12582
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7116 11762 7144 12106
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7208 11150 7236 12242
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7300 11082 7328 13670
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7392 12345 7420 12378
rect 7378 12336 7434 12345
rect 7378 12271 7434 12280
rect 7484 11558 7512 14350
rect 7760 13938 7788 14758
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 12481 7604 13806
rect 7562 12472 7618 12481
rect 7562 12407 7618 12416
rect 7760 12170 7788 13874
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7576 11898 7604 12106
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7576 11694 7604 11834
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7562 11520 7618 11529
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7116 10062 7144 10134
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7208 9897 7236 10542
rect 7194 9888 7250 9897
rect 7194 9823 7250 9832
rect 7300 9738 7328 11018
rect 7392 10985 7420 11222
rect 7378 10976 7434 10985
rect 7378 10911 7434 10920
rect 7484 10418 7512 11494
rect 7562 11455 7618 11464
rect 7576 11354 7604 11455
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7668 10674 7696 11834
rect 7760 10810 7788 12106
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7484 10390 7696 10418
rect 7470 10296 7526 10305
rect 7470 10231 7526 10240
rect 7484 10062 7512 10231
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7208 9710 7328 9738
rect 7208 9586 7236 9710
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6932 9472 7052 9500
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8498 6960 8910
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7024 8294 7052 9472
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 6840 8266 7052 8294
rect 6840 8129 6868 8266
rect 6826 8120 6882 8129
rect 6826 8055 6882 8064
rect 7010 8120 7066 8129
rect 7010 8055 7066 8064
rect 6840 7954 6868 8055
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 7546 6868 7754
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 7024 7313 7052 8055
rect 7116 7886 7144 8502
rect 7208 8129 7236 9522
rect 7288 9512 7340 9518
rect 7286 9480 7288 9489
rect 7340 9480 7342 9489
rect 7286 9415 7342 9424
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7300 8566 7328 9046
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7194 8120 7250 8129
rect 7194 8055 7250 8064
rect 7300 7888 7328 8230
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7288 7882 7340 7888
rect 7288 7824 7340 7830
rect 7010 7304 7066 7313
rect 7010 7239 7066 7248
rect 6826 6896 6882 6905
rect 6826 6831 6882 6840
rect 6840 6798 6868 6831
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6458 6960 6598
rect 7010 6488 7066 6497
rect 6920 6452 6972 6458
rect 7010 6423 7066 6432
rect 6920 6394 6972 6400
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6840 5409 6868 6258
rect 6932 5846 6960 6258
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6826 5400 6882 5409
rect 6826 5335 6882 5344
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 5368 4146 5396 4218
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 6288 4078 6316 4218
rect 6840 4146 6868 5335
rect 7024 5166 7052 6423
rect 7116 6322 7144 7822
rect 7194 7576 7250 7585
rect 7300 7546 7328 7824
rect 7194 7511 7250 7520
rect 7288 7540 7340 7546
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7208 5234 7236 7511
rect 7288 7482 7340 7488
rect 7300 6662 7328 7482
rect 7392 7002 7420 9930
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7484 8906 7512 9114
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7484 7888 7512 8842
rect 7576 8430 7604 9522
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 7882 7524 7888
rect 7472 7824 7524 7830
rect 7576 7868 7604 8366
rect 7668 7993 7696 10390
rect 7748 9920 7800 9926
rect 7852 9908 7880 15438
rect 7944 12434 7972 15558
rect 8036 13920 8064 15846
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 15026 8156 15302
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8128 14074 8156 14350
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8116 13932 8168 13938
rect 8036 13892 8116 13920
rect 8116 13874 8168 13880
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8036 12986 8064 13738
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7944 12406 8064 12434
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7944 11626 7972 12242
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7944 11354 7972 11562
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7930 11248 7986 11257
rect 7930 11183 7986 11192
rect 7944 10198 7972 11183
rect 7932 10192 7984 10198
rect 7932 10134 7984 10140
rect 7800 9880 7880 9908
rect 7748 9862 7800 9868
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7760 8673 7788 9658
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7930 9344 7986 9353
rect 7852 9042 7880 9318
rect 7930 9279 7986 9288
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7944 8974 7972 9279
rect 8036 9178 8064 12406
rect 8128 11898 8156 13874
rect 8220 13462 8248 14894
rect 8312 14074 8340 17190
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 15706 8432 16934
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8392 15496 8444 15502
rect 8390 15464 8392 15473
rect 8444 15464 8446 15473
rect 8390 15399 8446 15408
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8220 12850 8248 13398
rect 8312 13326 8340 13670
rect 8404 13394 8432 14962
rect 8496 14550 8524 17614
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8588 16658 8616 17070
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8496 14278 8524 14350
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8484 14000 8536 14006
rect 8588 13988 8616 16594
rect 8536 13960 8616 13988
rect 8484 13942 8536 13948
rect 8496 13433 8524 13942
rect 8482 13424 8538 13433
rect 8392 13388 8444 13394
rect 8482 13359 8538 13368
rect 8392 13330 8444 13336
rect 8300 13320 8352 13326
rect 8298 13288 8300 13297
rect 8484 13320 8536 13326
rect 8352 13288 8354 13297
rect 8298 13223 8354 13232
rect 8482 13288 8484 13297
rect 8576 13320 8628 13326
rect 8536 13288 8538 13297
rect 8576 13262 8628 13268
rect 8482 13223 8538 13232
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8206 12744 8262 12753
rect 8312 12714 8340 13126
rect 8588 12986 8616 13262
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8206 12679 8262 12688
rect 8300 12708 8352 12714
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8220 11150 8248 12679
rect 8300 12650 8352 12656
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8312 11150 8340 12650
rect 8404 12238 8432 12650
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11830 8432 12174
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10742 8156 10950
rect 8116 10736 8168 10742
rect 8116 10678 8168 10684
rect 8220 10577 8248 11086
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8206 10568 8262 10577
rect 8116 10532 8168 10538
rect 8206 10503 8262 10512
rect 8116 10474 8168 10480
rect 8128 10033 8156 10474
rect 8114 10024 8170 10033
rect 8114 9959 8170 9968
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8128 9450 8156 9862
rect 8220 9586 8248 10503
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7746 8664 7802 8673
rect 7746 8599 7802 8608
rect 7746 8528 7802 8537
rect 7746 8463 7748 8472
rect 7800 8463 7802 8472
rect 7748 8434 7800 8440
rect 7838 8392 7894 8401
rect 7838 8327 7894 8336
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7654 7984 7710 7993
rect 7654 7919 7710 7928
rect 7656 7880 7708 7886
rect 7576 7840 7656 7868
rect 7576 7732 7604 7840
rect 7656 7822 7708 7828
rect 7760 7818 7788 8230
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7484 7704 7604 7732
rect 7656 7744 7708 7750
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7392 5778 7420 6938
rect 7484 6798 7512 7704
rect 7656 7686 7708 7692
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 6798 7604 7278
rect 7668 7206 7696 7686
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7484 6186 7512 6734
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7378 5264 7434 5273
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7196 5228 7248 5234
rect 7378 5199 7380 5208
rect 7196 5170 7248 5176
rect 7432 5199 7434 5208
rect 7564 5228 7616 5234
rect 7380 5170 7432 5176
rect 7564 5170 7616 5176
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7116 4826 7144 5170
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6932 4214 6960 4558
rect 7024 4486 7052 4558
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 6840 3670 6868 4082
rect 7024 3738 7052 4422
rect 7484 4146 7512 5034
rect 7576 5030 7604 5170
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7668 4826 7696 5170
rect 7760 4826 7788 7754
rect 7852 6610 7880 8327
rect 7944 8265 7972 8774
rect 7930 8256 7986 8265
rect 7930 8191 7986 8200
rect 7944 6798 7972 8191
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7852 6582 7972 6610
rect 7838 6352 7894 6361
rect 7838 6287 7894 6296
rect 7852 6186 7880 6287
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7852 5778 7880 6122
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7852 5370 7880 5578
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7944 5030 7972 6582
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7760 4486 7788 4762
rect 7944 4622 7972 4966
rect 8036 4622 8064 9114
rect 8128 8362 8156 9386
rect 8220 8362 8248 9522
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8312 8294 8340 10950
rect 8404 10674 8432 11222
rect 8588 11150 8616 12786
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10062 8432 10406
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8574 10024 8630 10033
rect 8484 9988 8536 9994
rect 8574 9959 8576 9968
rect 8484 9930 8536 9936
rect 8628 9959 8630 9968
rect 8576 9930 8628 9936
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 8566 8432 9318
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8390 8392 8446 8401
rect 8390 8327 8392 8336
rect 8444 8327 8446 8336
rect 8392 8298 8444 8304
rect 8300 8288 8352 8294
rect 8114 8256 8170 8265
rect 8300 8230 8352 8236
rect 8114 8191 8170 8200
rect 8128 7864 8156 8191
rect 8312 7970 8340 8230
rect 8312 7942 8432 7970
rect 8404 7886 8432 7942
rect 8300 7880 8352 7886
rect 8116 7858 8168 7864
rect 8300 7822 8352 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8116 7800 8168 7806
rect 8128 7721 8156 7800
rect 8208 7744 8260 7750
rect 8114 7712 8170 7721
rect 8208 7686 8260 7692
rect 8114 7647 8170 7656
rect 8220 7449 8248 7686
rect 8206 7440 8262 7449
rect 8206 7375 8262 7384
rect 8312 7041 8340 7822
rect 8390 7304 8446 7313
rect 8390 7239 8446 7248
rect 8114 7032 8170 7041
rect 8114 6967 8170 6976
rect 8298 7032 8354 7041
rect 8298 6967 8354 6976
rect 8128 6390 8156 6967
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8220 6497 8248 6802
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8206 6488 8262 6497
rect 8206 6423 8262 6432
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8128 5778 8156 6326
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 8036 3602 8064 4558
rect 8312 4078 8340 6734
rect 8404 4214 8432 7239
rect 8496 6390 8524 9930
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8588 8974 8616 9454
rect 8680 9178 8708 17614
rect 8760 17604 8812 17610
rect 8760 17546 8812 17552
rect 8772 16182 8800 17546
rect 8852 17536 8904 17542
rect 8850 17504 8852 17513
rect 8904 17504 8906 17513
rect 8850 17439 8906 17448
rect 9048 17202 9076 17818
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9232 17338 9260 17614
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 17338 9352 17478
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9312 17332 9364 17338
rect 9600 17320 9628 18255
rect 10140 18226 10192 18232
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9784 17882 9812 18090
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9772 17332 9824 17338
rect 9600 17292 9772 17320
rect 9312 17274 9364 17280
rect 9772 17274 9824 17280
rect 9126 17232 9182 17241
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9036 17196 9088 17202
rect 9770 17232 9826 17241
rect 9126 17167 9182 17176
rect 9220 17196 9272 17202
rect 9036 17138 9088 17144
rect 8864 16697 8892 17138
rect 8956 16726 8984 17138
rect 9048 16946 9076 17138
rect 9140 17066 9168 17167
rect 9220 17138 9272 17144
rect 9312 17196 9364 17202
rect 9770 17167 9772 17176
rect 9312 17138 9364 17144
rect 9824 17167 9826 17176
rect 9772 17138 9824 17144
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9048 16918 9168 16946
rect 9140 16794 9168 16918
rect 9232 16833 9260 17138
rect 9218 16824 9274 16833
rect 9128 16788 9180 16794
rect 9324 16794 9352 17138
rect 9680 17128 9732 17134
rect 9416 17088 9680 17116
rect 9218 16759 9274 16768
rect 9312 16788 9364 16794
rect 9128 16730 9180 16736
rect 9312 16730 9364 16736
rect 8944 16720 8996 16726
rect 8850 16688 8906 16697
rect 8944 16662 8996 16668
rect 8850 16623 8906 16632
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 8852 16516 8904 16522
rect 8852 16458 8904 16464
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8772 14521 8800 15642
rect 8864 15337 8892 16458
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8850 15328 8906 15337
rect 8850 15263 8906 15272
rect 8850 15192 8906 15201
rect 8850 15127 8906 15136
rect 8758 14512 8814 14521
rect 8758 14447 8814 14456
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8772 14113 8800 14350
rect 8864 14278 8892 15127
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8758 14104 8814 14113
rect 8758 14039 8814 14048
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13530 8800 13874
rect 8864 13705 8892 14214
rect 8850 13696 8906 13705
rect 8850 13631 8906 13640
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8772 12374 8800 12650
rect 8864 12458 8892 13631
rect 8956 13274 8984 15438
rect 9036 15360 9088 15366
rect 9140 15348 9168 15506
rect 9088 15320 9168 15348
rect 9036 15302 9088 15308
rect 9140 15094 9168 15320
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9034 14376 9090 14385
rect 9034 14311 9036 14320
rect 9088 14311 9090 14320
rect 9036 14282 9088 14288
rect 9140 14278 9168 14894
rect 9232 14278 9260 16526
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9324 16017 9352 16118
rect 9310 16008 9366 16017
rect 9310 15943 9366 15952
rect 9416 15502 9444 17088
rect 9680 17070 9732 17076
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9680 16992 9732 16998
rect 9864 16992 9916 16998
rect 9732 16952 9864 16980
rect 9680 16934 9732 16940
rect 9864 16934 9916 16940
rect 9496 16584 9548 16590
rect 9494 16552 9496 16561
rect 9548 16552 9550 16561
rect 9494 16487 9550 16496
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9508 15706 9536 16050
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9496 15564 9548 15570
rect 9600 15552 9628 16934
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 15638 9720 16526
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9784 15910 9812 16458
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9876 15910 9904 16390
rect 9968 16114 9996 17614
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9680 15632 9732 15638
rect 9680 15574 9732 15580
rect 9548 15524 9628 15552
rect 9496 15506 9548 15512
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9508 15162 9536 15506
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9496 15156 9548 15162
rect 9416 15116 9496 15144
rect 9312 14884 9364 14890
rect 9312 14826 9364 14832
rect 9128 14272 9180 14278
rect 9126 14240 9128 14249
rect 9220 14272 9272 14278
rect 9180 14240 9182 14249
rect 9220 14214 9272 14220
rect 9126 14175 9182 14184
rect 9232 14090 9260 14214
rect 9140 14062 9260 14090
rect 9140 13938 9168 14062
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9048 13530 9076 13874
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9218 13424 9274 13433
rect 9218 13359 9220 13368
rect 9272 13359 9274 13368
rect 9220 13330 9272 13336
rect 8956 13246 9260 13274
rect 9232 13190 9260 13246
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9034 12608 9090 12617
rect 9034 12543 9090 12552
rect 8942 12472 8998 12481
rect 8864 12430 8942 12458
rect 9048 12442 9076 12543
rect 8942 12407 8998 12416
rect 9036 12436 9088 12442
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8956 12306 8984 12407
rect 9036 12378 9088 12384
rect 9140 12306 9168 13126
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9232 12753 9260 12786
rect 9218 12744 9274 12753
rect 9218 12679 9274 12688
rect 9218 12608 9274 12617
rect 9218 12543 9274 12552
rect 9232 12306 9260 12543
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 8850 12200 8906 12209
rect 8850 12135 8852 12144
rect 8904 12135 8906 12144
rect 8944 12164 8996 12170
rect 8852 12106 8904 12112
rect 8944 12106 8996 12112
rect 8864 11506 8892 12106
rect 8956 12073 8984 12106
rect 8942 12064 8998 12073
rect 8942 11999 8998 12008
rect 9034 11792 9090 11801
rect 9034 11727 9090 11736
rect 8864 11478 8984 11506
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8864 10849 8892 11086
rect 8850 10840 8906 10849
rect 8850 10775 8906 10784
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 10577 8892 10610
rect 8850 10568 8906 10577
rect 8850 10503 8906 10512
rect 8850 10160 8906 10169
rect 8850 10095 8906 10104
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8634 8800 8774
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8588 5914 8616 8298
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8496 5710 8524 5850
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8588 5234 8616 5714
rect 8680 5234 8708 7958
rect 8864 7886 8892 10095
rect 8956 9625 8984 11478
rect 9048 10538 9076 11727
rect 9140 11393 9168 12242
rect 9232 11529 9260 12242
rect 9218 11520 9274 11529
rect 9218 11455 9274 11464
rect 9126 11384 9182 11393
rect 9324 11354 9352 14826
rect 9416 14600 9444 15116
rect 9496 15098 9548 15104
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9508 14793 9536 14962
rect 9494 14784 9550 14793
rect 9494 14719 9550 14728
rect 9416 14572 9536 14600
rect 9402 14512 9458 14521
rect 9402 14447 9458 14456
rect 9416 12782 9444 14447
rect 9508 14414 9536 14572
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9600 14260 9628 15302
rect 9692 15162 9720 15438
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9692 14929 9720 14962
rect 9678 14920 9734 14929
rect 9678 14855 9734 14864
rect 9508 14232 9628 14260
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9416 11665 9444 12174
rect 9508 11744 9536 14232
rect 9588 13320 9640 13326
rect 9586 13288 9588 13297
rect 9640 13288 9642 13297
rect 9586 13223 9642 13232
rect 9600 12617 9628 13223
rect 9692 12986 9720 14855
rect 9784 13530 9812 15846
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9876 15026 9904 15574
rect 9968 15366 9996 16050
rect 10060 16046 10088 16390
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10060 15706 10088 15982
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 10060 15162 10088 15642
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9876 14074 9904 14962
rect 10152 14618 10180 18226
rect 10336 18222 10364 18362
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10244 17882 10272 18158
rect 11716 17882 11744 18702
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11900 18358 11928 18566
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11992 18086 12020 18158
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10232 17672 10284 17678
rect 10230 17640 10232 17649
rect 10416 17672 10468 17678
rect 10284 17640 10286 17649
rect 10416 17614 10468 17620
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10230 17575 10286 17584
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10244 16998 10272 17138
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10244 15366 10272 16526
rect 10336 16454 10364 17070
rect 10428 16794 10456 17614
rect 10612 17542 10640 17614
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10520 16794 10548 17478
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10324 16176 10376 16182
rect 10322 16144 10324 16153
rect 10376 16144 10378 16153
rect 10322 16079 10378 16088
rect 10520 16017 10548 16390
rect 10506 16008 10562 16017
rect 10416 15972 10468 15978
rect 10506 15943 10562 15952
rect 10416 15914 10468 15920
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9968 14074 9996 14282
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9862 13968 9918 13977
rect 9862 13903 9864 13912
rect 9916 13903 9918 13912
rect 9956 13932 10008 13938
rect 9864 13874 9916 13880
rect 9956 13874 10008 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9770 13424 9826 13433
rect 9770 13359 9826 13368
rect 9784 13258 9812 13359
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9876 13138 9904 13738
rect 9784 13110 9904 13138
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9586 12608 9642 12617
rect 9586 12543 9642 12552
rect 9784 12238 9812 13110
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11898 9720 12106
rect 9876 12102 9904 12650
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9680 11892 9732 11898
rect 9864 11892 9916 11898
rect 9680 11834 9732 11840
rect 9784 11852 9864 11880
rect 9508 11716 9628 11744
rect 9402 11656 9458 11665
rect 9402 11591 9458 11600
rect 9126 11319 9182 11328
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9220 11280 9272 11286
rect 9140 11240 9220 11268
rect 9140 10606 9168 11240
rect 9220 11222 9272 11228
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9048 10266 9076 10474
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9232 10198 9260 10950
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 8942 9616 8998 9625
rect 9232 9586 9260 10134
rect 8942 9551 8998 9560
rect 9220 9580 9272 9586
rect 8956 9518 8984 9551
rect 9220 9522 9272 9528
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 8673 8984 8910
rect 9034 8800 9090 8809
rect 9034 8735 9090 8744
rect 8942 8664 8998 8673
rect 8942 8599 8998 8608
rect 8956 8566 8984 8599
rect 9048 8566 9076 8735
rect 8944 8560 8996 8566
rect 8944 8502 8996 8508
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8956 8090 8984 8366
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9048 8265 9076 8298
rect 9034 8256 9090 8265
rect 9034 8191 9090 8200
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8944 7744 8996 7750
rect 8850 7712 8906 7721
rect 8944 7686 8996 7692
rect 8850 7647 8906 7656
rect 8956 7670 8985 7686
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8772 6458 8800 7346
rect 8864 7177 8892 7647
rect 8956 7449 8984 7670
rect 8942 7440 8998 7449
rect 9048 7410 9076 7822
rect 9140 7449 9168 8434
rect 9232 8412 9260 9522
rect 9324 9178 9352 11290
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9402 10296 9458 10305
rect 9402 10231 9404 10240
rect 9456 10231 9458 10240
rect 9404 10202 9456 10208
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9416 9926 9444 10066
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9508 9722 9536 11154
rect 9600 11150 9628 11716
rect 9588 11144 9640 11150
rect 9680 11144 9732 11150
rect 9588 11086 9640 11092
rect 9678 11112 9680 11121
rect 9732 11112 9734 11121
rect 9678 11047 9734 11056
rect 9784 11014 9812 11852
rect 9864 11834 9916 11840
rect 9968 11762 9996 13874
rect 10060 13326 10088 13874
rect 10244 13802 10272 15302
rect 10336 15201 10364 15438
rect 10428 15434 10456 15914
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10322 15192 10378 15201
rect 10322 15127 10378 15136
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10336 13841 10364 14962
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10428 14414 10456 14758
rect 10520 14521 10548 14962
rect 10506 14512 10562 14521
rect 10506 14447 10562 14456
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 14074 10548 14350
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10416 13864 10468 13870
rect 10322 13832 10378 13841
rect 10232 13796 10284 13802
rect 10416 13806 10468 13812
rect 10322 13767 10378 13776
rect 10232 13738 10284 13744
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10060 11762 10088 12922
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10244 12238 10272 12378
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9876 11642 9904 11698
rect 9876 11614 9996 11642
rect 9862 11520 9918 11529
rect 9862 11455 9918 11464
rect 9876 11014 9904 11455
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9600 9586 9628 10542
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 9382 9628 9522
rect 9588 9376 9640 9382
rect 9508 9336 9588 9364
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9416 8974 9444 9046
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9310 8800 9366 8809
rect 9310 8735 9366 8744
rect 9324 8634 9352 8735
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9416 8480 9444 8910
rect 9400 8452 9444 8480
rect 9400 8412 9428 8452
rect 9232 8384 9286 8412
rect 9400 8384 9444 8412
rect 9258 8294 9286 8384
rect 9232 8266 9286 8294
rect 9126 7440 9182 7449
rect 8942 7375 8998 7384
rect 9036 7404 9088 7410
rect 9126 7375 9182 7384
rect 9036 7346 9088 7352
rect 9036 7200 9088 7206
rect 8850 7168 8906 7177
rect 8850 7103 8906 7112
rect 9034 7168 9036 7177
rect 9088 7168 9090 7177
rect 9034 7103 9090 7112
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8772 5914 8800 6258
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8864 5710 8892 7103
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8944 6384 8996 6390
rect 8942 6352 8944 6361
rect 8996 6352 8998 6361
rect 8942 6287 8998 6296
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8944 6248 8996 6254
rect 9048 6225 9076 6258
rect 9140 6254 9168 6394
rect 9128 6248 9180 6254
rect 8944 6190 8996 6196
rect 9034 6216 9090 6225
rect 8956 5914 8984 6190
rect 9128 6190 9180 6196
rect 9034 6151 9090 6160
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8588 5030 8616 5170
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8680 4690 8708 5170
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8864 4826 8892 5102
rect 8956 4826 8984 5238
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8574 4584 8630 4593
rect 8574 4519 8630 4528
rect 8588 4486 8616 4519
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8300 4072 8352 4078
rect 8680 4026 8708 4626
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8772 4214 8800 4490
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8300 4014 8352 4020
rect 8588 4010 8708 4026
rect 8576 4004 8708 4010
rect 8628 3998 8708 4004
rect 8576 3946 8628 3952
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 9048 2446 9076 6054
rect 9140 5846 9168 6054
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9140 4622 9168 5238
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 4486 9168 4558
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9232 4146 9260 8266
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 5846 9352 6598
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9416 5642 9444 8384
rect 9508 7886 9536 9336
rect 9588 9318 9640 9324
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8566 9628 8842
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9586 8120 9642 8129
rect 9586 8055 9588 8064
rect 9640 8055 9642 8064
rect 9588 8026 9640 8032
rect 9586 7984 9642 7993
rect 9586 7919 9642 7928
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9508 6798 9536 7822
rect 9600 6882 9628 7919
rect 9692 7002 9720 9318
rect 9784 8956 9812 10950
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9876 10266 9904 10746
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9968 10146 9996 11614
rect 9876 10130 9996 10146
rect 9864 10124 9996 10130
rect 9916 10118 9996 10124
rect 9864 10066 9916 10072
rect 9956 10056 10008 10062
rect 9862 10024 9918 10033
rect 9956 9998 10008 10004
rect 9862 9959 9864 9968
rect 9916 9959 9918 9968
rect 9864 9930 9916 9936
rect 9968 9450 9996 9998
rect 10060 9654 10088 11698
rect 10138 11248 10194 11257
rect 10138 11183 10140 11192
rect 10192 11183 10194 11192
rect 10140 11154 10192 11160
rect 10244 11150 10272 12038
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10244 10441 10272 10678
rect 10336 10470 10364 13466
rect 10428 13462 10456 13806
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10414 13288 10470 13297
rect 10414 13223 10470 13232
rect 10428 12714 10456 13223
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10324 10464 10376 10470
rect 10230 10432 10286 10441
rect 10324 10406 10376 10412
rect 10230 10367 10286 10376
rect 10138 10160 10194 10169
rect 10138 10095 10194 10104
rect 10324 10124 10376 10130
rect 10152 10062 10180 10095
rect 10324 10066 10376 10072
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9956 8968 10008 8974
rect 9784 8928 9956 8956
rect 9956 8910 10008 8916
rect 9956 8832 10008 8838
rect 9954 8800 9956 8809
rect 10008 8800 10010 8809
rect 9954 8735 10010 8744
rect 9862 8664 9918 8673
rect 9862 8599 9864 8608
rect 9916 8599 9918 8608
rect 9864 8570 9916 8576
rect 9862 8528 9918 8537
rect 9862 8463 9864 8472
rect 9916 8463 9918 8472
rect 9864 8434 9916 8440
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9600 6854 9720 6882
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9600 6458 9628 6666
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9402 5400 9458 5409
rect 9508 5370 9536 6258
rect 9600 5914 9628 6258
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9402 5335 9458 5344
rect 9496 5364 9548 5370
rect 9416 5098 9444 5335
rect 9496 5306 9548 5312
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4622 9352 4966
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9600 4162 9628 5714
rect 9692 5114 9720 6854
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 5370 9812 6802
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9692 5086 9812 5114
rect 9876 5098 9904 8434
rect 9968 7970 9996 8735
rect 10060 8498 10088 9590
rect 10152 8974 10180 9862
rect 10244 9722 10272 9998
rect 10336 9926 10364 10066
rect 10324 9920 10376 9926
rect 10322 9888 10324 9897
rect 10376 9888 10378 9897
rect 10322 9823 10378 9832
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10428 9586 10456 12650
rect 10612 12442 10640 17478
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16590 10732 16934
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10796 16250 10824 17682
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10968 17672 11020 17678
rect 11244 17672 11296 17678
rect 10968 17614 11020 17620
rect 11242 17640 11244 17649
rect 11520 17672 11572 17678
rect 11296 17640 11298 17649
rect 10888 16697 10916 17614
rect 10980 17542 11008 17614
rect 11520 17614 11572 17620
rect 11242 17575 11298 17584
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 10874 16688 10930 16697
rect 10874 16623 10930 16632
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10876 16176 10928 16182
rect 10690 16144 10746 16153
rect 10876 16118 10928 16124
rect 10690 16079 10746 16088
rect 10704 15910 10732 16079
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10796 15722 10824 15982
rect 10704 15694 10824 15722
rect 10888 15706 10916 16118
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10876 15700 10928 15706
rect 10704 14958 10732 15694
rect 10876 15642 10928 15648
rect 10876 15496 10928 15502
rect 10874 15464 10876 15473
rect 10928 15464 10930 15473
rect 10874 15399 10930 15408
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10888 14498 10916 15098
rect 10980 14618 11008 15982
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11072 14822 11100 15438
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10888 14470 11008 14498
rect 10980 14346 11008 14470
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10796 13326 10824 13874
rect 10784 13320 10836 13326
rect 10704 13280 10784 13308
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10506 11248 10562 11257
rect 10506 11183 10562 11192
rect 10520 11150 10548 11183
rect 10508 11144 10560 11150
rect 10600 11144 10652 11150
rect 10508 11086 10560 11092
rect 10598 11112 10600 11121
rect 10652 11112 10654 11121
rect 10598 11047 10654 11056
rect 10598 10976 10654 10985
rect 10598 10911 10654 10920
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 10062 10548 10406
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10520 9926 10548 9998
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10506 9752 10562 9761
rect 10506 9687 10562 9696
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10230 9344 10286 9353
rect 10230 9279 10286 9288
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9968 7942 10088 7970
rect 10060 7886 10088 7942
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9968 7546 9996 7822
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9968 7206 9996 7482
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6497 9996 6598
rect 9954 6488 10010 6497
rect 9954 6423 10010 6432
rect 9968 5574 9996 6423
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 10060 5409 10088 7346
rect 10152 7342 10180 8910
rect 10244 8090 10272 9279
rect 10322 8936 10378 8945
rect 10322 8871 10378 8880
rect 10336 8838 10364 8871
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10324 8492 10376 8498
rect 10428 8480 10456 9386
rect 10520 8650 10548 9687
rect 10612 8974 10640 10911
rect 10704 10606 10732 13280
rect 10784 13262 10836 13268
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12986 10916 13126
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10796 12714 10824 12786
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10704 10033 10732 10066
rect 10796 10062 10824 12650
rect 10888 11150 10916 12786
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10674 10916 11086
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10888 10169 10916 10610
rect 10874 10160 10930 10169
rect 10874 10095 10930 10104
rect 10784 10056 10836 10062
rect 10690 10024 10746 10033
rect 10980 10010 11008 14282
rect 11072 13938 11100 14758
rect 11164 14346 11192 16050
rect 11256 15434 11284 16594
rect 11348 16250 11376 17478
rect 11532 16250 11560 17614
rect 11992 17610 12020 18022
rect 12636 17610 12664 18838
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 13360 18420 13412 18426
rect 13280 18380 13360 18408
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13004 17882 13032 18226
rect 13188 17882 13216 18226
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13280 17814 13308 18380
rect 13360 18362 13412 18368
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13740 17882 13768 18294
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 11704 17604 11756 17610
rect 11980 17604 12032 17610
rect 11756 17564 11980 17592
rect 11704 17546 11756 17552
rect 11980 17546 12032 17552
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12268 17338 12296 17478
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12070 17232 12126 17241
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11980 17196 12032 17202
rect 12070 17167 12072 17176
rect 11980 17138 12032 17144
rect 12124 17167 12126 17176
rect 12072 17138 12124 17144
rect 11716 17105 11744 17138
rect 11702 17096 11758 17105
rect 11612 17060 11664 17066
rect 11992 17066 12020 17138
rect 11702 17031 11758 17040
rect 11980 17060 12032 17066
rect 11612 17002 11664 17008
rect 11980 17002 12032 17008
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11348 14498 11376 16050
rect 11440 15570 11468 16118
rect 11624 15960 11652 17002
rect 12084 16794 12112 17138
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12348 16720 12400 16726
rect 12348 16662 12400 16668
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 16046 11744 16390
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11532 15932 11652 15960
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11532 15502 11560 15932
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11704 15496 11756 15502
rect 11808 15484 11836 16594
rect 11886 15872 11942 15881
rect 11886 15807 11942 15816
rect 11900 15502 11928 15807
rect 11756 15456 11836 15484
rect 11888 15496 11940 15502
rect 11704 15438 11756 15444
rect 11888 15438 11940 15444
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11256 14470 11376 14498
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13161 11192 13670
rect 11150 13152 11206 13161
rect 11150 13087 11206 13096
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11072 12306 11100 12854
rect 11150 12472 11206 12481
rect 11150 12407 11206 12416
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10784 9998 10836 10004
rect 10690 9959 10746 9968
rect 10888 9982 11008 10010
rect 11072 9994 11100 12242
rect 11164 12238 11192 12407
rect 11152 12232 11204 12238
rect 11256 12209 11284 14470
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 13297 11376 14350
rect 11428 14272 11480 14278
rect 11426 14240 11428 14249
rect 11520 14272 11572 14278
rect 11480 14240 11482 14249
rect 11520 14214 11572 14220
rect 11426 14175 11482 14184
rect 11440 13818 11468 14175
rect 11532 13938 11560 14214
rect 11624 14074 11652 14486
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11716 13938 11744 14894
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11440 13790 11560 13818
rect 11334 13288 11390 13297
rect 11334 13223 11390 13232
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11152 12174 11204 12180
rect 11242 12200 11298 12209
rect 11164 11937 11192 12174
rect 11242 12135 11298 12144
rect 11150 11928 11206 11937
rect 11150 11863 11206 11872
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11060 9988 11112 9994
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10520 8622 10640 8650
rect 10508 8492 10560 8498
rect 10428 8452 10508 8480
rect 10324 8434 10376 8440
rect 10508 8434 10560 8440
rect 10336 8401 10364 8434
rect 10322 8392 10378 8401
rect 10322 8327 10378 8336
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10428 7993 10456 8298
rect 10414 7984 10470 7993
rect 10414 7919 10470 7928
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 10244 7274 10272 7482
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10336 6914 10364 7754
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 6934 10456 7686
rect 10520 7478 10548 8434
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10244 6886 10364 6914
rect 10416 6928 10468 6934
rect 10244 6730 10272 6886
rect 10416 6870 10468 6876
rect 10520 6798 10548 7142
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10508 6792 10560 6798
rect 10612 6769 10640 8622
rect 10704 8498 10732 9114
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10690 8256 10746 8265
rect 10690 8191 10746 8200
rect 10704 7818 10732 8191
rect 10796 8022 10824 8774
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10888 7818 10916 9982
rect 11060 9930 11112 9936
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10692 7812 10744 7818
rect 10876 7812 10928 7818
rect 10692 7754 10744 7760
rect 10796 7772 10876 7800
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10704 7002 10732 7210
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10508 6734 10560 6740
rect 10598 6760 10654 6769
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10140 6384 10192 6390
rect 10138 6352 10140 6361
rect 10428 6361 10456 6734
rect 10192 6352 10194 6361
rect 10138 6287 10194 6296
rect 10414 6352 10470 6361
rect 10414 6287 10470 6296
rect 10520 5914 10548 6734
rect 10598 6695 10654 6704
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10322 5808 10378 5817
rect 10322 5743 10324 5752
rect 10376 5743 10378 5752
rect 10324 5714 10376 5720
rect 10232 5568 10284 5574
rect 10138 5536 10194 5545
rect 10232 5510 10284 5516
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10138 5471 10194 5480
rect 10046 5400 10102 5409
rect 10046 5335 10102 5344
rect 10060 5234 10088 5335
rect 10152 5302 10180 5471
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10244 5234 10272 5510
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9508 4134 9628 4162
rect 9508 4078 9536 4134
rect 9692 4078 9720 4966
rect 9784 4826 9812 5086
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 10138 4856 10194 4865
rect 9772 4820 9824 4826
rect 10138 4791 10194 4800
rect 9772 4762 9824 4768
rect 10152 4690 10180 4791
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9784 3942 9812 4422
rect 10152 4282 10180 4626
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 4282 10272 4422
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10336 4078 10364 5510
rect 10520 5098 10548 5850
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10428 4978 10456 5034
rect 10612 4978 10640 6695
rect 10796 6254 10824 7772
rect 10876 7754 10928 7760
rect 10980 7290 11008 9862
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 9489 11100 9522
rect 11058 9480 11114 9489
rect 11164 9450 11192 11630
rect 11058 9415 11114 9424
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11058 9208 11114 9217
rect 11058 9143 11060 9152
rect 11112 9143 11114 9152
rect 11060 9114 11112 9120
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 11072 8673 11100 8842
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11058 8664 11114 8673
rect 11164 8634 11192 8774
rect 11058 8599 11114 8608
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11150 8392 11206 8401
rect 11150 8327 11206 8336
rect 11058 7984 11114 7993
rect 11058 7919 11114 7928
rect 10888 7262 11008 7290
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10428 4950 10640 4978
rect 10704 4826 10732 6054
rect 10796 5778 10824 6190
rect 10888 6118 10916 7262
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 7002 11008 7142
rect 11072 7002 11100 7919
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11058 6896 11114 6905
rect 10980 6854 11058 6882
rect 10980 6730 11008 6854
rect 11164 6882 11192 8327
rect 11256 7886 11284 11834
rect 11348 11529 11376 12718
rect 11532 12322 11560 13790
rect 11716 12458 11744 13874
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11716 12430 11745 12458
rect 11717 12356 11745 12430
rect 11440 12294 11560 12322
rect 11624 12328 11745 12356
rect 11440 11898 11468 12294
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11532 11898 11560 12174
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11520 11552 11572 11558
rect 11334 11520 11390 11529
rect 11520 11494 11572 11500
rect 11334 11455 11390 11464
rect 11348 10062 11376 11455
rect 11532 11286 11560 11494
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11348 9674 11376 9998
rect 11348 9646 11468 9674
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11348 8498 11376 9046
rect 11440 8498 11468 9646
rect 11520 9376 11572 9382
rect 11518 9344 11520 9353
rect 11572 9344 11574 9353
rect 11518 9279 11574 9288
rect 11532 8566 11560 9279
rect 11624 8673 11652 12328
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11830 11744 12174
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11716 11354 11744 11630
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11610 8664 11666 8673
rect 11610 8599 11666 8608
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 7410 11284 7822
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11164 6854 11284 6882
rect 11058 6831 11114 6840
rect 11256 6798 11284 6854
rect 11060 6792 11112 6798
rect 11244 6792 11296 6798
rect 11112 6752 11192 6780
rect 11060 6734 11112 6740
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10966 5808 11022 5817
rect 10784 5772 10836 5778
rect 10966 5743 11022 5752
rect 10784 5714 10836 5720
rect 10980 5710 11008 5743
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 10874 5400 10930 5409
rect 10874 5335 10930 5344
rect 10888 5234 10916 5335
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 11072 4826 11100 5578
rect 11164 5148 11192 6752
rect 11244 6734 11296 6740
rect 11256 5216 11284 6734
rect 11348 6322 11376 8026
rect 11440 7392 11468 8434
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 8090 11560 8230
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11440 7364 11560 7392
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11440 6390 11468 6870
rect 11532 6390 11560 7364
rect 11624 6798 11652 8298
rect 11716 8090 11744 11290
rect 11808 11098 11836 13126
rect 11992 12424 12020 16594
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12072 16176 12124 16182
rect 12070 16144 12072 16153
rect 12124 16144 12126 16153
rect 12070 16079 12126 16088
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 14618 12112 15982
rect 12164 15904 12216 15910
rect 12268 15881 12296 16526
rect 12360 16425 12388 16662
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12346 16416 12402 16425
rect 12346 16351 12402 16360
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12164 15846 12216 15852
rect 12254 15872 12310 15881
rect 12176 15706 12204 15846
rect 12254 15807 12310 15816
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 15026 12204 15438
rect 12268 15366 12296 15642
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13326 12112 14010
rect 12176 13938 12204 14826
rect 12360 14822 12388 16118
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12254 14648 12310 14657
rect 12254 14583 12310 14592
rect 12268 14498 12296 14583
rect 12452 14498 12480 16594
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12544 15094 12572 15370
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12268 14470 12572 14498
rect 12268 14414 12296 14470
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12254 14104 12310 14113
rect 12360 14074 12388 14350
rect 12254 14039 12310 14048
rect 12348 14068 12400 14074
rect 12268 14006 12296 14039
rect 12348 14010 12400 14016
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12176 13734 12204 13874
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12268 13326 12296 13942
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12348 13864 12400 13870
rect 12346 13832 12348 13841
rect 12400 13832 12402 13841
rect 12452 13802 12480 13874
rect 12346 13767 12402 13776
rect 12440 13796 12492 13802
rect 12440 13738 12492 13744
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12360 13376 12388 13670
rect 12440 13388 12492 13394
rect 12360 13348 12440 13376
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12084 12714 12112 12854
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 12176 12434 12204 13126
rect 12360 12918 12388 13348
rect 12440 13330 12492 13336
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12544 12782 12572 14470
rect 12636 14414 12664 14758
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12622 13968 12678 13977
rect 12622 13903 12624 13912
rect 12676 13903 12678 13912
rect 12624 13874 12676 13880
rect 12636 13734 12664 13874
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12728 13546 12756 17614
rect 13280 17542 13308 17750
rect 13924 17678 13952 18702
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14384 17746 14412 18022
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17270 13308 17478
rect 14108 17338 14136 17614
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12820 16794 12848 17070
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 13176 16584 13228 16590
rect 13174 16552 13176 16561
rect 13268 16584 13320 16590
rect 13228 16552 13230 16561
rect 13268 16526 13320 16532
rect 13174 16487 13230 16496
rect 13188 16289 13216 16487
rect 13174 16280 13230 16289
rect 13280 16250 13308 16526
rect 13174 16215 13230 16224
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 12900 15360 12952 15366
rect 13096 15337 13124 15642
rect 12900 15302 12952 15308
rect 13082 15328 13138 15337
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12820 14550 12848 14962
rect 12912 14958 12940 15302
rect 13082 15263 13138 15272
rect 13096 15026 13124 15263
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12912 14600 12940 14894
rect 12912 14572 13124 14600
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 13938 12848 14350
rect 12898 14104 12954 14113
rect 12898 14039 12900 14048
rect 12952 14039 12954 14048
rect 12900 14010 12952 14016
rect 13004 13938 13032 14418
rect 12808 13932 12860 13938
rect 12992 13932 13044 13938
rect 12808 13874 12860 13880
rect 12912 13892 12992 13920
rect 12636 13518 12756 13546
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 11900 12396 12020 12424
rect 12084 12406 12204 12434
rect 12254 12472 12310 12481
rect 12254 12407 12310 12416
rect 11900 12306 11928 12396
rect 11978 12336 12034 12345
rect 11888 12300 11940 12306
rect 11978 12271 12034 12280
rect 11888 12242 11940 12248
rect 11992 12238 12020 12271
rect 11980 12232 12032 12238
rect 11886 12200 11942 12209
rect 11980 12174 12032 12180
rect 11886 12135 11888 12144
rect 11940 12135 11942 12144
rect 11888 12106 11940 12112
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11886 11928 11942 11937
rect 11886 11863 11942 11872
rect 11900 11762 11928 11863
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11992 11218 12020 12038
rect 12084 11354 12112 12406
rect 12268 12374 12296 12407
rect 12164 12368 12216 12374
rect 12162 12336 12164 12345
rect 12256 12368 12308 12374
rect 12216 12336 12218 12345
rect 12256 12310 12308 12316
rect 12162 12271 12218 12280
rect 12164 12232 12216 12238
rect 12440 12232 12492 12238
rect 12216 12192 12388 12220
rect 12164 12174 12216 12180
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11808 11070 12020 11098
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11808 10062 11836 10950
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11900 10266 11928 10610
rect 11992 10606 12020 11070
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 12084 10266 12112 10610
rect 12176 10538 12204 11562
rect 12164 10532 12216 10538
rect 12164 10474 12216 10480
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12176 10146 12204 10474
rect 12084 10118 12204 10146
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11702 7984 11758 7993
rect 11702 7919 11704 7928
rect 11756 7919 11758 7928
rect 11704 7890 11756 7896
rect 11808 7546 11836 9998
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 8498 11928 9522
rect 11978 9480 12034 9489
rect 11978 9415 12034 9424
rect 11992 9110 12020 9415
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8498 12020 8774
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11900 8401 11928 8434
rect 11886 8392 11942 8401
rect 11886 8327 11942 8336
rect 12084 7886 12112 10118
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12176 9110 12204 9386
rect 12268 9217 12296 9590
rect 12254 9208 12310 9217
rect 12254 9143 12310 9152
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12268 8809 12296 8978
rect 12254 8800 12310 8809
rect 12254 8735 12310 8744
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12176 7886 12204 8026
rect 12268 7886 12296 8735
rect 12360 8498 12388 12192
rect 12440 12174 12492 12180
rect 12452 11354 12480 12174
rect 12544 11665 12572 12718
rect 12530 11656 12586 11665
rect 12530 11591 12586 11600
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12452 9586 12480 11154
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12176 7750 12204 7822
rect 12268 7750 12296 7822
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11348 5370 11376 6258
rect 11532 6225 11560 6326
rect 11624 6254 11652 6598
rect 11808 6304 11836 7482
rect 12268 7392 12296 7686
rect 12360 7449 12388 8434
rect 12084 7364 12296 7392
rect 12346 7440 12402 7449
rect 12346 7375 12402 7384
rect 11888 6316 11940 6322
rect 11808 6276 11888 6304
rect 11888 6258 11940 6264
rect 11612 6248 11664 6254
rect 11518 6216 11574 6225
rect 12084 6202 12112 7364
rect 12360 6746 12388 7375
rect 11612 6190 11664 6196
rect 11518 6151 11574 6160
rect 11808 6174 12112 6202
rect 12176 6718 12388 6746
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11808 5302 11836 6174
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11256 5188 11468 5216
rect 11164 5120 11376 5148
rect 11348 5030 11376 5120
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10598 4720 10654 4729
rect 11348 4690 11376 4966
rect 11440 4690 11468 5188
rect 11808 5148 11836 5238
rect 12084 5216 12112 5510
rect 11992 5188 12112 5216
rect 11888 5160 11940 5166
rect 11808 5120 11888 5148
rect 11888 5102 11940 5108
rect 11518 4856 11574 4865
rect 11518 4791 11574 4800
rect 11796 4820 11848 4826
rect 10598 4655 10654 4664
rect 11336 4684 11388 4690
rect 10612 4554 10640 4655
rect 11336 4626 11388 4632
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11532 4622 11560 4791
rect 11796 4762 11848 4768
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 10704 4214 10732 4558
rect 11256 4282 11284 4558
rect 11808 4282 11836 4762
rect 11900 4690 11928 5102
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10324 4072 10376 4078
rect 10520 4049 10548 4082
rect 10324 4014 10376 4020
rect 10506 4040 10562 4049
rect 10506 3975 10562 3984
rect 9772 3936 9824 3942
rect 10508 3936 10560 3942
rect 9772 3878 9824 3884
rect 10506 3904 10508 3913
rect 10560 3904 10562 3913
rect 10506 3839 10562 3848
rect 11992 2446 12020 5188
rect 12176 4690 12204 6718
rect 12452 6372 12480 9522
rect 12544 9382 12572 11494
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12544 9042 12572 9114
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 7886 12572 8434
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12544 7478 12572 7822
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12452 6344 12572 6372
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12268 5302 12296 6258
rect 12346 6216 12402 6225
rect 12346 6151 12402 6160
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 4282 12112 4558
rect 12268 4486 12296 4966
rect 12360 4758 12388 6151
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12452 5302 12480 5510
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12544 4826 12572 6344
rect 12636 5710 12664 13518
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12850 12756 13126
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12728 12442 12756 12786
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12728 11898 12756 12106
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12820 11218 12848 13874
rect 12912 12850 12940 13892
rect 12992 13874 13044 13880
rect 13096 13802 13124 14572
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 14006 13216 14214
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 11937 12940 12786
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13096 12481 13124 12718
rect 13082 12472 13138 12481
rect 13082 12407 13138 12416
rect 13188 12306 13216 13942
rect 13280 13326 13308 16186
rect 13556 16114 13584 16934
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 16250 13952 16594
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 14016 16182 14044 16390
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13280 12850 13308 13262
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13372 12434 13400 15438
rect 13464 15366 13492 16050
rect 13556 15978 13584 16050
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13464 13394 13492 14894
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13556 13190 13584 15914
rect 13924 15609 13952 16050
rect 14002 16008 14058 16017
rect 14002 15943 14058 15952
rect 14016 15910 14044 15943
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13726 15600 13782 15609
rect 13726 15535 13782 15544
rect 13910 15600 13966 15609
rect 13910 15535 13966 15544
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13280 12406 13400 12434
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 12990 12200 13046 12209
rect 12990 12135 12992 12144
rect 13044 12135 13046 12144
rect 12992 12106 13044 12112
rect 12898 11928 12954 11937
rect 12898 11863 12954 11872
rect 13280 11778 13308 12406
rect 13450 11928 13506 11937
rect 13450 11863 13506 11872
rect 13464 11830 13492 11863
rect 12912 11762 13308 11778
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 12912 11756 13320 11762
rect 12912 11750 13268 11756
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12728 9586 12756 11086
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12820 9450 12848 9862
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 8022 12756 9318
rect 12820 8498 12848 9386
rect 12912 8945 12940 11750
rect 13268 11698 13320 11704
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13082 11656 13138 11665
rect 13082 11591 13138 11600
rect 13266 11656 13322 11665
rect 13372 11626 13400 11698
rect 13266 11591 13322 11600
rect 13360 11620 13412 11626
rect 13096 11218 13124 11591
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 13096 9926 13124 11154
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13174 9752 13230 9761
rect 12992 9716 13044 9722
rect 13174 9687 13230 9696
rect 12992 9658 13044 9664
rect 13004 9382 13032 9658
rect 13188 9586 13216 9687
rect 13176 9580 13228 9586
rect 13084 9570 13136 9576
rect 13176 9522 13228 9528
rect 13084 9512 13136 9518
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12898 8936 12954 8945
rect 12898 8871 12954 8880
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12808 8492 12860 8498
rect 12912 8480 12940 8774
rect 13004 8634 13032 9318
rect 13096 8974 13124 9512
rect 13188 9489 13216 9522
rect 13174 9480 13230 9489
rect 13174 9415 13230 9424
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12912 8452 13032 8480
rect 12808 8434 12860 8440
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12912 8090 12940 8298
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12728 7449 12756 7822
rect 12714 7440 12770 7449
rect 12714 7375 12770 7384
rect 12728 7041 12756 7375
rect 12820 7177 12848 7822
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12912 7478 12940 7754
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12806 7168 12862 7177
rect 12806 7103 12862 7112
rect 12714 7032 12770 7041
rect 12714 6967 12770 6976
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12912 6322 12940 6666
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12636 5234 12664 5646
rect 12728 5386 12756 5714
rect 12728 5370 12848 5386
rect 12728 5364 12860 5370
rect 12728 5358 12808 5364
rect 12808 5306 12860 5312
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 13004 4842 13032 8452
rect 13096 8430 13124 8910
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13096 7002 13124 8366
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13188 5710 13216 8774
rect 13280 7449 13308 11591
rect 13360 11562 13412 11568
rect 13372 9722 13400 11562
rect 13464 11150 13492 11766
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13556 11529 13584 11698
rect 13542 11520 13598 11529
rect 13542 11455 13598 11464
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13544 9512 13596 9518
rect 13648 9489 13676 13670
rect 13740 12764 13768 15535
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13924 13841 13952 14010
rect 14016 13938 14044 15846
rect 14108 15502 14136 17274
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14200 16522 14228 17138
rect 14476 16658 14504 17818
rect 15028 17746 15056 18158
rect 15120 17882 15148 18158
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14568 16538 14596 17138
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 14476 16510 14596 16538
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14200 15162 14228 16458
rect 14278 16416 14334 16425
rect 14278 16351 14334 16360
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14292 15042 14320 16351
rect 14476 16182 14504 16510
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14568 16250 14596 16390
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14292 15026 14412 15042
rect 14292 15020 14424 15026
rect 14292 15014 14372 15020
rect 14372 14962 14424 14968
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13910 13832 13966 13841
rect 13820 13796 13872 13802
rect 13910 13767 13912 13776
rect 13820 13738 13872 13744
rect 13964 13767 13966 13776
rect 13912 13738 13964 13744
rect 13832 13462 13860 13738
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13924 12986 13952 13126
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 14016 12866 14044 13126
rect 13924 12850 14044 12866
rect 13912 12844 14044 12850
rect 13964 12838 14044 12844
rect 13912 12786 13964 12792
rect 13820 12776 13872 12782
rect 13740 12736 13820 12764
rect 13820 12718 13872 12724
rect 14108 12306 14136 14282
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14188 13864 14240 13870
rect 14292 13841 14320 14010
rect 14188 13806 14240 13812
rect 14278 13832 14334 13841
rect 14096 12300 14148 12306
rect 14016 12260 14096 12288
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11150 13768 11494
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 14016 10674 14044 12260
rect 14096 12242 14148 12248
rect 14200 12170 14228 13806
rect 14278 13767 14334 13776
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14292 12646 14320 12854
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 11898 14228 12106
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13544 9454 13596 9460
rect 13634 9480 13690 9489
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 9110 13400 9386
rect 13556 9353 13584 9454
rect 13634 9415 13690 9424
rect 13636 9376 13688 9382
rect 13542 9344 13598 9353
rect 13636 9318 13688 9324
rect 13542 9279 13598 9288
rect 13542 9208 13598 9217
rect 13452 9172 13504 9178
rect 13542 9143 13598 9152
rect 13452 9114 13504 9120
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13266 7440 13322 7449
rect 13266 7375 13322 7384
rect 13464 7290 13492 9114
rect 13556 8430 13584 9143
rect 13648 9042 13676 9318
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13740 7886 13768 8298
rect 13728 7880 13780 7886
rect 13542 7848 13598 7857
rect 13728 7822 13780 7828
rect 13542 7783 13544 7792
rect 13596 7783 13598 7792
rect 13636 7812 13688 7818
rect 13544 7754 13596 7760
rect 13636 7754 13688 7760
rect 13648 7546 13676 7754
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13280 7262 13492 7290
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13280 7206 13308 7262
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13280 6497 13308 7142
rect 13372 6662 13400 7142
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13266 6488 13322 6497
rect 13266 6423 13322 6432
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13280 5914 13308 6258
rect 13464 6254 13492 6938
rect 13556 6934 13584 7278
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13740 6458 13768 7822
rect 13832 7546 13860 10542
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13924 8498 13952 9930
rect 14016 9586 14044 10610
rect 14108 10470 14136 10950
rect 14200 10810 14228 11086
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14108 9897 14136 9930
rect 14094 9888 14150 9897
rect 14094 9823 14150 9832
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13452 6248 13504 6254
rect 13728 6248 13780 6254
rect 13452 6190 13504 6196
rect 13726 6216 13728 6225
rect 13780 6216 13782 6225
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13358 5808 13414 5817
rect 13358 5743 13414 5752
rect 13372 5710 13400 5743
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13188 5234 13216 5646
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12912 4814 13032 4842
rect 12348 4752 12400 4758
rect 12440 4752 12492 4758
rect 12348 4694 12400 4700
rect 12438 4720 12440 4729
rect 12492 4720 12494 4729
rect 12438 4655 12494 4664
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12544 4282 12572 4762
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12912 4026 12940 4814
rect 13464 4554 13492 6190
rect 13726 6151 13782 6160
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5642 13676 6054
rect 13740 5658 13768 6151
rect 13740 5642 13860 5658
rect 13636 5636 13688 5642
rect 13740 5636 13872 5642
rect 13740 5630 13820 5636
rect 13636 5578 13688 5584
rect 13820 5578 13872 5584
rect 13728 5568 13780 5574
rect 13924 5545 13952 8434
rect 14016 7585 14044 9522
rect 14002 7576 14058 7585
rect 14002 7511 14058 7520
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 13728 5510 13780 5516
rect 13910 5536 13966 5545
rect 13636 5228 13688 5234
rect 13740 5216 13768 5510
rect 13910 5471 13966 5480
rect 13688 5188 13768 5216
rect 13912 5228 13964 5234
rect 13636 5170 13688 5176
rect 13912 5170 13964 5176
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13832 4622 13860 5034
rect 13924 4690 13952 5170
rect 14016 5166 14044 6870
rect 14108 6390 14136 9823
rect 14200 9178 14228 10746
rect 14292 9382 14320 12582
rect 14384 11150 14412 14962
rect 14464 14952 14516 14958
rect 14568 14940 14596 16186
rect 14660 16114 14688 17546
rect 15028 17338 15056 17682
rect 15396 17610 15424 18566
rect 16592 18290 16620 18702
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14936 16590 14964 16934
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14646 15464 14702 15473
rect 14646 15399 14702 15408
rect 14660 15162 14688 15399
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14516 14912 14596 14940
rect 14464 14894 14516 14900
rect 14476 14822 14504 14894
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14462 14240 14518 14249
rect 14462 14175 14518 14184
rect 14476 13938 14504 14175
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13326 14504 13670
rect 14568 13326 14596 13738
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14556 13320 14608 13326
rect 14752 13308 14780 15302
rect 14936 15026 14964 16526
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 15978 15332 16390
rect 15396 16182 15424 16526
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 15488 16046 15516 18226
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 15586 15240 15846
rect 15120 15570 15240 15586
rect 15108 15564 15240 15570
rect 15160 15558 15240 15564
rect 15108 15506 15160 15512
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14830 14920 14886 14929
rect 14830 14855 14886 14864
rect 14844 14550 14872 14855
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14936 13870 14964 14962
rect 15014 14376 15070 14385
rect 15014 14311 15016 14320
rect 15068 14311 15070 14320
rect 15016 14282 15068 14288
rect 15028 13870 15056 14282
rect 15212 13920 15240 15558
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15396 14618 15424 15370
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15382 14240 15438 14249
rect 15382 14175 15438 14184
rect 15292 13932 15344 13938
rect 15212 13892 15292 13920
rect 15292 13874 15344 13880
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14752 13280 14872 13308
rect 14556 13262 14608 13268
rect 14476 12850 14504 13262
rect 14844 12986 14872 13280
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14844 12889 14872 12922
rect 14830 12880 14886 12889
rect 14568 12850 14780 12866
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14568 12844 14792 12850
rect 14568 12838 14740 12844
rect 14568 12646 14596 12838
rect 14830 12815 14886 12824
rect 14740 12786 14792 12792
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14660 12238 14688 12582
rect 14738 12336 14794 12345
rect 14738 12271 14794 12280
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14554 11792 14610 11801
rect 14554 11727 14610 11736
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14476 10724 14504 11290
rect 14384 10696 14504 10724
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14200 8634 14228 8910
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14292 8498 14320 9318
rect 14384 8974 14412 10696
rect 14568 10674 14596 11727
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14660 10810 14688 11018
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14556 10668 14608 10674
rect 14476 10628 14556 10656
rect 14476 10033 14504 10628
rect 14556 10610 14608 10616
rect 14462 10024 14518 10033
rect 14462 9959 14518 9968
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14372 8424 14424 8430
rect 14370 8392 14372 8401
rect 14424 8392 14426 8401
rect 14370 8327 14426 8336
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14384 7546 14412 7754
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14384 6866 14412 7482
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14094 6080 14150 6089
rect 14094 6015 14150 6024
rect 14108 5914 14136 6015
rect 14476 5914 14504 9959
rect 14752 9194 14780 12271
rect 14844 11694 14872 12718
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 12374 14964 12582
rect 14924 12368 14976 12374
rect 14924 12310 14976 12316
rect 15028 12306 15056 13194
rect 15304 13190 15332 13874
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15120 12238 15148 12854
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12442 15240 12786
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 14936 12102 14964 12174
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 15120 11626 15148 12174
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11830 15240 12038
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 14830 11520 14886 11529
rect 14830 11455 14886 11464
rect 14844 11150 14872 11455
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15016 10736 15068 10742
rect 15014 10704 15016 10713
rect 15068 10704 15070 10713
rect 15014 10639 15070 10648
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15212 10418 15240 10746
rect 15304 10656 15332 13126
rect 15396 12782 15424 14175
rect 15488 13938 15516 15982
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 14890 15608 15846
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15580 13802 15608 14826
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15488 12374 15516 12718
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15396 11150 15424 12174
rect 15580 11898 15608 13738
rect 15672 13462 15700 15506
rect 15856 15502 15884 16594
rect 15948 16114 15976 17478
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15948 15706 15976 15914
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15396 10810 15424 11086
rect 15580 11082 15608 11834
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15304 10628 15516 10656
rect 15384 10532 15436 10538
rect 15384 10474 15436 10480
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14660 9166 14872 9194
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14568 8362 14596 8910
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14554 7984 14610 7993
rect 14554 7919 14610 7928
rect 14568 7274 14596 7919
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14568 5778 14596 6598
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14200 5681 14228 5714
rect 14280 5704 14332 5710
rect 14186 5672 14242 5681
rect 14280 5646 14332 5652
rect 14372 5704 14424 5710
rect 14660 5658 14688 9166
rect 14844 8974 14872 9166
rect 14936 8974 14964 9522
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14752 8634 14780 8910
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14844 8498 14872 8774
rect 14832 8492 14884 8498
rect 14752 8452 14832 8480
rect 14752 7750 14780 8452
rect 14832 8434 14884 8440
rect 15028 7954 15056 10406
rect 15120 8634 15148 10406
rect 15212 10390 15332 10418
rect 15304 10266 15332 10390
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15200 10192 15252 10198
rect 15198 10160 15200 10169
rect 15252 10160 15254 10169
rect 15396 10146 15424 10474
rect 15198 10095 15254 10104
rect 15304 10118 15424 10146
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14844 7546 14872 7822
rect 14936 7721 14964 7822
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 14922 7712 14978 7721
rect 14922 7647 14978 7656
rect 15028 7585 15056 7754
rect 15014 7576 15070 7585
rect 14832 7540 14884 7546
rect 15212 7546 15240 8502
rect 15014 7511 15070 7520
rect 15200 7540 15252 7546
rect 14832 7482 14884 7488
rect 15200 7482 15252 7488
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 14372 5646 14424 5652
rect 14186 5607 14242 5616
rect 14200 5234 14228 5607
rect 14292 5370 14320 5646
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14384 5234 14412 5646
rect 14476 5630 14688 5658
rect 14476 5234 14504 5630
rect 14752 5370 14780 7210
rect 15212 6934 15240 7482
rect 15304 7410 15332 10118
rect 15488 9330 15516 10628
rect 15580 10062 15608 11018
rect 15672 11014 15700 13398
rect 15856 13190 15884 15438
rect 16040 15026 16068 18226
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16224 17746 16252 18090
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16408 17338 16436 18226
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16224 14074 16252 15370
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12434 15884 13126
rect 15856 12406 16068 12434
rect 16040 12238 16068 12406
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15856 11898 15884 12106
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15948 11830 15976 12174
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 15844 11688 15896 11694
rect 15936 11688 15988 11694
rect 15844 11630 15896 11636
rect 15934 11656 15936 11665
rect 15988 11656 15990 11665
rect 15856 11354 15884 11630
rect 15934 11591 15990 11600
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 16040 11218 16068 12174
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 11393 16160 11698
rect 16118 11384 16174 11393
rect 16118 11319 16174 11328
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 16316 11150 16344 17070
rect 16500 14618 16528 17138
rect 16592 16674 16620 18226
rect 16684 17202 16712 18634
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17610 16804 18022
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 17202 17724 17478
rect 16672 17196 16724 17202
rect 17684 17196 17736 17202
rect 16724 17156 16804 17184
rect 16672 17138 16724 17144
rect 16776 16794 16804 17156
rect 17684 17138 17736 17144
rect 17696 17105 17724 17138
rect 17682 17096 17738 17105
rect 17682 17031 17738 17040
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16592 16658 16804 16674
rect 16592 16652 16816 16658
rect 16592 16646 16764 16652
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16120 11144 16172 11150
rect 15948 11092 16120 11098
rect 15948 11086 16172 11092
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 15948 11070 16160 11086
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15672 10130 15700 10950
rect 15752 10668 15804 10674
rect 15804 10628 15884 10656
rect 15752 10610 15804 10616
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15396 9302 15792 9330
rect 15396 8378 15424 9302
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15474 9072 15530 9081
rect 15474 9007 15530 9016
rect 15488 8974 15516 9007
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15580 8498 15608 9114
rect 15764 8974 15792 9302
rect 15856 9217 15884 10628
rect 15842 9208 15898 9217
rect 15842 9143 15898 9152
rect 15856 8974 15884 9143
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15672 8634 15700 8910
rect 15948 8634 15976 11070
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16224 10674 16252 10950
rect 16408 10742 16436 13942
rect 16500 13326 16528 14554
rect 16592 14498 16620 16646
rect 16764 16594 16816 16600
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16672 15904 16724 15910
rect 16670 15872 16672 15881
rect 16724 15872 16726 15881
rect 16670 15807 16726 15816
rect 16776 14958 16804 16118
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 15570 16896 15846
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16868 15162 16896 15506
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16960 15026 16988 15982
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16684 14793 16712 14826
rect 16670 14784 16726 14793
rect 16670 14719 16726 14728
rect 16592 14482 16712 14498
rect 16580 14476 16712 14482
rect 16632 14470 16712 14476
rect 16580 14418 16632 14424
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16592 11370 16620 14282
rect 16684 12850 16712 14470
rect 16776 13938 16804 14894
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16776 12986 16804 13874
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16868 12850 16896 13806
rect 16960 13394 16988 14962
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16684 12306 16712 12786
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16776 12170 16804 12582
rect 16960 12434 16988 13330
rect 17696 12918 17724 15302
rect 17880 14618 17908 15370
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 18050 14376 18106 14385
rect 17788 14074 17816 14350
rect 17960 14340 18012 14346
rect 18050 14311 18106 14320
rect 17960 14282 18012 14288
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17972 13705 18000 14282
rect 18064 14006 18092 14311
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 17958 13696 18014 13705
rect 17958 13631 18014 13640
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17328 12753 17356 12786
rect 17314 12744 17370 12753
rect 17314 12679 17370 12688
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 16868 12406 16988 12434
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16868 11558 16896 12406
rect 18064 12345 18092 12582
rect 18050 12336 18106 12345
rect 18050 12271 18106 12280
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17788 11762 17816 12038
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16500 11354 16620 11370
rect 16488 11348 16620 11354
rect 16540 11342 16620 11348
rect 16488 11290 16540 11296
rect 16578 11248 16634 11257
rect 16578 11183 16634 11192
rect 16592 10810 16620 11183
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16304 10736 16356 10742
rect 16304 10678 16356 10684
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16132 10198 16160 10610
rect 16224 10470 16252 10610
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 16120 9988 16172 9994
rect 16120 9930 16172 9936
rect 16040 9450 16068 9930
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15396 8350 15608 8378
rect 15384 8288 15436 8294
rect 15382 8256 15384 8265
rect 15436 8256 15438 8265
rect 15382 8191 15438 8200
rect 15396 8022 15424 8191
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7546 15424 7686
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15304 7313 15332 7346
rect 15290 7304 15346 7313
rect 15580 7274 15608 8350
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15290 7239 15346 7248
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15200 6928 15252 6934
rect 14922 6896 14978 6905
rect 15200 6870 15252 6876
rect 14922 6831 14978 6840
rect 15016 6860 15068 6866
rect 14936 6798 14964 6831
rect 15016 6802 15068 6808
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 15028 5273 15056 6802
rect 15476 6792 15528 6798
rect 15580 6780 15608 7210
rect 15528 6752 15608 6780
rect 15476 6734 15528 6740
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15120 6458 15148 6666
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15120 5574 15148 5646
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5302 15240 5510
rect 15200 5296 15252 5302
rect 15014 5264 15070 5273
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14556 5228 14608 5234
rect 15200 5238 15252 5244
rect 15014 5199 15016 5208
rect 14556 5170 14608 5176
rect 15068 5199 15070 5208
rect 15016 5170 15068 5176
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 14384 4826 14412 5170
rect 14476 4826 14504 5170
rect 14568 4865 14596 5170
rect 14554 4856 14610 4865
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14464 4820 14516 4826
rect 15212 4826 15240 5238
rect 15304 5234 15332 5782
rect 15488 5234 15516 5850
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 15580 5370 15608 5578
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 14554 4791 14610 4800
rect 15200 4820 15252 4826
rect 14464 4762 14516 4768
rect 15200 4762 15252 4768
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13004 4146 13032 4490
rect 13832 4282 13860 4558
rect 14476 4486 14504 4762
rect 15198 4720 15254 4729
rect 15198 4655 15254 4664
rect 15212 4486 15240 4655
rect 15304 4622 15332 4966
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13832 4162 13860 4218
rect 13832 4146 13952 4162
rect 14476 4146 14504 4422
rect 14568 4282 14596 4422
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13084 4140 13136 4146
rect 13832 4140 13964 4146
rect 13832 4134 13912 4140
rect 13084 4082 13136 4088
rect 13912 4082 13964 4088
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 13096 4026 13124 4082
rect 12912 4010 13124 4026
rect 14280 4072 14332 4078
rect 14568 4026 14596 4218
rect 15212 4214 15240 4422
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 14332 4020 14596 4026
rect 14280 4014 14596 4020
rect 12900 4004 13124 4010
rect 12952 3998 13124 4004
rect 14292 3998 14596 4014
rect 15396 4010 15424 5102
rect 15672 4826 15700 8298
rect 15764 6769 15792 8434
rect 16040 8430 16068 9386
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16040 7868 16068 8230
rect 16132 8022 16160 9930
rect 16224 9042 16252 10202
rect 16316 9994 16344 10678
rect 16684 10266 16712 11018
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16684 10130 16712 10202
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 16316 9178 16344 9930
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16224 8634 16252 8842
rect 16408 8809 16436 8910
rect 16394 8800 16450 8809
rect 16394 8735 16450 8744
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 16040 7840 16160 7868
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15750 6760 15806 6769
rect 15750 6695 15752 6704
rect 15804 6695 15806 6704
rect 15752 6666 15804 6672
rect 15750 6352 15806 6361
rect 15750 6287 15806 6296
rect 15764 6254 15792 6287
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15488 4622 15516 4694
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15580 4078 15608 4558
rect 15764 4554 15792 5646
rect 15856 5098 15884 7754
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15948 6798 15976 7278
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16026 6352 16082 6361
rect 16026 6287 16082 6296
rect 16040 6254 16068 6287
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16040 5914 16068 6190
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16132 5710 16160 7840
rect 16224 6322 16252 8570
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 7818 16344 8230
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16408 6798 16436 8735
rect 16500 6934 16528 9998
rect 16670 9752 16726 9761
rect 16670 9687 16726 9696
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16592 9081 16620 9114
rect 16684 9110 16712 9687
rect 16672 9104 16724 9110
rect 16578 9072 16634 9081
rect 16672 9046 16724 9052
rect 16578 9007 16634 9016
rect 16592 8922 16620 9007
rect 16592 8894 16712 8922
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16592 8498 16620 8774
rect 16684 8634 16712 8894
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16684 7954 16712 8366
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6390 16436 6598
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16486 6352 16542 6361
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16212 6180 16264 6186
rect 16316 6168 16344 6258
rect 16264 6140 16344 6168
rect 16212 6122 16264 6128
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 15948 5574 15976 5646
rect 16224 5642 16252 6122
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 15936 5568 15988 5574
rect 16224 5545 16252 5578
rect 15936 5510 15988 5516
rect 16210 5536 16266 5545
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15948 4282 15976 5510
rect 16210 5471 16266 5480
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16316 4146 16344 5714
rect 16408 4622 16436 6326
rect 16486 6287 16488 6296
rect 16540 6287 16542 6296
rect 16488 6258 16540 6264
rect 16776 5710 16804 11494
rect 16868 10606 16896 11494
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16960 10062 16988 11562
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17052 10266 17080 10610
rect 17236 10606 17264 11290
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17420 10742 17448 10950
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16856 9648 16908 9654
rect 16854 9616 16856 9625
rect 16908 9616 16910 9625
rect 16854 9551 16910 9560
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16868 9178 16896 9454
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16868 8430 16896 9114
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16856 8288 16908 8294
rect 16854 8256 16856 8265
rect 16908 8256 16910 8265
rect 16854 8191 16910 8200
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16868 6610 16896 7754
rect 16960 6798 16988 9998
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 8650 17080 9862
rect 17236 9704 17264 10542
rect 17420 10180 17448 10678
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17696 10441 17724 10610
rect 17682 10432 17738 10441
rect 17682 10367 17738 10376
rect 17420 10152 17540 10180
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17144 9676 17264 9704
rect 17144 8974 17172 9676
rect 17222 9616 17278 9625
rect 17222 9551 17278 9560
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17130 8664 17186 8673
rect 17052 8622 17130 8650
rect 17130 8599 17186 8608
rect 17144 8498 17172 8599
rect 17236 8498 17264 9551
rect 17328 9518 17356 9998
rect 17420 9586 17448 9998
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17420 9160 17448 9522
rect 17512 9518 17540 10152
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17604 9761 17632 9998
rect 17590 9752 17646 9761
rect 17590 9687 17646 9696
rect 17590 9616 17646 9625
rect 17590 9551 17646 9560
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17328 9132 17448 9160
rect 17328 8838 17356 9132
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17420 8498 17448 8978
rect 17512 8974 17540 9454
rect 17604 8974 17632 9551
rect 17788 9382 17816 11562
rect 17972 11150 18000 12038
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17868 10056 17920 10062
rect 17866 10024 17868 10033
rect 17920 10024 17922 10033
rect 17866 9959 17922 9968
rect 18064 9586 18092 10610
rect 18156 9654 18184 11154
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17684 9104 17736 9110
rect 17684 9046 17736 9052
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 16868 6582 16988 6610
rect 16854 6488 16910 6497
rect 16854 6423 16910 6432
rect 16868 6390 16896 6423
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16856 6248 16908 6254
rect 16960 6236 16988 6582
rect 17052 6458 17080 6734
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16908 6208 16988 6236
rect 16856 6190 16908 6196
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16408 4146 16436 4558
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15384 4004 15436 4010
rect 12900 3946 12952 3952
rect 15384 3946 15436 3952
rect 16776 3942 16804 5646
rect 16868 5030 16896 6190
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16960 5234 16988 5646
rect 17052 5302 17080 6394
rect 17144 5710 17172 7686
rect 17328 6322 17356 8434
rect 17512 8090 17540 8910
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17604 7750 17632 8774
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17420 6322 17448 6802
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17604 6322 17632 6598
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17328 5914 17356 6258
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17144 5574 17172 5646
rect 17696 5642 17724 9046
rect 17788 8498 17816 9318
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18064 7585 18092 7686
rect 18050 7576 18106 7585
rect 18050 7511 18106 7520
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4690 16896 4966
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16960 4622 16988 5170
rect 17052 4758 17080 5238
rect 17144 5216 17172 5510
rect 17224 5228 17276 5234
rect 17144 5188 17224 5216
rect 17224 5170 17276 5176
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16960 4146 16988 4558
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 9048 800 9076 2246
rect 11624 800 11652 2246
rect 9034 0 9090 800
rect 11610 0 11666 800
<< via2 >>
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 5170 18264 5226 18320
rect 1490 16360 1546 16416
rect 1306 15700 1362 15736
rect 1306 15680 1308 15700
rect 1308 15680 1360 15700
rect 1360 15680 1362 15700
rect 846 14456 902 14512
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1306 13640 1362 13696
rect 1122 11600 1178 11656
rect 1490 9560 1546 9616
rect 2686 14864 2742 14920
rect 2686 14456 2742 14512
rect 2226 13368 2282 13424
rect 2134 9968 2190 10024
rect 1490 8200 1546 8256
rect 3054 15444 3056 15464
rect 3056 15444 3108 15464
rect 3108 15444 3110 15464
rect 3054 15408 3110 15444
rect 4066 17584 4122 17640
rect 3238 14048 3294 14104
rect 2870 12960 2926 13016
rect 3146 12844 3202 12880
rect 3146 12824 3148 12844
rect 3148 12824 3200 12844
rect 3200 12824 3202 12844
rect 2870 12280 2926 12336
rect 2594 9424 2650 9480
rect 2318 9016 2374 9072
rect 1858 7520 1914 7576
rect 846 6704 902 6760
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 3974 14492 3976 14512
rect 3976 14492 4028 14512
rect 4028 14492 4030 14512
rect 3974 14456 4030 14492
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 3974 14320 4030 14376
rect 3882 13932 3938 13968
rect 3882 13912 3884 13932
rect 3884 13912 3936 13932
rect 3936 13912 3938 13932
rect 3882 12280 3938 12336
rect 3790 12144 3846 12200
rect 3698 10668 3754 10704
rect 3698 10648 3700 10668
rect 3700 10648 3752 10668
rect 3752 10648 3754 10668
rect 3606 9596 3608 9616
rect 3608 9596 3660 9616
rect 3660 9596 3662 9616
rect 3606 9560 3662 9596
rect 3422 7792 3478 7848
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 5354 17040 5410 17096
rect 4894 16516 4950 16552
rect 4894 16496 4896 16516
rect 4896 16496 4948 16516
rect 4948 16496 4950 16516
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4710 15700 4766 15736
rect 4710 15680 4712 15700
rect 4712 15680 4764 15700
rect 4764 15680 4766 15700
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 5722 16360 5778 16416
rect 5630 15952 5686 16008
rect 5538 15544 5594 15600
rect 5170 14728 5226 14784
rect 5262 14592 5318 14648
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4250 12280 4306 12336
rect 4158 11756 4214 11792
rect 4158 11736 4160 11756
rect 4160 11736 4212 11756
rect 4212 11736 4214 11756
rect 4526 12008 4582 12064
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4250 11600 4306 11656
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 5170 11600 5226 11656
rect 4986 11076 5042 11112
rect 4986 11056 4988 11076
rect 4988 11056 5040 11076
rect 5040 11056 5042 11076
rect 3974 10512 4030 10568
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4342 10104 4398 10160
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3882 8472 3938 8528
rect 4342 8916 4344 8936
rect 4344 8916 4396 8936
rect 4396 8916 4398 8936
rect 4342 8880 4398 8916
rect 3330 4664 3386 4720
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4986 10240 5042 10296
rect 4802 10104 4858 10160
rect 5446 11736 5502 11792
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5170 9324 5172 9344
rect 5172 9324 5224 9344
rect 5224 9324 5226 9344
rect 5170 9288 5226 9324
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4618 8472 4674 8528
rect 4618 8234 4674 8290
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4342 7928 4398 7984
rect 4894 8200 4950 8256
rect 4986 8084 5042 8120
rect 4986 8064 4988 8084
rect 4988 8064 5040 8084
rect 5040 8064 5042 8084
rect 5262 8336 5318 8392
rect 5538 10784 5594 10840
rect 7102 17040 7158 17096
rect 7286 17448 7342 17504
rect 7562 17176 7618 17232
rect 6182 14048 6238 14104
rect 6550 15580 6552 15600
rect 6552 15580 6604 15600
rect 6604 15580 6606 15600
rect 6550 15544 6606 15580
rect 6734 15544 6790 15600
rect 6090 13912 6146 13968
rect 6090 13640 6146 13696
rect 6090 12588 6092 12608
rect 6092 12588 6144 12608
rect 6144 12588 6146 12608
rect 6090 12552 6146 12588
rect 5814 10376 5870 10432
rect 5722 8608 5778 8664
rect 5630 7928 5686 7984
rect 4066 7248 4122 7304
rect 4710 7384 4766 7440
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 5078 7404 5134 7440
rect 5078 7384 5080 7404
rect 5080 7384 5132 7404
rect 5132 7384 5134 7404
rect 5538 7656 5594 7712
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4342 6740 4344 6760
rect 4344 6740 4396 6760
rect 4396 6740 4398 6760
rect 4066 6432 4122 6488
rect 4342 6704 4398 6740
rect 4710 6296 4766 6352
rect 4710 6160 4766 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5170 7248 5226 7304
rect 5262 6840 5318 6896
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 5262 6296 5318 6352
rect 5998 11600 6054 11656
rect 5906 9324 5908 9344
rect 5908 9324 5960 9344
rect 5960 9324 5962 9344
rect 5906 9288 5962 9324
rect 6366 13776 6422 13832
rect 6550 12552 6606 12608
rect 6550 12416 6606 12472
rect 6366 12144 6422 12200
rect 6366 11872 6422 11928
rect 6274 11328 6330 11384
rect 6366 11192 6422 11248
rect 6182 10512 6238 10568
rect 7286 16224 7342 16280
rect 7194 15680 7250 15736
rect 7654 16496 7710 16552
rect 7470 16088 7526 16144
rect 9586 18264 9642 18320
rect 6734 11056 6790 11112
rect 6734 9968 6790 10024
rect 6734 9832 6790 9888
rect 6642 9696 6698 9752
rect 6550 9152 6606 9208
rect 5630 6976 5686 7032
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 5446 5344 5502 5400
rect 6090 8744 6146 8800
rect 6182 8472 6238 8528
rect 6274 7948 6330 7984
rect 6274 7928 6276 7948
rect 6276 7928 6328 7948
rect 6328 7928 6330 7948
rect 6366 7792 6422 7848
rect 6274 7520 6330 7576
rect 5906 6452 5962 6488
rect 5906 6432 5908 6452
rect 5908 6432 5960 6452
rect 5960 6432 5962 6452
rect 6642 8880 6698 8936
rect 6366 6160 6422 6216
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 6458 4664 6514 4720
rect 6274 4564 6276 4584
rect 6276 4564 6328 4584
rect 6328 4564 6330 4584
rect 6274 4528 6330 4564
rect 7378 12280 7434 12336
rect 7562 12416 7618 12472
rect 7194 9832 7250 9888
rect 7378 10920 7434 10976
rect 7562 11464 7618 11520
rect 7470 10240 7526 10296
rect 6826 8064 6882 8120
rect 7010 8064 7066 8120
rect 7286 9460 7288 9480
rect 7288 9460 7340 9480
rect 7340 9460 7342 9480
rect 7286 9424 7342 9460
rect 7194 8064 7250 8120
rect 7010 7248 7066 7304
rect 6826 6840 6882 6896
rect 7010 6432 7066 6488
rect 6826 5344 6882 5400
rect 7194 7520 7250 7576
rect 7930 11192 7986 11248
rect 7930 9288 7986 9344
rect 8390 15444 8392 15464
rect 8392 15444 8444 15464
rect 8444 15444 8446 15464
rect 8390 15408 8446 15444
rect 8482 13368 8538 13424
rect 8298 13268 8300 13288
rect 8300 13268 8352 13288
rect 8352 13268 8354 13288
rect 8298 13232 8354 13268
rect 8482 13268 8484 13288
rect 8484 13268 8536 13288
rect 8536 13268 8538 13288
rect 8482 13232 8538 13268
rect 8206 12688 8262 12744
rect 8206 10512 8262 10568
rect 8114 9968 8170 10024
rect 7746 8608 7802 8664
rect 7746 8492 7802 8528
rect 7746 8472 7748 8492
rect 7748 8472 7800 8492
rect 7800 8472 7802 8492
rect 7838 8336 7894 8392
rect 7654 7928 7710 7984
rect 7378 5228 7434 5264
rect 7378 5208 7380 5228
rect 7380 5208 7432 5228
rect 7432 5208 7434 5228
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 7930 8200 7986 8256
rect 7838 6296 7894 6352
rect 8574 9988 8630 10024
rect 8574 9968 8576 9988
rect 8576 9968 8628 9988
rect 8628 9968 8630 9988
rect 8390 8356 8446 8392
rect 8390 8336 8392 8356
rect 8392 8336 8444 8356
rect 8444 8336 8446 8356
rect 8114 8200 8170 8256
rect 8114 7656 8170 7712
rect 8206 7384 8262 7440
rect 8390 7248 8446 7304
rect 8114 6976 8170 7032
rect 8298 6976 8354 7032
rect 8206 6432 8262 6488
rect 8850 17484 8852 17504
rect 8852 17484 8904 17504
rect 8904 17484 8906 17504
rect 8850 17448 8906 17484
rect 9126 17176 9182 17232
rect 9770 17196 9826 17232
rect 9770 17176 9772 17196
rect 9772 17176 9824 17196
rect 9824 17176 9826 17196
rect 9218 16768 9274 16824
rect 8850 16632 8906 16688
rect 8850 15272 8906 15328
rect 8850 15136 8906 15192
rect 8758 14456 8814 14512
rect 8758 14048 8814 14104
rect 8850 13640 8906 13696
rect 9034 14340 9090 14376
rect 9034 14320 9036 14340
rect 9036 14320 9088 14340
rect 9088 14320 9090 14340
rect 9310 15952 9366 16008
rect 9494 16532 9496 16552
rect 9496 16532 9548 16552
rect 9548 16532 9550 16552
rect 9494 16496 9550 16532
rect 9126 14220 9128 14240
rect 9128 14220 9180 14240
rect 9180 14220 9182 14240
rect 9126 14184 9182 14220
rect 9218 13388 9274 13424
rect 9218 13368 9220 13388
rect 9220 13368 9272 13388
rect 9272 13368 9274 13388
rect 9034 12552 9090 12608
rect 8942 12416 8998 12472
rect 9218 12688 9274 12744
rect 9218 12552 9274 12608
rect 8850 12164 8906 12200
rect 8850 12144 8852 12164
rect 8852 12144 8904 12164
rect 8904 12144 8906 12164
rect 8942 12008 8998 12064
rect 9034 11736 9090 11792
rect 8850 10784 8906 10840
rect 8850 10512 8906 10568
rect 8850 10104 8906 10160
rect 9218 11464 9274 11520
rect 9126 11328 9182 11384
rect 9494 14728 9550 14784
rect 9402 14456 9458 14512
rect 9678 14864 9734 14920
rect 9586 13268 9588 13288
rect 9588 13268 9640 13288
rect 9640 13268 9642 13288
rect 9586 13232 9642 13268
rect 10230 17620 10232 17640
rect 10232 17620 10284 17640
rect 10284 17620 10286 17640
rect 10230 17584 10286 17620
rect 10322 16124 10324 16144
rect 10324 16124 10376 16144
rect 10376 16124 10378 16144
rect 10322 16088 10378 16124
rect 10506 15952 10562 16008
rect 9862 13932 9918 13968
rect 9862 13912 9864 13932
rect 9864 13912 9916 13932
rect 9916 13912 9918 13932
rect 9770 13368 9826 13424
rect 9586 12552 9642 12608
rect 9402 11600 9458 11656
rect 8942 9560 8998 9616
rect 9034 8744 9090 8800
rect 8942 8608 8998 8664
rect 9034 8200 9090 8256
rect 8850 7656 8906 7712
rect 8942 7384 8998 7440
rect 9402 10260 9458 10296
rect 9402 10240 9404 10260
rect 9404 10240 9456 10260
rect 9456 10240 9458 10260
rect 9678 11092 9680 11112
rect 9680 11092 9732 11112
rect 9732 11092 9734 11112
rect 9678 11056 9734 11092
rect 10322 15136 10378 15192
rect 10506 14456 10562 14512
rect 10322 13776 10378 13832
rect 9862 11464 9918 11520
rect 9310 8744 9366 8800
rect 9126 7384 9182 7440
rect 8850 7112 8906 7168
rect 9034 7148 9036 7168
rect 9036 7148 9088 7168
rect 9088 7148 9090 7168
rect 9034 7112 9090 7148
rect 8942 6332 8944 6352
rect 8944 6332 8996 6352
rect 8996 6332 8998 6352
rect 8942 6296 8998 6332
rect 9034 6160 9090 6216
rect 8574 4528 8630 4584
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9586 8084 9642 8120
rect 9586 8064 9588 8084
rect 9588 8064 9640 8084
rect 9640 8064 9642 8084
rect 9586 7928 9642 7984
rect 9862 9988 9918 10024
rect 9862 9968 9864 9988
rect 9864 9968 9916 9988
rect 9916 9968 9918 9988
rect 10138 11212 10194 11248
rect 10138 11192 10140 11212
rect 10140 11192 10192 11212
rect 10192 11192 10194 11212
rect 10414 13232 10470 13288
rect 10230 10376 10286 10432
rect 10138 10104 10194 10160
rect 9954 8780 9956 8800
rect 9956 8780 10008 8800
rect 10008 8780 10010 8800
rect 9954 8744 10010 8780
rect 9862 8628 9918 8664
rect 9862 8608 9864 8628
rect 9864 8608 9916 8628
rect 9916 8608 9918 8628
rect 9862 8492 9918 8528
rect 9862 8472 9864 8492
rect 9864 8472 9916 8492
rect 9916 8472 9918 8492
rect 9402 5344 9458 5400
rect 10322 9868 10324 9888
rect 10324 9868 10376 9888
rect 10376 9868 10378 9888
rect 10322 9832 10378 9868
rect 11242 17620 11244 17640
rect 11244 17620 11296 17640
rect 11296 17620 11298 17640
rect 11242 17584 11298 17620
rect 10874 16632 10930 16688
rect 10690 16088 10746 16144
rect 10874 15444 10876 15464
rect 10876 15444 10928 15464
rect 10928 15444 10930 15464
rect 10874 15408 10930 15444
rect 10506 11192 10562 11248
rect 10598 11092 10600 11112
rect 10600 11092 10652 11112
rect 10652 11092 10654 11112
rect 10598 11056 10654 11092
rect 10598 10920 10654 10976
rect 10506 9696 10562 9752
rect 10230 9288 10286 9344
rect 9954 6432 10010 6488
rect 10322 8880 10378 8936
rect 10874 10104 10930 10160
rect 10690 9968 10746 10024
rect 12070 17196 12126 17232
rect 12070 17176 12072 17196
rect 12072 17176 12124 17196
rect 12124 17176 12126 17196
rect 11702 17040 11758 17096
rect 11886 15816 11942 15872
rect 11150 13096 11206 13152
rect 11150 12416 11206 12472
rect 11426 14220 11428 14240
rect 11428 14220 11480 14240
rect 11480 14220 11482 14240
rect 11426 14184 11482 14220
rect 11334 13232 11390 13288
rect 11242 12144 11298 12200
rect 11150 11872 11206 11928
rect 10322 8336 10378 8392
rect 10414 7928 10470 7984
rect 10690 8200 10746 8256
rect 10138 6332 10140 6352
rect 10140 6332 10192 6352
rect 10192 6332 10194 6352
rect 10138 6296 10194 6332
rect 10414 6296 10470 6352
rect 10598 6704 10654 6760
rect 10322 5772 10378 5808
rect 10322 5752 10324 5772
rect 10324 5752 10376 5772
rect 10376 5752 10378 5772
rect 10138 5480 10194 5536
rect 10046 5344 10102 5400
rect 10138 4800 10194 4856
rect 11058 9424 11114 9480
rect 11058 9172 11114 9208
rect 11058 9152 11060 9172
rect 11060 9152 11112 9172
rect 11112 9152 11114 9172
rect 11058 8608 11114 8664
rect 11150 8336 11206 8392
rect 11058 7928 11114 7984
rect 11058 6840 11114 6896
rect 11334 11464 11390 11520
rect 11518 9324 11520 9344
rect 11520 9324 11572 9344
rect 11572 9324 11574 9344
rect 11518 9288 11574 9324
rect 11610 8608 11666 8664
rect 10966 5752 11022 5808
rect 10874 5344 10930 5400
rect 12070 16124 12072 16144
rect 12072 16124 12124 16144
rect 12124 16124 12126 16144
rect 12070 16088 12126 16124
rect 12346 16360 12402 16416
rect 12254 15816 12310 15872
rect 12254 14592 12310 14648
rect 12254 14048 12310 14104
rect 12346 13812 12348 13832
rect 12348 13812 12400 13832
rect 12400 13812 12402 13832
rect 12346 13776 12402 13812
rect 12622 13932 12678 13968
rect 12622 13912 12624 13932
rect 12624 13912 12676 13932
rect 12676 13912 12678 13932
rect 13174 16532 13176 16552
rect 13176 16532 13228 16552
rect 13228 16532 13230 16552
rect 13174 16496 13230 16532
rect 13174 16224 13230 16280
rect 13082 15272 13138 15328
rect 12898 14068 12954 14104
rect 12898 14048 12900 14068
rect 12900 14048 12952 14068
rect 12952 14048 12954 14068
rect 12254 12416 12310 12472
rect 11978 12280 12034 12336
rect 11886 12164 11942 12200
rect 11886 12144 11888 12164
rect 11888 12144 11940 12164
rect 11940 12144 11942 12164
rect 11886 11872 11942 11928
rect 12162 12316 12164 12336
rect 12164 12316 12216 12336
rect 12216 12316 12218 12336
rect 12162 12280 12218 12316
rect 11702 7948 11758 7984
rect 11702 7928 11704 7948
rect 11704 7928 11756 7948
rect 11756 7928 11758 7948
rect 11978 9424 12034 9480
rect 11886 8336 11942 8392
rect 12254 9152 12310 9208
rect 12254 8744 12310 8800
rect 12530 11600 12586 11656
rect 12346 7384 12402 7440
rect 11518 6160 11574 6216
rect 10598 4664 10654 4720
rect 11518 4800 11574 4856
rect 10506 3984 10562 4040
rect 10506 3884 10508 3904
rect 10508 3884 10560 3904
rect 10560 3884 10562 3904
rect 10506 3848 10562 3884
rect 12346 6160 12402 6216
rect 13082 12416 13138 12472
rect 14002 15952 14058 16008
rect 13726 15544 13782 15600
rect 13910 15544 13966 15600
rect 12990 12164 13046 12200
rect 12990 12144 12992 12164
rect 12992 12144 13044 12164
rect 13044 12144 13046 12164
rect 12898 11872 12954 11928
rect 13450 11872 13506 11928
rect 13082 11600 13138 11656
rect 13266 11600 13322 11656
rect 13174 9696 13230 9752
rect 12898 8880 12954 8936
rect 13174 9424 13230 9480
rect 12714 7384 12770 7440
rect 12806 7112 12862 7168
rect 12714 6976 12770 7032
rect 13542 11464 13598 11520
rect 14278 16360 14334 16416
rect 13910 13796 13966 13832
rect 13910 13776 13912 13796
rect 13912 13776 13964 13796
rect 13964 13776 13966 13796
rect 14278 13776 14334 13832
rect 13634 9424 13690 9480
rect 13542 9288 13598 9344
rect 13542 9152 13598 9208
rect 13266 7384 13322 7440
rect 13542 7812 13598 7848
rect 13542 7792 13544 7812
rect 13544 7792 13596 7812
rect 13596 7792 13598 7812
rect 13266 6432 13322 6488
rect 14094 9832 14150 9888
rect 13726 6196 13728 6216
rect 13728 6196 13780 6216
rect 13780 6196 13782 6216
rect 13358 5752 13414 5808
rect 12438 4700 12440 4720
rect 12440 4700 12492 4720
rect 12492 4700 12494 4720
rect 12438 4664 12494 4700
rect 13726 6160 13782 6196
rect 14002 7520 14058 7576
rect 13910 5480 13966 5536
rect 14646 15408 14702 15464
rect 14462 14184 14518 14240
rect 14830 14864 14886 14920
rect 15014 14340 15070 14376
rect 15014 14320 15016 14340
rect 15016 14320 15068 14340
rect 15068 14320 15070 14340
rect 15382 14184 15438 14240
rect 14830 12824 14886 12880
rect 14738 12280 14794 12336
rect 14554 11736 14610 11792
rect 14462 9968 14518 10024
rect 14370 8372 14372 8392
rect 14372 8372 14424 8392
rect 14424 8372 14426 8392
rect 14370 8336 14426 8372
rect 14094 6024 14150 6080
rect 14830 11464 14886 11520
rect 15014 10684 15016 10704
rect 15016 10684 15068 10704
rect 15068 10684 15070 10704
rect 15014 10648 15070 10684
rect 14554 7928 14610 7984
rect 14186 5616 14242 5672
rect 15198 10140 15200 10160
rect 15200 10140 15252 10160
rect 15252 10140 15254 10160
rect 15198 10104 15254 10140
rect 14922 7656 14978 7712
rect 15014 7520 15070 7576
rect 15934 11636 15936 11656
rect 15936 11636 15988 11656
rect 15988 11636 15990 11656
rect 15934 11600 15990 11636
rect 16118 11328 16174 11384
rect 17682 17040 17738 17096
rect 15474 9016 15530 9072
rect 15842 9152 15898 9208
rect 16670 15852 16672 15872
rect 16672 15852 16724 15872
rect 16724 15852 16726 15872
rect 16670 15816 16726 15852
rect 16670 14728 16726 14784
rect 18050 14320 18106 14376
rect 17958 13640 18014 13696
rect 17314 12688 17370 12744
rect 18050 12280 18106 12336
rect 16578 11192 16634 11248
rect 15382 8236 15384 8256
rect 15384 8236 15436 8256
rect 15436 8236 15438 8256
rect 15382 8200 15438 8236
rect 15290 7248 15346 7304
rect 14922 6840 14978 6896
rect 15014 5228 15070 5264
rect 15014 5208 15016 5228
rect 15016 5208 15068 5228
rect 15068 5208 15070 5228
rect 14554 4800 14610 4856
rect 15198 4664 15254 4720
rect 16394 8744 16450 8800
rect 15750 6724 15806 6760
rect 15750 6704 15752 6724
rect 15752 6704 15804 6724
rect 15804 6704 15806 6724
rect 15750 6296 15806 6352
rect 16026 6296 16082 6352
rect 16670 9696 16726 9752
rect 16578 9016 16634 9072
rect 16210 5480 16266 5536
rect 16486 6316 16542 6352
rect 16486 6296 16488 6316
rect 16488 6296 16540 6316
rect 16540 6296 16542 6316
rect 16854 9596 16856 9616
rect 16856 9596 16908 9616
rect 16908 9596 16910 9616
rect 16854 9560 16910 9596
rect 16854 8236 16856 8256
rect 16856 8236 16908 8256
rect 16908 8236 16910 8256
rect 16854 8200 16910 8236
rect 17682 10376 17738 10432
rect 17222 9560 17278 9616
rect 17130 8608 17186 8664
rect 17590 9696 17646 9752
rect 17590 9560 17646 9616
rect 17866 10004 17868 10024
rect 17868 10004 17920 10024
rect 17920 10004 17922 10024
rect 17866 9968 17922 10004
rect 16854 6432 16910 6488
rect 18050 7520 18106 7576
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 5165 18322 5231 18325
rect 8334 18322 8340 18324
rect 5165 18320 8340 18322
rect 5165 18264 5170 18320
rect 5226 18264 8340 18320
rect 5165 18262 8340 18264
rect 5165 18259 5231 18262
rect 8334 18260 8340 18262
rect 8404 18322 8410 18324
rect 9581 18322 9647 18325
rect 8404 18320 9647 18322
rect 8404 18264 9586 18320
rect 9642 18264 9647 18320
rect 8404 18262 9647 18264
rect 8404 18260 8410 18262
rect 9581 18259 9647 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 4061 17642 4127 17645
rect 8886 17642 8892 17644
rect 4061 17640 8892 17642
rect 4061 17584 4066 17640
rect 4122 17584 8892 17640
rect 4061 17582 8892 17584
rect 4061 17579 4127 17582
rect 8886 17580 8892 17582
rect 8956 17642 8962 17644
rect 10225 17642 10291 17645
rect 8956 17640 10291 17642
rect 8956 17584 10230 17640
rect 10286 17584 10291 17640
rect 8956 17582 10291 17584
rect 8956 17580 8962 17582
rect 10225 17579 10291 17582
rect 10358 17580 10364 17644
rect 10428 17642 10434 17644
rect 11237 17642 11303 17645
rect 10428 17640 11303 17642
rect 10428 17584 11242 17640
rect 11298 17584 11303 17640
rect 10428 17582 11303 17584
rect 10428 17580 10434 17582
rect 7281 17506 7347 17509
rect 8845 17506 8911 17509
rect 10366 17506 10426 17580
rect 11237 17579 11303 17582
rect 7281 17504 10426 17506
rect 7281 17448 7286 17504
rect 7342 17448 8850 17504
rect 8906 17448 10426 17504
rect 7281 17446 10426 17448
rect 7281 17443 7347 17446
rect 8845 17443 8911 17446
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 7557 17234 7623 17237
rect 9121 17234 9187 17237
rect 7557 17232 9187 17234
rect 7557 17176 7562 17232
rect 7618 17176 9126 17232
rect 9182 17176 9187 17232
rect 7557 17174 9187 17176
rect 7557 17171 7623 17174
rect 9121 17171 9187 17174
rect 9765 17234 9831 17237
rect 12065 17234 12131 17237
rect 9765 17232 12131 17234
rect 9765 17176 9770 17232
rect 9826 17176 12070 17232
rect 12126 17176 12131 17232
rect 9765 17174 12131 17176
rect 9765 17171 9831 17174
rect 12065 17171 12131 17174
rect 5349 17098 5415 17101
rect 7097 17098 7163 17101
rect 11697 17100 11763 17101
rect 8150 17098 8156 17100
rect 5349 17096 8156 17098
rect 5349 17040 5354 17096
rect 5410 17040 7102 17096
rect 7158 17040 8156 17096
rect 5349 17038 8156 17040
rect 5349 17035 5415 17038
rect 7097 17035 7163 17038
rect 8150 17036 8156 17038
rect 8220 17036 8226 17100
rect 11646 17036 11652 17100
rect 11716 17098 11763 17100
rect 11716 17096 11808 17098
rect 11758 17040 11808 17096
rect 11716 17038 11808 17040
rect 11716 17036 11763 17038
rect 17166 17036 17172 17100
rect 17236 17098 17242 17100
rect 17677 17098 17743 17101
rect 17236 17096 17743 17098
rect 17236 17040 17682 17096
rect 17738 17040 17743 17096
rect 17236 17038 17743 17040
rect 17236 17036 17242 17038
rect 11697 17035 11763 17036
rect 17677 17035 17743 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 9070 16764 9076 16828
rect 9140 16826 9146 16828
rect 9213 16826 9279 16829
rect 9140 16824 9279 16826
rect 9140 16768 9218 16824
rect 9274 16768 9279 16824
rect 9140 16766 9279 16768
rect 9140 16764 9146 16766
rect 9213 16763 9279 16766
rect 8845 16690 8911 16693
rect 9254 16690 9260 16692
rect 8845 16688 9260 16690
rect 8845 16632 8850 16688
rect 8906 16632 9260 16688
rect 8845 16630 9260 16632
rect 8845 16627 8911 16630
rect 9254 16628 9260 16630
rect 9324 16628 9330 16692
rect 10869 16690 10935 16693
rect 11462 16690 11468 16692
rect 10869 16688 11468 16690
rect 10869 16632 10874 16688
rect 10930 16632 11468 16688
rect 10869 16630 11468 16632
rect 10869 16627 10935 16630
rect 11462 16628 11468 16630
rect 11532 16628 11538 16692
rect 4889 16554 4955 16557
rect 7649 16554 7715 16557
rect 4889 16552 7715 16554
rect 4889 16496 4894 16552
rect 4950 16496 7654 16552
rect 7710 16496 7715 16552
rect 4889 16494 7715 16496
rect 4889 16491 4955 16494
rect 7649 16491 7715 16494
rect 9489 16554 9555 16557
rect 9622 16554 9628 16556
rect 9489 16552 9628 16554
rect 9489 16496 9494 16552
rect 9550 16496 9628 16552
rect 9489 16494 9628 16496
rect 9489 16491 9555 16494
rect 9622 16492 9628 16494
rect 9692 16492 9698 16556
rect 13169 16554 13235 16557
rect 15878 16554 15884 16556
rect 13169 16552 15884 16554
rect 13169 16496 13174 16552
rect 13230 16496 15884 16552
rect 13169 16494 15884 16496
rect 13169 16491 13235 16494
rect 15878 16492 15884 16494
rect 15948 16492 15954 16556
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 5717 16420 5783 16421
rect 5717 16418 5764 16420
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 5672 16416 5764 16418
rect 5672 16360 5722 16416
rect 5672 16358 5764 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 5717 16356 5764 16358
rect 5828 16356 5834 16420
rect 12341 16418 12407 16421
rect 14273 16418 14339 16421
rect 12341 16416 14339 16418
rect 12341 16360 12346 16416
rect 12402 16360 14278 16416
rect 14334 16360 14339 16416
rect 12341 16358 14339 16360
rect 5717 16355 5783 16356
rect 12341 16355 12407 16358
rect 14273 16355 14339 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 7281 16282 7347 16285
rect 13169 16282 13235 16285
rect 7281 16280 13235 16282
rect 7281 16224 7286 16280
rect 7342 16224 13174 16280
rect 13230 16224 13235 16280
rect 7281 16222 13235 16224
rect 7281 16219 7347 16222
rect 13169 16219 13235 16222
rect 7465 16146 7531 16149
rect 9806 16146 9812 16148
rect 7465 16144 9812 16146
rect 7465 16088 7470 16144
rect 7526 16088 9812 16144
rect 7465 16086 9812 16088
rect 7465 16083 7531 16086
rect 9806 16084 9812 16086
rect 9876 16146 9882 16148
rect 10317 16146 10383 16149
rect 9876 16144 10383 16146
rect 9876 16088 10322 16144
rect 10378 16088 10383 16144
rect 9876 16086 10383 16088
rect 9876 16084 9882 16086
rect 10317 16083 10383 16086
rect 10685 16146 10751 16149
rect 12065 16146 12131 16149
rect 10685 16144 12131 16146
rect 10685 16088 10690 16144
rect 10746 16088 12070 16144
rect 12126 16088 12131 16144
rect 10685 16086 12131 16088
rect 10685 16083 10751 16086
rect 12065 16083 12131 16086
rect 3366 15948 3372 16012
rect 3436 16010 3442 16012
rect 5625 16010 5691 16013
rect 9305 16010 9371 16013
rect 3436 16008 9371 16010
rect 3436 15952 5630 16008
rect 5686 15952 9310 16008
rect 9366 15952 9371 16008
rect 3436 15950 9371 15952
rect 3436 15948 3442 15950
rect 5625 15947 5691 15950
rect 9305 15947 9371 15950
rect 10501 16010 10567 16013
rect 13997 16010 14063 16013
rect 10501 16008 14063 16010
rect 10501 15952 10506 16008
rect 10562 15952 14002 16008
rect 14058 15952 14063 16008
rect 10501 15950 14063 15952
rect 10501 15947 10567 15950
rect 13997 15947 14063 15950
rect 11881 15874 11947 15877
rect 12249 15874 12315 15877
rect 16665 15874 16731 15877
rect 16798 15874 16804 15876
rect 11881 15872 16804 15874
rect 11881 15816 11886 15872
rect 11942 15816 12254 15872
rect 12310 15816 16670 15872
rect 16726 15816 16804 15872
rect 11881 15814 16804 15816
rect 11881 15811 11947 15814
rect 12249 15811 12315 15814
rect 16665 15811 16731 15814
rect 16798 15812 16804 15814
rect 16868 15812 16874 15876
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 4705 15738 4771 15741
rect 7189 15738 7255 15741
rect 4705 15736 7255 15738
rect 4705 15680 4710 15736
rect 4766 15680 7194 15736
rect 7250 15680 7255 15736
rect 4705 15678 7255 15680
rect 4705 15675 4771 15678
rect 7189 15675 7255 15678
rect 5533 15602 5599 15605
rect 6545 15602 6611 15605
rect 5533 15600 6611 15602
rect 5533 15544 5538 15600
rect 5594 15544 6550 15600
rect 6606 15544 6611 15600
rect 5533 15542 6611 15544
rect 5533 15539 5599 15542
rect 6545 15539 6611 15542
rect 6729 15602 6795 15605
rect 13721 15602 13787 15605
rect 13905 15602 13971 15605
rect 6729 15600 13971 15602
rect 6729 15544 6734 15600
rect 6790 15544 13726 15600
rect 13782 15544 13910 15600
rect 13966 15544 13971 15600
rect 6729 15542 13971 15544
rect 6729 15539 6795 15542
rect 13721 15539 13787 15542
rect 13905 15539 13971 15542
rect 3049 15466 3115 15469
rect 8385 15466 8451 15469
rect 3049 15464 8451 15466
rect 3049 15408 3054 15464
rect 3110 15408 8390 15464
rect 8446 15408 8451 15464
rect 3049 15406 8451 15408
rect 3049 15403 3115 15406
rect 8385 15403 8451 15406
rect 10869 15466 10935 15469
rect 14641 15466 14707 15469
rect 10869 15464 14707 15466
rect 10869 15408 10874 15464
rect 10930 15408 14646 15464
rect 14702 15408 14707 15464
rect 10869 15406 14707 15408
rect 10869 15403 10935 15406
rect 14641 15403 14707 15406
rect 8845 15330 8911 15333
rect 13077 15330 13143 15333
rect 8845 15328 13143 15330
rect 8845 15272 8850 15328
rect 8906 15272 13082 15328
rect 13138 15272 13143 15328
rect 8845 15270 13143 15272
rect 8845 15267 8911 15270
rect 13077 15267 13143 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 8845 15194 8911 15197
rect 10317 15194 10383 15197
rect 8845 15192 10383 15194
rect 8845 15136 8850 15192
rect 8906 15136 10322 15192
rect 10378 15136 10383 15192
rect 8845 15134 10383 15136
rect 8845 15131 8911 15134
rect 10317 15131 10383 15134
rect 2681 14922 2747 14925
rect 2814 14922 2820 14924
rect 2681 14920 2820 14922
rect 2681 14864 2686 14920
rect 2742 14864 2820 14920
rect 2681 14862 2820 14864
rect 2681 14859 2747 14862
rect 2814 14860 2820 14862
rect 2884 14860 2890 14924
rect 9673 14922 9739 14925
rect 14825 14922 14891 14925
rect 9673 14920 14891 14922
rect 9673 14864 9678 14920
rect 9734 14864 14830 14920
rect 14886 14864 14891 14920
rect 9673 14862 14891 14864
rect 9673 14859 9739 14862
rect 14825 14859 14891 14862
rect 5165 14786 5231 14789
rect 9489 14786 9555 14789
rect 9990 14786 9996 14788
rect 5165 14784 9996 14786
rect 5165 14728 5170 14784
rect 5226 14728 9494 14784
rect 9550 14728 9996 14784
rect 5165 14726 9996 14728
rect 5165 14723 5231 14726
rect 9489 14723 9555 14726
rect 9990 14724 9996 14726
rect 10060 14724 10066 14788
rect 15878 14724 15884 14788
rect 15948 14786 15954 14788
rect 16665 14786 16731 14789
rect 15948 14784 16731 14786
rect 15948 14728 16670 14784
rect 16726 14728 16731 14784
rect 15948 14726 16731 14728
rect 15948 14724 15954 14726
rect 16665 14723 16731 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 5257 14650 5323 14653
rect 12249 14650 12315 14653
rect 5257 14648 12315 14650
rect 5257 14592 5262 14648
rect 5318 14592 12254 14648
rect 12310 14592 12315 14648
rect 5257 14590 12315 14592
rect 5257 14587 5323 14590
rect 12249 14587 12315 14590
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 2681 14514 2747 14517
rect 3969 14514 4035 14517
rect 2681 14512 4035 14514
rect 2681 14456 2686 14512
rect 2742 14456 3974 14512
rect 4030 14456 4035 14512
rect 2681 14454 4035 14456
rect 2681 14451 2747 14454
rect 3969 14451 4035 14454
rect 8753 14514 8819 14517
rect 9397 14514 9463 14517
rect 8753 14512 9463 14514
rect 8753 14456 8758 14512
rect 8814 14456 9402 14512
rect 9458 14456 9463 14512
rect 8753 14454 9463 14456
rect 8753 14451 8819 14454
rect 9397 14451 9463 14454
rect 10501 14514 10567 14517
rect 10726 14514 10732 14516
rect 10501 14512 10732 14514
rect 10501 14456 10506 14512
rect 10562 14456 10732 14512
rect 10501 14454 10732 14456
rect 10501 14451 10567 14454
rect 10726 14452 10732 14454
rect 10796 14452 10802 14516
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 3969 14378 4035 14381
rect 9029 14378 9095 14381
rect 15009 14378 15075 14381
rect 3969 14376 15075 14378
rect 3969 14320 3974 14376
rect 4030 14320 9034 14376
rect 9090 14320 15014 14376
rect 15070 14320 15075 14376
rect 3969 14318 15075 14320
rect 0 14288 800 14318
rect 3969 14315 4035 14318
rect 9029 14315 9095 14318
rect 15009 14315 15075 14318
rect 18045 14378 18111 14381
rect 18812 14378 19612 14408
rect 18045 14376 19612 14378
rect 18045 14320 18050 14376
rect 18106 14320 19612 14376
rect 18045 14318 19612 14320
rect 18045 14315 18111 14318
rect 18812 14288 19612 14318
rect 8150 14180 8156 14244
rect 8220 14242 8226 14244
rect 9121 14242 9187 14245
rect 8220 14240 9187 14242
rect 8220 14184 9126 14240
rect 9182 14184 9187 14240
rect 8220 14182 9187 14184
rect 8220 14180 8226 14182
rect 9121 14179 9187 14182
rect 11421 14242 11487 14245
rect 11646 14242 11652 14244
rect 11421 14240 11652 14242
rect 11421 14184 11426 14240
rect 11482 14184 11652 14240
rect 11421 14182 11652 14184
rect 11421 14179 11487 14182
rect 11646 14180 11652 14182
rect 11716 14242 11722 14244
rect 14457 14242 14523 14245
rect 15377 14242 15443 14245
rect 11716 14240 15443 14242
rect 11716 14184 14462 14240
rect 14518 14184 15382 14240
rect 15438 14184 15443 14240
rect 11716 14182 15443 14184
rect 11716 14180 11722 14182
rect 14457 14179 14523 14182
rect 15377 14179 15443 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 3233 14106 3299 14109
rect 3734 14106 3740 14108
rect 3233 14104 3740 14106
rect 3233 14048 3238 14104
rect 3294 14048 3740 14104
rect 3233 14046 3740 14048
rect 3233 14043 3299 14046
rect 3734 14044 3740 14046
rect 3804 14044 3810 14108
rect 6177 14106 6243 14109
rect 6177 14104 6930 14106
rect 6177 14048 6182 14104
rect 6238 14048 6930 14104
rect 6177 14046 6930 14048
rect 6177 14043 6243 14046
rect 3877 13970 3943 13973
rect 6085 13970 6151 13973
rect 3877 13968 6151 13970
rect 3877 13912 3882 13968
rect 3938 13912 6090 13968
rect 6146 13912 6151 13968
rect 3877 13910 6151 13912
rect 6870 13970 6930 14046
rect 8518 14044 8524 14108
rect 8588 14106 8594 14108
rect 8753 14106 8819 14109
rect 8588 14104 8819 14106
rect 8588 14048 8758 14104
rect 8814 14048 8819 14104
rect 8588 14046 8819 14048
rect 8588 14044 8594 14046
rect 8753 14043 8819 14046
rect 12249 14106 12315 14109
rect 12893 14106 12959 14109
rect 12249 14104 12959 14106
rect 12249 14048 12254 14104
rect 12310 14048 12898 14104
rect 12954 14048 12959 14104
rect 12249 14046 12959 14048
rect 12249 14043 12315 14046
rect 12893 14043 12959 14046
rect 9857 13970 9923 13973
rect 12617 13970 12683 13973
rect 6870 13968 12683 13970
rect 6870 13912 9862 13968
rect 9918 13912 12622 13968
rect 12678 13912 12683 13968
rect 6870 13910 12683 13912
rect 3877 13907 3943 13910
rect 6085 13907 6151 13910
rect 9857 13907 9923 13910
rect 12617 13907 12683 13910
rect 6126 13772 6132 13836
rect 6196 13834 6202 13836
rect 6361 13834 6427 13837
rect 6196 13832 6427 13834
rect 6196 13776 6366 13832
rect 6422 13776 6427 13832
rect 6196 13774 6427 13776
rect 6196 13772 6202 13774
rect 6361 13771 6427 13774
rect 10174 13772 10180 13836
rect 10244 13834 10250 13836
rect 10317 13834 10383 13837
rect 10244 13832 10383 13834
rect 10244 13776 10322 13832
rect 10378 13776 10383 13832
rect 10244 13774 10383 13776
rect 10244 13772 10250 13774
rect 10317 13771 10383 13774
rect 12341 13834 12407 13837
rect 13905 13834 13971 13837
rect 12341 13832 13971 13834
rect 12341 13776 12346 13832
rect 12402 13776 13910 13832
rect 13966 13776 13971 13832
rect 12341 13774 13971 13776
rect 12341 13771 12407 13774
rect 13905 13771 13971 13774
rect 14273 13834 14339 13837
rect 14958 13834 14964 13836
rect 14273 13832 14964 13834
rect 14273 13776 14278 13832
rect 14334 13776 14964 13832
rect 14273 13774 14964 13776
rect 14273 13771 14339 13774
rect 14958 13772 14964 13774
rect 15028 13772 15034 13836
rect 0 13698 800 13728
rect 1301 13698 1367 13701
rect 0 13696 1367 13698
rect 0 13640 1306 13696
rect 1362 13640 1367 13696
rect 0 13638 1367 13640
rect 0 13608 800 13638
rect 1301 13635 1367 13638
rect 6085 13698 6151 13701
rect 8845 13698 8911 13701
rect 6085 13696 8911 13698
rect 6085 13640 6090 13696
rect 6146 13640 8850 13696
rect 8906 13640 8911 13696
rect 6085 13638 8911 13640
rect 6085 13635 6151 13638
rect 8845 13635 8911 13638
rect 17953 13698 18019 13701
rect 18812 13698 19612 13728
rect 17953 13696 19612 13698
rect 17953 13640 17958 13696
rect 18014 13640 19612 13696
rect 17953 13638 19612 13640
rect 17953 13635 18019 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 18812 13608 19612 13638
rect 4210 13567 4526 13568
rect 5758 13500 5764 13564
rect 5828 13562 5834 13564
rect 11646 13562 11652 13564
rect 5828 13502 11652 13562
rect 5828 13500 5834 13502
rect 11646 13500 11652 13502
rect 11716 13500 11722 13564
rect 2221 13426 2287 13429
rect 7966 13426 7972 13428
rect 2221 13424 7972 13426
rect 2221 13368 2226 13424
rect 2282 13368 7972 13424
rect 2221 13366 7972 13368
rect 2221 13363 2287 13366
rect 7966 13364 7972 13366
rect 8036 13364 8042 13428
rect 8477 13426 8543 13429
rect 9213 13426 9279 13429
rect 8477 13424 9279 13426
rect 8477 13368 8482 13424
rect 8538 13368 9218 13424
rect 9274 13368 9279 13424
rect 8477 13366 9279 13368
rect 8477 13363 8543 13366
rect 9213 13363 9279 13366
rect 9622 13364 9628 13428
rect 9692 13426 9698 13428
rect 9765 13426 9831 13429
rect 9692 13424 9831 13426
rect 9692 13368 9770 13424
rect 9826 13368 9831 13424
rect 9692 13366 9831 13368
rect 9692 13364 9698 13366
rect 9765 13363 9831 13366
rect 8293 13290 8359 13293
rect 4708 13288 8359 13290
rect 4708 13232 8298 13288
rect 8354 13232 8359 13288
rect 4708 13230 8359 13232
rect 3734 13092 3740 13156
rect 3804 13154 3810 13156
rect 4708 13154 4768 13230
rect 8293 13227 8359 13230
rect 8477 13290 8543 13293
rect 9581 13290 9647 13293
rect 8477 13288 9647 13290
rect 8477 13232 8482 13288
rect 8538 13232 9586 13288
rect 9642 13232 9647 13288
rect 8477 13230 9647 13232
rect 8477 13227 8543 13230
rect 9581 13227 9647 13230
rect 10409 13290 10475 13293
rect 11329 13290 11395 13293
rect 10409 13288 11395 13290
rect 10409 13232 10414 13288
rect 10470 13232 11334 13288
rect 11390 13232 11395 13288
rect 10409 13230 11395 13232
rect 10409 13227 10475 13230
rect 11329 13227 11395 13230
rect 11145 13156 11211 13157
rect 11094 13154 11100 13156
rect 3804 13094 4768 13154
rect 11054 13094 11100 13154
rect 11164 13152 11211 13156
rect 11206 13096 11211 13152
rect 3804 13092 3810 13094
rect 11094 13092 11100 13094
rect 11164 13092 11211 13096
rect 11145 13091 11211 13092
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 2865 13018 2931 13021
rect 2865 13016 4124 13018
rect 2865 12960 2870 13016
rect 2926 12960 4124 13016
rect 2865 12958 4124 12960
rect 2865 12955 2931 12958
rect 3141 12882 3207 12885
rect 3366 12882 3372 12884
rect 3141 12880 3372 12882
rect 3141 12824 3146 12880
rect 3202 12824 3372 12880
rect 3141 12822 3372 12824
rect 3141 12819 3207 12822
rect 3366 12820 3372 12822
rect 3436 12882 3442 12884
rect 3918 12882 3924 12884
rect 3436 12822 3924 12882
rect 3436 12820 3442 12822
rect 3918 12820 3924 12822
rect 3988 12820 3994 12884
rect 4064 12882 4124 12958
rect 7046 12882 7052 12884
rect 4064 12822 7052 12882
rect 7046 12820 7052 12822
rect 7116 12820 7122 12884
rect 8334 12882 8340 12884
rect 8204 12822 8340 12882
rect 8204 12749 8264 12822
rect 8334 12820 8340 12822
rect 8404 12820 8410 12884
rect 13854 12820 13860 12884
rect 13924 12882 13930 12884
rect 14825 12882 14891 12885
rect 13924 12880 14891 12882
rect 13924 12824 14830 12880
rect 14886 12824 14891 12880
rect 13924 12822 14891 12824
rect 13924 12820 13930 12822
rect 14825 12819 14891 12822
rect 8201 12744 8267 12749
rect 8201 12688 8206 12744
rect 8262 12688 8267 12744
rect 8201 12683 8267 12688
rect 8334 12684 8340 12748
rect 8404 12746 8410 12748
rect 9213 12746 9279 12749
rect 8404 12744 9279 12746
rect 8404 12688 9218 12744
rect 9274 12688 9279 12744
rect 8404 12686 9279 12688
rect 8404 12684 8410 12686
rect 9213 12683 9279 12686
rect 17309 12746 17375 12749
rect 17534 12746 17540 12748
rect 17309 12744 17540 12746
rect 17309 12688 17314 12744
rect 17370 12688 17540 12744
rect 17309 12686 17540 12688
rect 17309 12683 17375 12686
rect 17534 12684 17540 12686
rect 17604 12684 17610 12748
rect 5390 12548 5396 12612
rect 5460 12610 5466 12612
rect 6085 12610 6151 12613
rect 5460 12608 6151 12610
rect 5460 12552 6090 12608
rect 6146 12552 6151 12608
rect 5460 12550 6151 12552
rect 5460 12548 5466 12550
rect 6085 12547 6151 12550
rect 6545 12610 6611 12613
rect 9029 12612 9095 12613
rect 9029 12610 9076 12612
rect 6545 12608 7850 12610
rect 6545 12552 6550 12608
rect 6606 12552 7850 12608
rect 6545 12550 7850 12552
rect 8984 12608 9076 12610
rect 8984 12552 9034 12608
rect 8984 12550 9076 12552
rect 6545 12547 6611 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 6545 12474 6611 12477
rect 7557 12474 7623 12477
rect 6545 12472 7623 12474
rect 6545 12416 6550 12472
rect 6606 12416 7562 12472
rect 7618 12416 7623 12472
rect 6545 12414 7623 12416
rect 6545 12411 6611 12414
rect 7557 12411 7623 12414
rect 2865 12340 2931 12341
rect 2814 12338 2820 12340
rect 2774 12278 2820 12338
rect 2884 12336 2931 12340
rect 2926 12280 2931 12336
rect 2814 12276 2820 12278
rect 2884 12276 2931 12280
rect 2865 12275 2931 12276
rect 3877 12338 3943 12341
rect 4245 12338 4311 12341
rect 3877 12336 4311 12338
rect 3877 12280 3882 12336
rect 3938 12280 4250 12336
rect 4306 12280 4311 12336
rect 3877 12278 4311 12280
rect 3877 12275 3943 12278
rect 4245 12275 4311 12278
rect 7046 12276 7052 12340
rect 7116 12338 7122 12340
rect 7373 12338 7439 12341
rect 7116 12336 7439 12338
rect 7116 12280 7378 12336
rect 7434 12280 7439 12336
rect 7116 12278 7439 12280
rect 7790 12338 7850 12550
rect 9029 12548 9076 12550
rect 9140 12548 9146 12612
rect 9213 12610 9279 12613
rect 9581 12610 9647 12613
rect 9213 12608 9647 12610
rect 9213 12552 9218 12608
rect 9274 12552 9586 12608
rect 9642 12552 9647 12608
rect 9213 12550 9647 12552
rect 9029 12547 9095 12548
rect 9213 12547 9279 12550
rect 9581 12547 9647 12550
rect 8937 12474 9003 12477
rect 9070 12474 9076 12476
rect 8937 12472 9076 12474
rect 8937 12416 8942 12472
rect 8998 12416 9076 12472
rect 8937 12414 9076 12416
rect 8937 12411 9003 12414
rect 9070 12412 9076 12414
rect 9140 12412 9146 12476
rect 11145 12474 11211 12477
rect 12249 12474 12315 12477
rect 11145 12472 12315 12474
rect 11145 12416 11150 12472
rect 11206 12416 12254 12472
rect 12310 12416 12315 12472
rect 11145 12414 12315 12416
rect 11145 12411 11211 12414
rect 12249 12411 12315 12414
rect 12382 12412 12388 12476
rect 12452 12474 12458 12476
rect 13077 12474 13143 12477
rect 12452 12472 13143 12474
rect 12452 12416 13082 12472
rect 13138 12416 13143 12472
rect 12452 12414 13143 12416
rect 12452 12412 12458 12414
rect 13077 12411 13143 12414
rect 11278 12338 11284 12340
rect 7790 12278 11284 12338
rect 7116 12276 7122 12278
rect 7373 12275 7439 12278
rect 11278 12276 11284 12278
rect 11348 12338 11354 12340
rect 11973 12338 12039 12341
rect 11348 12336 12039 12338
rect 11348 12280 11978 12336
rect 12034 12280 12039 12336
rect 11348 12278 12039 12280
rect 11348 12276 11354 12278
rect 11973 12275 12039 12278
rect 12157 12338 12223 12341
rect 14733 12338 14799 12341
rect 12157 12336 14799 12338
rect 12157 12280 12162 12336
rect 12218 12280 14738 12336
rect 14794 12280 14799 12336
rect 12157 12278 14799 12280
rect 12157 12275 12223 12278
rect 14733 12275 14799 12278
rect 18045 12338 18111 12341
rect 18812 12338 19612 12368
rect 18045 12336 19612 12338
rect 18045 12280 18050 12336
rect 18106 12280 19612 12336
rect 18045 12278 19612 12280
rect 18045 12275 18111 12278
rect 18812 12248 19612 12278
rect 3785 12202 3851 12205
rect 6361 12202 6427 12205
rect 3785 12200 6427 12202
rect 3785 12144 3790 12200
rect 3846 12144 6366 12200
rect 6422 12144 6427 12200
rect 3785 12142 6427 12144
rect 3785 12139 3851 12142
rect 6361 12139 6427 12142
rect 8845 12202 8911 12205
rect 10174 12202 10180 12204
rect 8845 12200 10180 12202
rect 8845 12144 8850 12200
rect 8906 12144 10180 12200
rect 8845 12142 10180 12144
rect 8845 12139 8911 12142
rect 10174 12140 10180 12142
rect 10244 12140 10250 12204
rect 11237 12202 11303 12205
rect 11881 12202 11947 12205
rect 12985 12202 13051 12205
rect 11237 12200 13051 12202
rect 11237 12144 11242 12200
rect 11298 12144 11886 12200
rect 11942 12144 12990 12200
rect 13046 12144 13051 12200
rect 11237 12142 13051 12144
rect 11237 12139 11303 12142
rect 11881 12139 11947 12142
rect 12985 12139 13051 12142
rect 4521 12066 4587 12069
rect 4654 12066 4660 12068
rect 4521 12064 4660 12066
rect 4521 12008 4526 12064
rect 4582 12008 4660 12064
rect 4521 12006 4660 12008
rect 4521 12003 4587 12006
rect 4654 12004 4660 12006
rect 4724 12004 4730 12068
rect 8937 12066 9003 12069
rect 5260 12064 9003 12066
rect 5260 12008 8942 12064
rect 8998 12008 9003 12064
rect 5260 12006 9003 12008
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 4153 11794 4219 11797
rect 5260 11794 5320 12006
rect 8937 12003 9003 12006
rect 6361 11930 6427 11933
rect 11145 11930 11211 11933
rect 6361 11928 11211 11930
rect 6361 11872 6366 11928
rect 6422 11872 11150 11928
rect 11206 11872 11211 11928
rect 6361 11870 11211 11872
rect 6361 11867 6427 11870
rect 11145 11867 11211 11870
rect 11881 11930 11947 11933
rect 12893 11930 12959 11933
rect 13445 11930 13511 11933
rect 11881 11928 13511 11930
rect 11881 11872 11886 11928
rect 11942 11872 12898 11928
rect 12954 11872 13450 11928
rect 13506 11872 13511 11928
rect 11881 11870 13511 11872
rect 11881 11867 11947 11870
rect 12893 11867 12959 11870
rect 13445 11867 13511 11870
rect 4153 11792 5320 11794
rect 4153 11736 4158 11792
rect 4214 11736 5320 11792
rect 4153 11734 5320 11736
rect 5441 11794 5507 11797
rect 9029 11796 9095 11797
rect 5441 11792 6056 11794
rect 5441 11736 5446 11792
rect 5502 11736 6056 11792
rect 5441 11734 6056 11736
rect 4153 11731 4219 11734
rect 5441 11731 5507 11734
rect 0 11658 800 11688
rect 5996 11661 6056 11734
rect 9029 11792 9076 11796
rect 9140 11794 9146 11796
rect 14549 11794 14615 11797
rect 9029 11736 9034 11792
rect 9029 11732 9076 11736
rect 9140 11734 9186 11794
rect 9400 11792 14615 11794
rect 9400 11736 14554 11792
rect 14610 11736 14615 11792
rect 9400 11734 14615 11736
rect 9140 11732 9146 11734
rect 9029 11731 9095 11732
rect 9400 11661 9460 11734
rect 14549 11731 14615 11734
rect 1117 11658 1183 11661
rect 0 11656 1183 11658
rect 0 11600 1122 11656
rect 1178 11600 1183 11656
rect 0 11598 1183 11600
rect 0 11568 800 11598
rect 1117 11595 1183 11598
rect 4245 11658 4311 11661
rect 5165 11658 5231 11661
rect 5390 11658 5396 11660
rect 4245 11656 4722 11658
rect 4245 11600 4250 11656
rect 4306 11600 4722 11656
rect 4245 11598 4722 11600
rect 4245 11595 4311 11598
rect 4662 11522 4722 11598
rect 5165 11656 5396 11658
rect 5165 11600 5170 11656
rect 5226 11600 5396 11656
rect 5165 11598 5396 11600
rect 5165 11595 5231 11598
rect 5390 11596 5396 11598
rect 5460 11596 5466 11660
rect 5993 11658 6059 11661
rect 9397 11658 9463 11661
rect 5993 11656 9463 11658
rect 5993 11600 5998 11656
rect 6054 11600 9402 11656
rect 9458 11600 9463 11656
rect 5993 11598 9463 11600
rect 5993 11595 6059 11598
rect 9397 11595 9463 11598
rect 12525 11658 12591 11661
rect 13077 11658 13143 11661
rect 12525 11656 13143 11658
rect 12525 11600 12530 11656
rect 12586 11600 13082 11656
rect 13138 11600 13143 11656
rect 12525 11598 13143 11600
rect 12525 11595 12591 11598
rect 13077 11595 13143 11598
rect 13261 11658 13327 11661
rect 15929 11660 15995 11661
rect 15878 11658 15884 11660
rect 13261 11656 15884 11658
rect 15948 11658 15995 11660
rect 15948 11656 16040 11658
rect 13261 11600 13266 11656
rect 13322 11600 15884 11656
rect 15990 11600 16040 11656
rect 13261 11598 15884 11600
rect 13261 11595 13327 11598
rect 15878 11596 15884 11598
rect 15948 11598 16040 11600
rect 15948 11596 15995 11598
rect 15929 11595 15995 11596
rect 5390 11522 5396 11524
rect 4662 11462 5396 11522
rect 5390 11460 5396 11462
rect 5460 11522 5466 11524
rect 7557 11522 7623 11525
rect 9213 11522 9279 11525
rect 9857 11522 9923 11525
rect 5460 11520 7623 11522
rect 5460 11464 7562 11520
rect 7618 11464 7623 11520
rect 5460 11462 7623 11464
rect 5460 11460 5466 11462
rect 7557 11459 7623 11462
rect 8250 11520 9923 11522
rect 8250 11464 9218 11520
rect 9274 11464 9862 11520
rect 9918 11464 9923 11520
rect 8250 11462 9923 11464
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 6269 11386 6335 11389
rect 8250 11386 8310 11462
rect 9213 11459 9279 11462
rect 9857 11459 9923 11462
rect 11329 11522 11395 11525
rect 13537 11522 13603 11525
rect 14825 11522 14891 11525
rect 11329 11520 14891 11522
rect 11329 11464 11334 11520
rect 11390 11464 13542 11520
rect 13598 11464 14830 11520
rect 14886 11464 14891 11520
rect 11329 11462 14891 11464
rect 11329 11459 11395 11462
rect 13537 11459 13603 11462
rect 14825 11459 14891 11462
rect 6269 11384 8310 11386
rect 6269 11328 6274 11384
rect 6330 11328 8310 11384
rect 6269 11326 8310 11328
rect 9121 11386 9187 11389
rect 16113 11388 16179 11389
rect 9438 11386 9444 11388
rect 9121 11384 9444 11386
rect 9121 11328 9126 11384
rect 9182 11328 9444 11384
rect 9121 11326 9444 11328
rect 6269 11323 6335 11326
rect 9121 11323 9187 11326
rect 9438 11324 9444 11326
rect 9508 11324 9514 11388
rect 16062 11386 16068 11388
rect 16022 11326 16068 11386
rect 16132 11384 16179 11388
rect 16174 11328 16179 11384
rect 16062 11324 16068 11326
rect 16132 11324 16179 11328
rect 16113 11323 16179 11324
rect 6361 11250 6427 11253
rect 5398 11248 6427 11250
rect 5398 11192 6366 11248
rect 6422 11192 6427 11248
rect 5398 11190 6427 11192
rect 4654 11052 4660 11116
rect 4724 11114 4730 11116
rect 4981 11114 5047 11117
rect 5398 11114 5458 11190
rect 6361 11187 6427 11190
rect 7925 11250 7991 11253
rect 8150 11250 8156 11252
rect 7925 11248 8156 11250
rect 7925 11192 7930 11248
rect 7986 11192 8156 11248
rect 7925 11190 8156 11192
rect 7925 11187 7991 11190
rect 8150 11188 8156 11190
rect 8220 11188 8226 11252
rect 8886 11188 8892 11252
rect 8956 11250 8962 11252
rect 10133 11250 10199 11253
rect 8956 11248 10199 11250
rect 8956 11192 10138 11248
rect 10194 11192 10199 11248
rect 8956 11190 10199 11192
rect 8956 11188 8962 11190
rect 10133 11187 10199 11190
rect 10501 11250 10567 11253
rect 16573 11250 16639 11253
rect 10501 11248 16639 11250
rect 10501 11192 10506 11248
rect 10562 11192 16578 11248
rect 16634 11192 16639 11248
rect 10501 11190 16639 11192
rect 10501 11187 10567 11190
rect 16573 11187 16639 11190
rect 4724 11112 5458 11114
rect 4724 11056 4986 11112
rect 5042 11056 5458 11112
rect 4724 11054 5458 11056
rect 6729 11114 6795 11117
rect 9673 11114 9739 11117
rect 10593 11116 10659 11117
rect 10542 11114 10548 11116
rect 6729 11112 9739 11114
rect 6729 11056 6734 11112
rect 6790 11056 9678 11112
rect 9734 11056 9739 11112
rect 6729 11054 9739 11056
rect 10502 11054 10548 11114
rect 10612 11112 10659 11116
rect 10654 11056 10659 11112
rect 4724 11052 4730 11054
rect 4981 11051 5047 11054
rect 6729 11051 6795 11054
rect 9673 11051 9739 11054
rect 10542 11052 10548 11054
rect 10612 11052 10659 11056
rect 10593 11051 10659 11052
rect 7373 10978 7439 10981
rect 9806 10978 9812 10980
rect 7373 10976 9812 10978
rect 7373 10920 7378 10976
rect 7434 10920 9812 10976
rect 7373 10918 9812 10920
rect 7373 10915 7439 10918
rect 9806 10916 9812 10918
rect 9876 10978 9882 10980
rect 10593 10978 10659 10981
rect 9876 10976 10659 10978
rect 9876 10920 10598 10976
rect 10654 10920 10659 10976
rect 9876 10918 10659 10920
rect 9876 10916 9882 10918
rect 10593 10915 10659 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 5533 10842 5599 10845
rect 8845 10842 8911 10845
rect 5533 10840 8911 10842
rect 5533 10784 5538 10840
rect 5594 10784 8850 10840
rect 8906 10784 8911 10840
rect 5533 10782 8911 10784
rect 5533 10779 5599 10782
rect 8845 10779 8911 10782
rect 3693 10706 3759 10709
rect 8518 10706 8524 10708
rect 3693 10704 8524 10706
rect 3693 10648 3698 10704
rect 3754 10648 8524 10704
rect 3693 10646 8524 10648
rect 3693 10643 3759 10646
rect 8518 10644 8524 10646
rect 8588 10706 8594 10708
rect 15009 10706 15075 10709
rect 8588 10704 15075 10706
rect 8588 10648 15014 10704
rect 15070 10648 15075 10704
rect 8588 10646 15075 10648
rect 8588 10644 8594 10646
rect 15009 10643 15075 10646
rect 3969 10570 4035 10573
rect 5942 10570 5948 10572
rect 3969 10568 5948 10570
rect 3969 10512 3974 10568
rect 4030 10512 5948 10568
rect 3969 10510 5948 10512
rect 3969 10507 4035 10510
rect 5942 10508 5948 10510
rect 6012 10570 6018 10572
rect 6177 10570 6243 10573
rect 6012 10568 6243 10570
rect 6012 10512 6182 10568
rect 6238 10512 6243 10568
rect 6012 10510 6243 10512
rect 6012 10508 6018 10510
rect 6177 10507 6243 10510
rect 8201 10570 8267 10573
rect 8845 10570 8911 10573
rect 8201 10568 8911 10570
rect 8201 10512 8206 10568
rect 8262 10512 8850 10568
rect 8906 10512 8911 10568
rect 8201 10510 8911 10512
rect 8201 10507 8267 10510
rect 8845 10507 8911 10510
rect 5809 10434 5875 10437
rect 10225 10434 10291 10437
rect 5809 10432 10291 10434
rect 5809 10376 5814 10432
rect 5870 10376 10230 10432
rect 10286 10376 10291 10432
rect 5809 10374 10291 10376
rect 5809 10371 5875 10374
rect 10225 10371 10291 10374
rect 11646 10372 11652 10436
rect 11716 10434 11722 10436
rect 17677 10434 17743 10437
rect 11716 10432 17743 10434
rect 11716 10376 17682 10432
rect 17738 10376 17743 10432
rect 11716 10374 17743 10376
rect 11716 10372 11722 10374
rect 17677 10371 17743 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4981 10298 5047 10301
rect 7465 10298 7531 10301
rect 4981 10296 7531 10298
rect 4981 10240 4986 10296
rect 5042 10240 7470 10296
rect 7526 10240 7531 10296
rect 4981 10238 7531 10240
rect 4981 10235 5047 10238
rect 7465 10235 7531 10238
rect 9254 10236 9260 10300
rect 9324 10298 9330 10300
rect 9397 10298 9463 10301
rect 9324 10296 9463 10298
rect 9324 10240 9402 10296
rect 9458 10240 9463 10296
rect 9324 10238 9463 10240
rect 9324 10236 9330 10238
rect 9397 10235 9463 10238
rect 3734 10100 3740 10164
rect 3804 10162 3810 10164
rect 4337 10162 4403 10165
rect 3804 10160 4403 10162
rect 3804 10104 4342 10160
rect 4398 10104 4403 10160
rect 3804 10102 4403 10104
rect 3804 10100 3810 10102
rect 4337 10099 4403 10102
rect 4797 10162 4863 10165
rect 8845 10162 8911 10165
rect 9990 10162 9996 10164
rect 4797 10160 6930 10162
rect 4797 10104 4802 10160
rect 4858 10104 6930 10160
rect 4797 10102 6930 10104
rect 4797 10099 4863 10102
rect 2129 10026 2195 10029
rect 6729 10026 6795 10029
rect 2129 10024 6795 10026
rect 2129 9968 2134 10024
rect 2190 9968 6734 10024
rect 6790 9968 6795 10024
rect 2129 9966 6795 9968
rect 2129 9963 2195 9966
rect 6729 9963 6795 9966
rect 6729 9890 6795 9893
rect 6870 9890 6930 10102
rect 8845 10160 9996 10162
rect 8845 10104 8850 10160
rect 8906 10104 9996 10160
rect 8845 10102 9996 10104
rect 8845 10099 8911 10102
rect 9990 10100 9996 10102
rect 10060 10162 10066 10164
rect 10133 10162 10199 10165
rect 10060 10160 10199 10162
rect 10060 10104 10138 10160
rect 10194 10104 10199 10160
rect 10060 10102 10199 10104
rect 10060 10100 10066 10102
rect 10133 10099 10199 10102
rect 10869 10164 10935 10165
rect 15193 10164 15259 10165
rect 10869 10160 10916 10164
rect 10980 10162 10986 10164
rect 10869 10104 10874 10160
rect 10869 10100 10916 10104
rect 10980 10102 11026 10162
rect 10980 10100 10986 10102
rect 15142 10100 15148 10164
rect 15212 10162 15259 10164
rect 15212 10160 15304 10162
rect 15254 10104 15304 10160
rect 15212 10102 15304 10104
rect 15212 10100 15259 10102
rect 10869 10099 10935 10100
rect 15193 10099 15259 10100
rect 8109 10026 8175 10029
rect 8569 10026 8635 10029
rect 8109 10024 8635 10026
rect 8109 9968 8114 10024
rect 8170 9968 8574 10024
rect 8630 9968 8635 10024
rect 8109 9966 8635 9968
rect 8109 9963 8175 9966
rect 8569 9963 8635 9966
rect 9857 10026 9923 10029
rect 10685 10026 10751 10029
rect 9857 10024 10751 10026
rect 9857 9968 9862 10024
rect 9918 9968 10690 10024
rect 10746 9968 10751 10024
rect 9857 9966 10751 9968
rect 9857 9963 9923 9966
rect 10685 9963 10751 9966
rect 14457 10026 14523 10029
rect 17861 10026 17927 10029
rect 14457 10024 17927 10026
rect 14457 9968 14462 10024
rect 14518 9968 17866 10024
rect 17922 9968 17927 10024
rect 14457 9966 17927 9968
rect 14457 9963 14523 9966
rect 17861 9963 17927 9966
rect 7189 9890 7255 9893
rect 6729 9888 7255 9890
rect 6729 9832 6734 9888
rect 6790 9832 7194 9888
rect 7250 9832 7255 9888
rect 6729 9830 7255 9832
rect 6729 9827 6795 9830
rect 7189 9827 7255 9830
rect 10317 9890 10383 9893
rect 14089 9890 14155 9893
rect 10317 9888 14155 9890
rect 10317 9832 10322 9888
rect 10378 9832 14094 9888
rect 14150 9832 14155 9888
rect 10317 9830 14155 9832
rect 10317 9827 10383 9830
rect 14089 9827 14155 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 6637 9756 6703 9757
rect 6637 9752 6684 9756
rect 6748 9754 6754 9756
rect 10501 9754 10567 9757
rect 11094 9754 11100 9756
rect 6637 9696 6642 9752
rect 6637 9692 6684 9696
rect 6748 9694 6794 9754
rect 10501 9752 11100 9754
rect 10501 9696 10506 9752
rect 10562 9696 11100 9752
rect 10501 9694 11100 9696
rect 6748 9692 6754 9694
rect 6637 9691 6703 9692
rect 10501 9691 10567 9694
rect 11094 9692 11100 9694
rect 11164 9692 11170 9756
rect 13169 9754 13235 9757
rect 16665 9754 16731 9757
rect 17585 9754 17651 9757
rect 13169 9752 17651 9754
rect 13169 9696 13174 9752
rect 13230 9696 16670 9752
rect 16726 9696 17590 9752
rect 17646 9696 17651 9752
rect 13169 9694 17651 9696
rect 13169 9691 13235 9694
rect 16665 9691 16731 9694
rect 17585 9691 17651 9694
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 3601 9618 3667 9621
rect 8937 9618 9003 9621
rect 16849 9618 16915 9621
rect 17217 9620 17283 9621
rect 17585 9620 17651 9621
rect 17166 9618 17172 9620
rect 3601 9616 7666 9618
rect 3601 9560 3606 9616
rect 3662 9560 7666 9616
rect 3601 9558 7666 9560
rect 3601 9555 3667 9558
rect 2589 9482 2655 9485
rect 7281 9482 7347 9485
rect 2589 9480 7347 9482
rect 2589 9424 2594 9480
rect 2650 9424 7286 9480
rect 7342 9424 7347 9480
rect 2589 9422 7347 9424
rect 7606 9482 7666 9558
rect 8937 9616 16915 9618
rect 8937 9560 8942 9616
rect 8998 9560 16854 9616
rect 16910 9560 16915 9616
rect 8937 9558 16915 9560
rect 17126 9558 17172 9618
rect 17236 9616 17283 9620
rect 17534 9618 17540 9620
rect 17278 9560 17283 9616
rect 8937 9555 9003 9558
rect 16849 9555 16915 9558
rect 17166 9556 17172 9558
rect 17236 9556 17283 9560
rect 17494 9558 17540 9618
rect 17604 9616 17651 9620
rect 17646 9560 17651 9616
rect 17534 9556 17540 9558
rect 17604 9556 17651 9560
rect 17217 9555 17283 9556
rect 17585 9555 17651 9556
rect 11053 9482 11119 9485
rect 7606 9480 11119 9482
rect 7606 9424 11058 9480
rect 11114 9424 11119 9480
rect 7606 9422 11119 9424
rect 2589 9419 2655 9422
rect 7281 9419 7347 9422
rect 11053 9419 11119 9422
rect 11973 9482 12039 9485
rect 13169 9482 13235 9485
rect 11973 9480 13235 9482
rect 11973 9424 11978 9480
rect 12034 9424 13174 9480
rect 13230 9424 13235 9480
rect 11973 9422 13235 9424
rect 11973 9419 12039 9422
rect 13169 9419 13235 9422
rect 13629 9484 13695 9485
rect 13629 9480 13676 9484
rect 13740 9482 13746 9484
rect 13629 9424 13634 9480
rect 13629 9420 13676 9424
rect 13740 9422 13786 9482
rect 13740 9420 13746 9422
rect 13629 9419 13695 9420
rect 5165 9346 5231 9349
rect 5390 9346 5396 9348
rect 5165 9344 5396 9346
rect 5165 9288 5170 9344
rect 5226 9288 5396 9344
rect 5165 9286 5396 9288
rect 5165 9283 5231 9286
rect 5390 9284 5396 9286
rect 5460 9284 5466 9348
rect 5901 9346 5967 9349
rect 7925 9346 7991 9349
rect 5901 9344 7991 9346
rect 5901 9288 5906 9344
rect 5962 9288 7930 9344
rect 7986 9288 7991 9344
rect 5901 9286 7991 9288
rect 5901 9283 5967 9286
rect 7925 9283 7991 9286
rect 9438 9284 9444 9348
rect 9508 9346 9514 9348
rect 10225 9346 10291 9349
rect 9508 9344 10291 9346
rect 9508 9288 10230 9344
rect 10286 9288 10291 9344
rect 9508 9286 10291 9288
rect 9508 9284 9514 9286
rect 10225 9283 10291 9286
rect 11513 9346 11579 9349
rect 13537 9346 13603 9349
rect 11513 9344 13603 9346
rect 11513 9288 11518 9344
rect 11574 9288 13542 9344
rect 13598 9288 13603 9344
rect 11513 9286 13603 9288
rect 11513 9283 11579 9286
rect 13537 9283 13603 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 6545 9210 6611 9213
rect 7046 9210 7052 9212
rect 6545 9208 7052 9210
rect 6545 9152 6550 9208
rect 6606 9152 7052 9208
rect 6545 9150 7052 9152
rect 6545 9147 6611 9150
rect 7046 9148 7052 9150
rect 7116 9148 7122 9212
rect 11053 9210 11119 9213
rect 11462 9210 11468 9212
rect 11053 9208 11468 9210
rect 11053 9152 11058 9208
rect 11114 9152 11468 9208
rect 11053 9150 11468 9152
rect 11053 9147 11119 9150
rect 11462 9148 11468 9150
rect 11532 9148 11538 9212
rect 12249 9210 12315 9213
rect 13537 9210 13603 9213
rect 15837 9210 15903 9213
rect 12249 9208 15903 9210
rect 12249 9152 12254 9208
rect 12310 9152 13542 9208
rect 13598 9152 15842 9208
rect 15898 9152 15903 9208
rect 12249 9150 15903 9152
rect 12249 9147 12315 9150
rect 13537 9147 13603 9150
rect 15837 9147 15903 9150
rect 2313 9074 2379 9077
rect 15469 9074 15535 9077
rect 16573 9074 16639 9077
rect 2313 9072 16639 9074
rect 2313 9016 2318 9072
rect 2374 9016 15474 9072
rect 15530 9016 16578 9072
rect 16634 9016 16639 9072
rect 2313 9014 16639 9016
rect 2313 9011 2379 9014
rect 15469 9011 15535 9014
rect 16573 9011 16639 9014
rect 4337 8938 4403 8941
rect 6637 8938 6703 8941
rect 10317 8940 10383 8941
rect 10317 8938 10364 8940
rect 4337 8936 6703 8938
rect 4337 8880 4342 8936
rect 4398 8880 6642 8936
rect 6698 8880 6703 8936
rect 4337 8878 6703 8880
rect 10272 8936 10364 8938
rect 10428 8938 10434 8940
rect 11094 8938 11100 8940
rect 10272 8880 10322 8936
rect 10272 8878 10364 8880
rect 4337 8875 4403 8878
rect 6637 8875 6703 8878
rect 10317 8876 10364 8878
rect 10428 8878 11100 8938
rect 10428 8876 10434 8878
rect 11094 8876 11100 8878
rect 11164 8876 11170 8940
rect 12893 8938 12959 8941
rect 11286 8936 12959 8938
rect 11286 8880 12898 8936
rect 12954 8880 12959 8936
rect 11286 8878 12959 8880
rect 10317 8875 10383 8876
rect 5942 8740 5948 8804
rect 6012 8802 6018 8804
rect 6085 8802 6151 8805
rect 6012 8800 6151 8802
rect 6012 8744 6090 8800
rect 6146 8744 6151 8800
rect 6012 8742 6151 8744
rect 6012 8740 6018 8742
rect 6085 8739 6151 8742
rect 9029 8802 9095 8805
rect 9305 8802 9371 8805
rect 9029 8800 9371 8802
rect 9029 8744 9034 8800
rect 9090 8744 9310 8800
rect 9366 8744 9371 8800
rect 9029 8742 9371 8744
rect 9029 8739 9095 8742
rect 9305 8739 9371 8742
rect 9949 8802 10015 8805
rect 11286 8802 11346 8878
rect 12893 8875 12959 8878
rect 9949 8800 11346 8802
rect 9949 8744 9954 8800
rect 10010 8744 11346 8800
rect 9949 8742 11346 8744
rect 12249 8802 12315 8805
rect 16389 8802 16455 8805
rect 12249 8800 16455 8802
rect 12249 8744 12254 8800
rect 12310 8744 16394 8800
rect 16450 8744 16455 8800
rect 12249 8742 16455 8744
rect 9949 8739 10015 8742
rect 12249 8739 12315 8742
rect 16389 8739 16455 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 5717 8666 5783 8669
rect 7741 8666 7807 8669
rect 5717 8664 7807 8666
rect 5717 8608 5722 8664
rect 5778 8608 7746 8664
rect 7802 8608 7807 8664
rect 5717 8606 7807 8608
rect 5717 8603 5783 8606
rect 7741 8603 7807 8606
rect 8937 8666 9003 8669
rect 9857 8666 9923 8669
rect 8937 8664 9923 8666
rect 8937 8608 8942 8664
rect 8998 8608 9862 8664
rect 9918 8608 9923 8664
rect 8937 8606 9923 8608
rect 8937 8603 9003 8606
rect 9857 8603 9923 8606
rect 11053 8666 11119 8669
rect 11605 8666 11671 8669
rect 17125 8666 17191 8669
rect 11053 8664 17191 8666
rect 11053 8608 11058 8664
rect 11114 8608 11610 8664
rect 11666 8608 17130 8664
rect 17186 8608 17191 8664
rect 11053 8606 17191 8608
rect 11053 8603 11119 8606
rect 11605 8603 11671 8606
rect 17125 8603 17191 8606
rect 3877 8530 3943 8533
rect 4613 8530 4679 8533
rect 6177 8530 6243 8533
rect 7741 8530 7807 8533
rect 3877 8528 5320 8530
rect 3877 8472 3882 8528
rect 3938 8472 4618 8528
rect 4674 8472 5320 8528
rect 3877 8470 5320 8472
rect 3877 8467 3943 8470
rect 4613 8467 4679 8470
rect 5260 8397 5320 8470
rect 6177 8528 7807 8530
rect 6177 8472 6182 8528
rect 6238 8472 7746 8528
rect 7802 8472 7807 8528
rect 6177 8470 7807 8472
rect 6177 8467 6243 8470
rect 7741 8467 7807 8470
rect 9857 8530 9923 8533
rect 16062 8530 16068 8532
rect 9857 8528 16068 8530
rect 9857 8472 9862 8528
rect 9918 8472 16068 8528
rect 9857 8470 16068 8472
rect 9857 8467 9923 8470
rect 16062 8468 16068 8470
rect 16132 8468 16138 8532
rect 5257 8394 5323 8397
rect 6678 8394 6684 8396
rect 5257 8392 6684 8394
rect 5257 8336 5262 8392
rect 5318 8336 6684 8392
rect 5257 8334 6684 8336
rect 5257 8331 5323 8334
rect 6678 8332 6684 8334
rect 6748 8394 6754 8396
rect 7833 8394 7899 8397
rect 6748 8392 7899 8394
rect 6748 8336 7838 8392
rect 7894 8336 7899 8392
rect 6748 8334 7899 8336
rect 6748 8332 6754 8334
rect 7833 8331 7899 8334
rect 8385 8394 8451 8397
rect 10317 8394 10383 8397
rect 8385 8392 10383 8394
rect 8385 8336 8390 8392
rect 8446 8336 10322 8392
rect 10378 8336 10383 8392
rect 8385 8334 10383 8336
rect 8385 8331 8451 8334
rect 10317 8331 10383 8334
rect 11145 8394 11211 8397
rect 11278 8394 11284 8396
rect 11145 8392 11284 8394
rect 11145 8336 11150 8392
rect 11206 8336 11284 8392
rect 11145 8334 11284 8336
rect 11145 8331 11211 8334
rect 11278 8332 11284 8334
rect 11348 8332 11354 8396
rect 11881 8394 11947 8397
rect 14365 8394 14431 8397
rect 11881 8392 14431 8394
rect 11881 8336 11886 8392
rect 11942 8336 14370 8392
rect 14426 8336 14431 8392
rect 11881 8334 14431 8336
rect 11881 8331 11947 8334
rect 14365 8331 14431 8334
rect 4613 8292 4679 8295
rect 4613 8290 4722 8292
rect 0 8258 800 8288
rect 1485 8258 1551 8261
rect 0 8256 1551 8258
rect 0 8200 1490 8256
rect 1546 8200 1551 8256
rect 4613 8234 4618 8290
rect 4674 8234 4722 8290
rect 4613 8229 4722 8234
rect 0 8198 1551 8200
rect 0 8168 800 8198
rect 1485 8195 1551 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4337 7986 4403 7989
rect 4662 7986 4722 8229
rect 4889 8258 4955 8261
rect 7925 8258 7991 8261
rect 4889 8256 7991 8258
rect 4889 8200 4894 8256
rect 4950 8200 7930 8256
rect 7986 8200 7991 8256
rect 4889 8198 7991 8200
rect 4889 8195 4955 8198
rect 7925 8195 7991 8198
rect 8109 8258 8175 8261
rect 9029 8258 9095 8261
rect 10685 8260 10751 8261
rect 10685 8258 10732 8260
rect 8109 8256 9095 8258
rect 8109 8200 8114 8256
rect 8170 8200 9034 8256
rect 9090 8200 9095 8256
rect 8109 8198 9095 8200
rect 10644 8256 10732 8258
rect 10796 8258 10802 8260
rect 15377 8258 15443 8261
rect 16849 8260 16915 8261
rect 16798 8258 16804 8260
rect 10796 8256 15443 8258
rect 10644 8200 10690 8256
rect 10796 8200 15382 8256
rect 15438 8200 15443 8256
rect 10644 8198 10732 8200
rect 8109 8195 8175 8198
rect 9029 8195 9095 8198
rect 10685 8196 10732 8198
rect 10796 8198 15443 8200
rect 16758 8198 16804 8258
rect 16868 8256 16915 8260
rect 16910 8200 16915 8256
rect 10796 8196 10802 8198
rect 10685 8195 10751 8196
rect 15377 8195 15443 8198
rect 16798 8196 16804 8198
rect 16868 8196 16915 8200
rect 16849 8195 16915 8196
rect 4981 8122 5047 8125
rect 6821 8122 6887 8125
rect 4981 8120 6887 8122
rect 4981 8064 4986 8120
rect 5042 8064 6826 8120
rect 6882 8064 6887 8120
rect 4981 8062 6887 8064
rect 4981 8059 5047 8062
rect 6821 8059 6887 8062
rect 7005 8122 7071 8125
rect 7189 8122 7255 8125
rect 7005 8120 7255 8122
rect 7005 8064 7010 8120
rect 7066 8064 7194 8120
rect 7250 8064 7255 8120
rect 7005 8062 7255 8064
rect 7005 8059 7071 8062
rect 7189 8059 7255 8062
rect 9581 8122 9647 8125
rect 12566 8122 12572 8124
rect 9581 8120 12572 8122
rect 9581 8064 9586 8120
rect 9642 8064 12572 8120
rect 9581 8062 12572 8064
rect 9581 8059 9647 8062
rect 12566 8060 12572 8062
rect 12636 8060 12642 8124
rect 4337 7984 4722 7986
rect 4337 7928 4342 7984
rect 4398 7928 4722 7984
rect 4337 7926 4722 7928
rect 5625 7986 5691 7989
rect 6126 7986 6132 7988
rect 5625 7984 6132 7986
rect 5625 7928 5630 7984
rect 5686 7928 6132 7984
rect 5625 7926 6132 7928
rect 4337 7923 4403 7926
rect 5625 7923 5691 7926
rect 6126 7924 6132 7926
rect 6196 7924 6202 7988
rect 6269 7986 6335 7989
rect 7649 7986 7715 7989
rect 9581 7986 9647 7989
rect 10409 7986 10475 7989
rect 11053 7986 11119 7989
rect 6269 7984 11119 7986
rect 6269 7928 6274 7984
rect 6330 7928 7654 7984
rect 7710 7928 9586 7984
rect 9642 7928 10414 7984
rect 10470 7928 11058 7984
rect 11114 7928 11119 7984
rect 6269 7926 11119 7928
rect 6269 7923 6335 7926
rect 7649 7923 7715 7926
rect 9581 7923 9647 7926
rect 10409 7923 10475 7926
rect 11053 7923 11119 7926
rect 11697 7986 11763 7989
rect 14549 7986 14615 7989
rect 11697 7984 14615 7986
rect 11697 7928 11702 7984
rect 11758 7928 14554 7984
rect 14610 7928 14615 7984
rect 11697 7926 14615 7928
rect 11697 7923 11763 7926
rect 14549 7923 14615 7926
rect 3417 7850 3483 7853
rect 6361 7850 6427 7853
rect 13537 7850 13603 7853
rect 3417 7848 5320 7850
rect 3417 7792 3422 7848
rect 3478 7792 5320 7848
rect 3417 7790 5320 7792
rect 3417 7787 3483 7790
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 1853 7578 1919 7581
rect 0 7576 1919 7578
rect 0 7520 1858 7576
rect 1914 7520 1919 7576
rect 0 7518 1919 7520
rect 5260 7578 5320 7790
rect 6361 7848 13603 7850
rect 6361 7792 6366 7848
rect 6422 7792 13542 7848
rect 13598 7792 13603 7848
rect 6361 7790 13603 7792
rect 6361 7787 6427 7790
rect 13537 7787 13603 7790
rect 5533 7714 5599 7717
rect 8109 7714 8175 7717
rect 5533 7712 8175 7714
rect 5533 7656 5538 7712
rect 5594 7656 8114 7712
rect 8170 7656 8175 7712
rect 5533 7654 8175 7656
rect 5533 7651 5599 7654
rect 8109 7651 8175 7654
rect 8845 7714 8911 7717
rect 14917 7714 14983 7717
rect 8845 7712 14983 7714
rect 8845 7656 8850 7712
rect 8906 7656 14922 7712
rect 14978 7656 14983 7712
rect 8845 7654 14983 7656
rect 8845 7651 8911 7654
rect 14917 7651 14983 7654
rect 6269 7578 6335 7581
rect 5260 7576 6335 7578
rect 5260 7520 6274 7576
rect 6330 7520 6335 7576
rect 5260 7518 6335 7520
rect 0 7488 800 7518
rect 1853 7515 1919 7518
rect 6269 7515 6335 7518
rect 7189 7578 7255 7581
rect 13997 7578 14063 7581
rect 15009 7578 15075 7581
rect 7189 7576 15075 7578
rect 7189 7520 7194 7576
rect 7250 7520 14002 7576
rect 14058 7520 15014 7576
rect 15070 7520 15075 7576
rect 7189 7518 15075 7520
rect 7189 7515 7255 7518
rect 13997 7515 14063 7518
rect 15009 7515 15075 7518
rect 18045 7578 18111 7581
rect 18812 7578 19612 7608
rect 18045 7576 19612 7578
rect 18045 7520 18050 7576
rect 18106 7520 19612 7576
rect 18045 7518 19612 7520
rect 18045 7515 18111 7518
rect 18812 7488 19612 7518
rect 4705 7442 4771 7445
rect 5073 7442 5139 7445
rect 4705 7440 5139 7442
rect 4705 7384 4710 7440
rect 4766 7384 5078 7440
rect 5134 7384 5139 7440
rect 4705 7382 5139 7384
rect 4705 7379 4771 7382
rect 5073 7379 5139 7382
rect 8201 7442 8267 7445
rect 8937 7442 9003 7445
rect 8201 7440 9003 7442
rect 8201 7384 8206 7440
rect 8262 7384 8942 7440
rect 8998 7384 9003 7440
rect 8201 7382 9003 7384
rect 8201 7379 8267 7382
rect 8937 7379 9003 7382
rect 9121 7442 9187 7445
rect 12341 7442 12407 7445
rect 9121 7440 12407 7442
rect 9121 7384 9126 7440
rect 9182 7384 12346 7440
rect 12402 7384 12407 7440
rect 9121 7382 12407 7384
rect 9121 7379 9187 7382
rect 12341 7379 12407 7382
rect 12709 7442 12775 7445
rect 13261 7442 13327 7445
rect 12709 7440 13327 7442
rect 12709 7384 12714 7440
rect 12770 7384 13266 7440
rect 13322 7384 13327 7440
rect 12709 7382 13327 7384
rect 12709 7379 12775 7382
rect 13261 7379 13327 7382
rect 4061 7306 4127 7309
rect 5165 7306 5231 7309
rect 4061 7304 5231 7306
rect 4061 7248 4066 7304
rect 4122 7248 5170 7304
rect 5226 7248 5231 7304
rect 4061 7246 5231 7248
rect 4061 7243 4127 7246
rect 5165 7243 5231 7246
rect 7005 7306 7071 7309
rect 8385 7306 8451 7309
rect 15285 7306 15351 7309
rect 7005 7304 15351 7306
rect 7005 7248 7010 7304
rect 7066 7248 8390 7304
rect 8446 7248 15290 7304
rect 15346 7248 15351 7304
rect 7005 7246 15351 7248
rect 7005 7243 7071 7246
rect 8385 7243 8451 7246
rect 15285 7243 15351 7246
rect 7966 7108 7972 7172
rect 8036 7170 8042 7172
rect 8845 7170 8911 7173
rect 8036 7168 8911 7170
rect 8036 7112 8850 7168
rect 8906 7112 8911 7168
rect 8036 7110 8911 7112
rect 8036 7108 8042 7110
rect 8845 7107 8911 7110
rect 9029 7170 9095 7173
rect 12801 7170 12867 7173
rect 9029 7168 12867 7170
rect 9029 7112 9034 7168
rect 9090 7112 12806 7168
rect 12862 7112 12867 7168
rect 9029 7110 12867 7112
rect 9029 7107 9095 7110
rect 12801 7107 12867 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 5625 7034 5691 7037
rect 8109 7034 8175 7037
rect 8293 7036 8359 7037
rect 8293 7034 8340 7036
rect 5625 7032 5826 7034
rect 5625 6976 5630 7032
rect 5686 6976 5826 7032
rect 5625 6974 5826 6976
rect 5625 6971 5691 6974
rect 0 6898 800 6928
rect 5257 6898 5323 6901
rect 5766 6898 5826 6974
rect 8109 7032 8340 7034
rect 8109 6976 8114 7032
rect 8170 6976 8298 7032
rect 8109 6974 8340 6976
rect 8109 6971 8175 6974
rect 8293 6972 8340 6974
rect 8404 6972 8410 7036
rect 12709 7034 12775 7037
rect 9630 7032 12775 7034
rect 9630 6976 12714 7032
rect 12770 6976 12775 7032
rect 9630 6974 12775 6976
rect 8293 6971 8359 6972
rect 0 6808 858 6898
rect 5257 6896 5826 6898
rect 5257 6840 5262 6896
rect 5318 6840 5826 6896
rect 5257 6838 5826 6840
rect 5257 6835 5323 6838
rect 798 6765 858 6808
rect 798 6760 907 6765
rect 798 6704 846 6760
rect 902 6704 907 6760
rect 798 6702 907 6704
rect 841 6699 907 6702
rect 4337 6762 4403 6765
rect 5390 6762 5396 6764
rect 4337 6760 5396 6762
rect 4337 6704 4342 6760
rect 4398 6704 5396 6760
rect 4337 6702 5396 6704
rect 4337 6699 4403 6702
rect 5390 6700 5396 6702
rect 5460 6762 5466 6764
rect 5766 6762 5826 6838
rect 6821 6898 6887 6901
rect 9630 6898 9690 6974
rect 12709 6971 12775 6974
rect 6821 6896 9690 6898
rect 6821 6840 6826 6896
rect 6882 6840 9690 6896
rect 6821 6838 9690 6840
rect 11053 6898 11119 6901
rect 14917 6900 14983 6901
rect 11646 6898 11652 6900
rect 11053 6896 11652 6898
rect 11053 6840 11058 6896
rect 11114 6840 11652 6896
rect 11053 6838 11652 6840
rect 6821 6835 6887 6838
rect 11053 6835 11119 6838
rect 11646 6836 11652 6838
rect 11716 6836 11722 6900
rect 14917 6898 14964 6900
rect 14872 6896 14964 6898
rect 14872 6840 14922 6896
rect 14872 6838 14964 6840
rect 14917 6836 14964 6838
rect 15028 6836 15034 6900
rect 14917 6835 14983 6836
rect 10593 6762 10659 6765
rect 15745 6762 15811 6765
rect 5460 6702 5642 6762
rect 5766 6760 10659 6762
rect 5766 6704 10598 6760
rect 10654 6704 10659 6760
rect 5766 6702 10659 6704
rect 5460 6700 5466 6702
rect 5582 6626 5642 6702
rect 10593 6699 10659 6702
rect 12390 6760 15811 6762
rect 12390 6704 15750 6760
rect 15806 6704 15811 6760
rect 12390 6702 15811 6704
rect 12390 6626 12450 6702
rect 15745 6699 15811 6702
rect 5582 6566 12450 6626
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 3918 6428 3924 6492
rect 3988 6490 3994 6492
rect 4061 6490 4127 6493
rect 3988 6488 4127 6490
rect 3988 6432 4066 6488
rect 4122 6432 4127 6488
rect 3988 6430 4127 6432
rect 3988 6428 3994 6430
rect 4061 6427 4127 6430
rect 5901 6490 5967 6493
rect 7005 6490 7071 6493
rect 8201 6490 8267 6493
rect 5901 6488 8267 6490
rect 5901 6432 5906 6488
rect 5962 6432 7010 6488
rect 7066 6432 8206 6488
rect 8262 6432 8267 6488
rect 5901 6430 8267 6432
rect 5901 6427 5967 6430
rect 7005 6427 7071 6430
rect 8201 6427 8267 6430
rect 9949 6490 10015 6493
rect 13261 6490 13327 6493
rect 16849 6490 16915 6493
rect 9949 6488 13327 6490
rect 9949 6432 9954 6488
rect 10010 6432 13266 6488
rect 13322 6432 13327 6488
rect 9949 6430 13327 6432
rect 9949 6427 10015 6430
rect 13261 6427 13327 6430
rect 15748 6488 16915 6490
rect 15748 6432 16854 6488
rect 16910 6432 16915 6488
rect 15748 6430 16915 6432
rect 15748 6357 15808 6430
rect 16849 6427 16915 6430
rect 4705 6354 4771 6357
rect 5257 6354 5323 6357
rect 7833 6354 7899 6357
rect 4705 6352 7899 6354
rect 4705 6296 4710 6352
rect 4766 6296 5262 6352
rect 5318 6296 7838 6352
rect 7894 6296 7899 6352
rect 4705 6294 7899 6296
rect 4705 6291 4771 6294
rect 5257 6291 5323 6294
rect 7833 6291 7899 6294
rect 8937 6354 9003 6357
rect 10133 6354 10199 6357
rect 8937 6352 10199 6354
rect 8937 6296 8942 6352
rect 8998 6296 10138 6352
rect 10194 6296 10199 6352
rect 8937 6294 10199 6296
rect 8937 6291 9003 6294
rect 10133 6291 10199 6294
rect 10409 6354 10475 6357
rect 13670 6354 13676 6356
rect 10409 6352 13676 6354
rect 10409 6296 10414 6352
rect 10470 6296 13676 6352
rect 10409 6294 13676 6296
rect 10409 6291 10475 6294
rect 13670 6292 13676 6294
rect 13740 6354 13746 6356
rect 15745 6354 15811 6357
rect 16021 6356 16087 6357
rect 16021 6354 16068 6356
rect 13740 6352 15811 6354
rect 13740 6296 15750 6352
rect 15806 6296 15811 6352
rect 13740 6294 15811 6296
rect 15976 6352 16068 6354
rect 16132 6354 16138 6356
rect 16481 6354 16547 6357
rect 16132 6352 16547 6354
rect 15976 6296 16026 6352
rect 16132 6296 16486 6352
rect 16542 6296 16547 6352
rect 15976 6294 16068 6296
rect 13740 6292 13746 6294
rect 15745 6291 15811 6294
rect 16021 6292 16068 6294
rect 16132 6294 16547 6296
rect 16132 6292 16138 6294
rect 16021 6291 16087 6292
rect 16481 6291 16547 6294
rect 4705 6218 4771 6221
rect 6361 6218 6427 6221
rect 4705 6216 6427 6218
rect 4705 6160 4710 6216
rect 4766 6160 6366 6216
rect 6422 6160 6427 6216
rect 4705 6158 6427 6160
rect 4705 6155 4771 6158
rect 6361 6155 6427 6158
rect 9029 6218 9095 6221
rect 11513 6218 11579 6221
rect 12341 6218 12407 6221
rect 13721 6218 13787 6221
rect 9029 6216 11346 6218
rect 9029 6160 9034 6216
rect 9090 6160 11346 6216
rect 9029 6158 11346 6160
rect 9029 6155 9095 6158
rect 11286 6082 11346 6158
rect 11513 6216 13787 6218
rect 11513 6160 11518 6216
rect 11574 6160 12346 6216
rect 12402 6160 13726 6216
rect 13782 6160 13787 6216
rect 11513 6158 13787 6160
rect 11513 6155 11579 6158
rect 12341 6155 12407 6158
rect 13721 6155 13787 6158
rect 14089 6082 14155 6085
rect 11286 6080 14155 6082
rect 11286 6024 14094 6080
rect 14150 6024 14155 6080
rect 11286 6022 14155 6024
rect 14089 6019 14155 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 10317 5810 10383 5813
rect 10961 5810 11027 5813
rect 10317 5808 11027 5810
rect 10317 5752 10322 5808
rect 10378 5752 10966 5808
rect 11022 5752 11027 5808
rect 10317 5750 11027 5752
rect 10317 5747 10383 5750
rect 10961 5747 11027 5750
rect 11094 5748 11100 5812
rect 11164 5810 11170 5812
rect 13353 5810 13419 5813
rect 11164 5808 13419 5810
rect 11164 5752 13358 5808
rect 13414 5752 13419 5808
rect 11164 5750 13419 5752
rect 11164 5748 11170 5750
rect 13353 5747 13419 5750
rect 14181 5674 14247 5677
rect 9630 5672 14247 5674
rect 9630 5616 14186 5672
rect 14242 5616 14247 5672
rect 9630 5614 14247 5616
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 5441 5402 5507 5405
rect 6821 5402 6887 5405
rect 5441 5400 6887 5402
rect 5441 5344 5446 5400
rect 5502 5344 6826 5400
rect 6882 5344 6887 5400
rect 5441 5342 6887 5344
rect 5441 5339 5507 5342
rect 6821 5339 6887 5342
rect 9397 5402 9463 5405
rect 9630 5402 9690 5614
rect 14181 5611 14247 5614
rect 10133 5538 10199 5541
rect 13905 5538 13971 5541
rect 16205 5538 16271 5541
rect 10133 5536 16271 5538
rect 10133 5480 10138 5536
rect 10194 5480 13910 5536
rect 13966 5480 16210 5536
rect 16266 5480 16271 5536
rect 10133 5478 16271 5480
rect 10133 5475 10199 5478
rect 13905 5475 13971 5478
rect 16205 5475 16271 5478
rect 9397 5400 9690 5402
rect 9397 5344 9402 5400
rect 9458 5344 9690 5400
rect 9397 5342 9690 5344
rect 10041 5402 10107 5405
rect 10869 5402 10935 5405
rect 10041 5400 10935 5402
rect 10041 5344 10046 5400
rect 10102 5344 10874 5400
rect 10930 5344 10935 5400
rect 10041 5342 10935 5344
rect 9397 5339 9463 5342
rect 10041 5339 10107 5342
rect 10869 5339 10935 5342
rect 7373 5266 7439 5269
rect 15009 5266 15075 5269
rect 7373 5264 15075 5266
rect 7373 5208 7378 5264
rect 7434 5208 15014 5264
rect 15070 5208 15075 5264
rect 7373 5206 15075 5208
rect 7373 5203 7439 5206
rect 15009 5203 15075 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 10133 4858 10199 4861
rect 10910 4858 10916 4860
rect 10133 4856 10916 4858
rect 10133 4800 10138 4856
rect 10194 4800 10916 4856
rect 10133 4798 10916 4800
rect 10133 4795 10199 4798
rect 10910 4796 10916 4798
rect 10980 4858 10986 4860
rect 11513 4858 11579 4861
rect 14549 4858 14615 4861
rect 10980 4856 14615 4858
rect 10980 4800 11518 4856
rect 11574 4800 14554 4856
rect 14610 4800 14615 4856
rect 10980 4798 14615 4800
rect 10980 4796 10986 4798
rect 11513 4795 11579 4798
rect 14549 4795 14615 4798
rect 3325 4722 3391 4725
rect 6453 4722 6519 4725
rect 3325 4720 6519 4722
rect 3325 4664 3330 4720
rect 3386 4664 6458 4720
rect 6514 4664 6519 4720
rect 3325 4662 6519 4664
rect 3325 4659 3391 4662
rect 6453 4659 6519 4662
rect 10593 4722 10659 4725
rect 12433 4722 12499 4725
rect 15193 4724 15259 4725
rect 15142 4722 15148 4724
rect 10593 4720 12499 4722
rect 10593 4664 10598 4720
rect 10654 4664 12438 4720
rect 12494 4664 12499 4720
rect 10593 4662 12499 4664
rect 15102 4662 15148 4722
rect 15212 4720 15259 4724
rect 15254 4664 15259 4720
rect 10593 4659 10659 4662
rect 12433 4659 12499 4662
rect 15142 4660 15148 4662
rect 15212 4660 15259 4664
rect 15193 4659 15259 4660
rect 6269 4586 6335 4589
rect 8569 4586 8635 4589
rect 6269 4584 8635 4586
rect 6269 4528 6274 4584
rect 6330 4528 8574 4584
rect 8630 4528 8635 4584
rect 6269 4526 8635 4528
rect 6269 4523 6335 4526
rect 8569 4523 8635 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 10501 4042 10567 4045
rect 13854 4042 13860 4044
rect 10501 4040 13860 4042
rect 10501 3984 10506 4040
rect 10562 3984 13860 4040
rect 10501 3982 13860 3984
rect 10501 3979 10567 3982
rect 13854 3980 13860 3982
rect 13924 3980 13930 4044
rect 10501 3908 10567 3909
rect 10501 3906 10548 3908
rect 10456 3904 10548 3906
rect 10456 3848 10506 3904
rect 10456 3846 10548 3848
rect 10501 3844 10548 3846
rect 10612 3844 10618 3908
rect 10501 3843 10567 3844
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 8340 18260 8404 18324
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 8892 17580 8956 17644
rect 10364 17580 10428 17644
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 8156 17036 8220 17100
rect 11652 17096 11716 17100
rect 11652 17040 11702 17096
rect 11702 17040 11716 17096
rect 11652 17036 11716 17040
rect 17172 17036 17236 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 9076 16764 9140 16828
rect 9260 16628 9324 16692
rect 11468 16628 11532 16692
rect 9628 16492 9692 16556
rect 15884 16492 15948 16556
rect 5764 16416 5828 16420
rect 5764 16360 5778 16416
rect 5778 16360 5828 16416
rect 5764 16356 5828 16360
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 9812 16084 9876 16148
rect 3372 15948 3436 16012
rect 16804 15812 16868 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 2820 14860 2884 14924
rect 9996 14724 10060 14788
rect 15884 14724 15948 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 10732 14452 10796 14516
rect 8156 14180 8220 14244
rect 11652 14180 11716 14244
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 3740 14044 3804 14108
rect 8524 14044 8588 14108
rect 6132 13772 6196 13836
rect 10180 13772 10244 13836
rect 14964 13772 15028 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 5764 13500 5828 13564
rect 11652 13500 11716 13564
rect 7972 13364 8036 13428
rect 9628 13364 9692 13428
rect 3740 13092 3804 13156
rect 11100 13152 11164 13156
rect 11100 13096 11150 13152
rect 11150 13096 11164 13152
rect 11100 13092 11164 13096
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 3372 12820 3436 12884
rect 3924 12820 3988 12884
rect 7052 12820 7116 12884
rect 8340 12820 8404 12884
rect 13860 12820 13924 12884
rect 8340 12684 8404 12748
rect 17540 12684 17604 12748
rect 5396 12548 5460 12612
rect 9076 12608 9140 12612
rect 9076 12552 9090 12608
rect 9090 12552 9140 12608
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 2820 12336 2884 12340
rect 2820 12280 2870 12336
rect 2870 12280 2884 12336
rect 2820 12276 2884 12280
rect 7052 12276 7116 12340
rect 9076 12548 9140 12552
rect 9076 12412 9140 12476
rect 12388 12412 12452 12476
rect 11284 12276 11348 12340
rect 10180 12140 10244 12204
rect 4660 12004 4724 12068
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 9076 11792 9140 11796
rect 9076 11736 9090 11792
rect 9090 11736 9140 11792
rect 9076 11732 9140 11736
rect 5396 11596 5460 11660
rect 15884 11656 15948 11660
rect 15884 11600 15934 11656
rect 15934 11600 15948 11656
rect 15884 11596 15948 11600
rect 5396 11460 5460 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 9444 11324 9508 11388
rect 16068 11384 16132 11388
rect 16068 11328 16118 11384
rect 16118 11328 16132 11384
rect 16068 11324 16132 11328
rect 4660 11052 4724 11116
rect 8156 11188 8220 11252
rect 8892 11188 8956 11252
rect 10548 11112 10612 11116
rect 10548 11056 10598 11112
rect 10598 11056 10612 11112
rect 10548 11052 10612 11056
rect 9812 10916 9876 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 8524 10644 8588 10708
rect 5948 10508 6012 10572
rect 11652 10372 11716 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 9260 10236 9324 10300
rect 3740 10100 3804 10164
rect 9996 10100 10060 10164
rect 10916 10160 10980 10164
rect 10916 10104 10930 10160
rect 10930 10104 10980 10160
rect 10916 10100 10980 10104
rect 15148 10160 15212 10164
rect 15148 10104 15198 10160
rect 15198 10104 15212 10160
rect 15148 10100 15212 10104
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 6684 9752 6748 9756
rect 6684 9696 6698 9752
rect 6698 9696 6748 9752
rect 6684 9692 6748 9696
rect 11100 9692 11164 9756
rect 17172 9616 17236 9620
rect 17172 9560 17222 9616
rect 17222 9560 17236 9616
rect 17172 9556 17236 9560
rect 17540 9616 17604 9620
rect 17540 9560 17590 9616
rect 17590 9560 17604 9616
rect 17540 9556 17604 9560
rect 13676 9480 13740 9484
rect 13676 9424 13690 9480
rect 13690 9424 13740 9480
rect 13676 9420 13740 9424
rect 5396 9284 5460 9348
rect 9444 9284 9508 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 7052 9148 7116 9212
rect 11468 9148 11532 9212
rect 10364 8936 10428 8940
rect 10364 8880 10378 8936
rect 10378 8880 10428 8936
rect 10364 8876 10428 8880
rect 11100 8876 11164 8940
rect 5948 8740 6012 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 16068 8468 16132 8532
rect 6684 8332 6748 8396
rect 11284 8332 11348 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 10732 8256 10796 8260
rect 10732 8200 10746 8256
rect 10746 8200 10796 8256
rect 10732 8196 10796 8200
rect 16804 8256 16868 8260
rect 16804 8200 16854 8256
rect 16854 8200 16868 8256
rect 16804 8196 16868 8200
rect 12572 8060 12636 8124
rect 6132 7924 6196 7988
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 7972 7108 8036 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 8340 7032 8404 7036
rect 8340 6976 8354 7032
rect 8354 6976 8404 7032
rect 8340 6972 8404 6976
rect 5396 6700 5460 6764
rect 11652 6836 11716 6900
rect 14964 6896 15028 6900
rect 14964 6840 14978 6896
rect 14978 6840 15028 6896
rect 14964 6836 15028 6840
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 3924 6428 3988 6492
rect 13676 6292 13740 6356
rect 16068 6352 16132 6356
rect 16068 6296 16082 6352
rect 16082 6296 16132 6352
rect 16068 6292 16132 6296
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 11100 5748 11164 5812
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 10916 4796 10980 4860
rect 15148 4720 15212 4724
rect 15148 4664 15198 4720
rect 15198 4664 15212 4720
rect 15148 4660 15212 4664
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 13860 3980 13924 4044
rect 10548 3904 10612 3908
rect 10548 3848 10562 3904
rect 10562 3848 10612 3904
rect 10548 3844 10612 3848
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 19072 4528 19088
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 3371 16012 3437 16013
rect 3371 15948 3372 16012
rect 3436 15948 3437 16012
rect 3371 15947 3437 15948
rect 2819 14924 2885 14925
rect 2819 14860 2820 14924
rect 2884 14860 2885 14924
rect 2819 14859 2885 14860
rect 2822 12341 2882 14859
rect 3374 12885 3434 15947
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 3739 14108 3805 14109
rect 3739 14044 3740 14108
rect 3804 14044 3805 14108
rect 3739 14043 3805 14044
rect 3742 13157 3802 14043
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 3739 13156 3805 13157
rect 3739 13092 3740 13156
rect 3804 13092 3805 13156
rect 3739 13091 3805 13092
rect 3371 12884 3437 12885
rect 3371 12820 3372 12884
rect 3436 12820 3437 12884
rect 3371 12819 3437 12820
rect 2819 12340 2885 12341
rect 2819 12276 2820 12340
rect 2884 12276 2885 12340
rect 2819 12275 2885 12276
rect 3742 10165 3802 13091
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 3739 10164 3805 10165
rect 3739 10100 3740 10164
rect 3804 10100 3805 10164
rect 3739 10099 3805 10100
rect 3926 6493 3986 12819
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4868 18528 5188 19088
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 8339 18324 8405 18325
rect 8339 18260 8340 18324
rect 8404 18260 8405 18324
rect 8339 18259 8405 18260
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 8155 17100 8221 17101
rect 8155 17036 8156 17100
rect 8220 17036 8221 17100
rect 8155 17035 8221 17036
rect 5763 16420 5829 16421
rect 5763 16356 5764 16420
rect 5828 16356 5829 16420
rect 5763 16355 5829 16356
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 5766 13565 5826 16355
rect 8158 14245 8218 17035
rect 8155 14244 8221 14245
rect 8155 14180 8156 14244
rect 8220 14180 8221 14244
rect 8155 14179 8221 14180
rect 6131 13836 6197 13837
rect 6131 13772 6132 13836
rect 6196 13772 6197 13836
rect 6131 13771 6197 13772
rect 5763 13564 5829 13565
rect 5763 13500 5764 13564
rect 5828 13500 5829 13564
rect 5763 13499 5829 13500
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4659 12068 4725 12069
rect 4659 12004 4660 12068
rect 4724 12004 4725 12068
rect 4659 12003 4725 12004
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4662 11117 4722 12003
rect 4868 12000 5188 13024
rect 5395 12612 5461 12613
rect 5395 12548 5396 12612
rect 5460 12548 5461 12612
rect 5395 12547 5461 12548
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4659 11116 4725 11117
rect 4659 11052 4660 11116
rect 4724 11052 4725 11116
rect 4659 11051 4725 11052
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 3923 6492 3989 6493
rect 3923 6428 3924 6492
rect 3988 6428 3989 6492
rect 3923 6427 3989 6428
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 10912 5188 11936
rect 5398 11661 5458 12547
rect 5395 11660 5461 11661
rect 5395 11596 5396 11660
rect 5460 11596 5461 11660
rect 5395 11595 5461 11596
rect 5395 11524 5461 11525
rect 5395 11460 5396 11524
rect 5460 11460 5461 11524
rect 5395 11459 5461 11460
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 5398 9349 5458 11459
rect 5947 10572 6013 10573
rect 5947 10508 5948 10572
rect 6012 10508 6013 10572
rect 5947 10507 6013 10508
rect 5395 9348 5461 9349
rect 5395 9284 5396 9348
rect 5460 9284 5461 9348
rect 5395 9283 5461 9284
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 5398 6765 5458 9283
rect 5950 8805 6010 10507
rect 5947 8804 6013 8805
rect 5947 8740 5948 8804
rect 6012 8740 6013 8804
rect 5947 8739 6013 8740
rect 6134 7989 6194 13771
rect 7971 13428 8037 13429
rect 7971 13364 7972 13428
rect 8036 13364 8037 13428
rect 7971 13363 8037 13364
rect 7051 12884 7117 12885
rect 7051 12820 7052 12884
rect 7116 12820 7117 12884
rect 7051 12819 7117 12820
rect 7054 12341 7114 12819
rect 7051 12340 7117 12341
rect 7051 12276 7052 12340
rect 7116 12276 7117 12340
rect 7051 12275 7117 12276
rect 6683 9756 6749 9757
rect 6683 9692 6684 9756
rect 6748 9692 6749 9756
rect 6683 9691 6749 9692
rect 6686 8397 6746 9691
rect 7054 9213 7114 12275
rect 7051 9212 7117 9213
rect 7051 9148 7052 9212
rect 7116 9148 7117 9212
rect 7051 9147 7117 9148
rect 6683 8396 6749 8397
rect 6683 8332 6684 8396
rect 6748 8332 6749 8396
rect 6683 8331 6749 8332
rect 6131 7988 6197 7989
rect 6131 7924 6132 7988
rect 6196 7924 6197 7988
rect 6131 7923 6197 7924
rect 7974 7173 8034 13363
rect 8158 11253 8218 14179
rect 8342 12885 8402 18259
rect 8891 17644 8957 17645
rect 8891 17580 8892 17644
rect 8956 17580 8957 17644
rect 8891 17579 8957 17580
rect 10363 17644 10429 17645
rect 10363 17580 10364 17644
rect 10428 17580 10429 17644
rect 10363 17579 10429 17580
rect 8523 14108 8589 14109
rect 8523 14044 8524 14108
rect 8588 14044 8589 14108
rect 8523 14043 8589 14044
rect 8339 12884 8405 12885
rect 8339 12820 8340 12884
rect 8404 12820 8405 12884
rect 8339 12819 8405 12820
rect 8339 12748 8405 12749
rect 8339 12684 8340 12748
rect 8404 12684 8405 12748
rect 8339 12683 8405 12684
rect 8155 11252 8221 11253
rect 8155 11188 8156 11252
rect 8220 11188 8221 11252
rect 8155 11187 8221 11188
rect 7971 7172 8037 7173
rect 7971 7108 7972 7172
rect 8036 7108 8037 7172
rect 7971 7107 8037 7108
rect 8342 7037 8402 12683
rect 8526 10709 8586 14043
rect 8894 11253 8954 17579
rect 9075 16828 9141 16829
rect 9075 16764 9076 16828
rect 9140 16764 9141 16828
rect 9075 16763 9141 16764
rect 9078 12613 9138 16763
rect 9259 16692 9325 16693
rect 9259 16628 9260 16692
rect 9324 16628 9325 16692
rect 9259 16627 9325 16628
rect 9075 12612 9141 12613
rect 9075 12548 9076 12612
rect 9140 12548 9141 12612
rect 9075 12547 9141 12548
rect 9075 12476 9141 12477
rect 9075 12412 9076 12476
rect 9140 12412 9141 12476
rect 9075 12411 9141 12412
rect 9078 11797 9138 12411
rect 9075 11796 9141 11797
rect 9075 11732 9076 11796
rect 9140 11732 9141 11796
rect 9075 11731 9141 11732
rect 8891 11252 8957 11253
rect 8891 11188 8892 11252
rect 8956 11188 8957 11252
rect 8891 11187 8957 11188
rect 8523 10708 8589 10709
rect 8523 10644 8524 10708
rect 8588 10644 8589 10708
rect 8523 10643 8589 10644
rect 9262 10301 9322 16627
rect 9627 16556 9693 16557
rect 9627 16492 9628 16556
rect 9692 16492 9693 16556
rect 9627 16491 9693 16492
rect 9630 13429 9690 16491
rect 9811 16148 9877 16149
rect 9811 16084 9812 16148
rect 9876 16084 9877 16148
rect 9811 16083 9877 16084
rect 9627 13428 9693 13429
rect 9627 13364 9628 13428
rect 9692 13364 9693 13428
rect 9627 13363 9693 13364
rect 9443 11388 9509 11389
rect 9443 11324 9444 11388
rect 9508 11324 9509 11388
rect 9443 11323 9509 11324
rect 9259 10300 9325 10301
rect 9259 10236 9260 10300
rect 9324 10236 9325 10300
rect 9259 10235 9325 10236
rect 9446 9349 9506 11323
rect 9814 10981 9874 16083
rect 9995 14788 10061 14789
rect 9995 14724 9996 14788
rect 10060 14724 10061 14788
rect 9995 14723 10061 14724
rect 9811 10980 9877 10981
rect 9811 10916 9812 10980
rect 9876 10916 9877 10980
rect 9811 10915 9877 10916
rect 9998 10165 10058 14723
rect 10179 13836 10245 13837
rect 10179 13772 10180 13836
rect 10244 13772 10245 13836
rect 10179 13771 10245 13772
rect 10182 12205 10242 13771
rect 10179 12204 10245 12205
rect 10179 12140 10180 12204
rect 10244 12140 10245 12204
rect 10179 12139 10245 12140
rect 9995 10164 10061 10165
rect 9995 10100 9996 10164
rect 10060 10100 10061 10164
rect 9995 10099 10061 10100
rect 9443 9348 9509 9349
rect 9443 9284 9444 9348
rect 9508 9284 9509 9348
rect 9443 9283 9509 9284
rect 10366 8941 10426 17579
rect 11651 17100 11717 17101
rect 11651 17036 11652 17100
rect 11716 17036 11717 17100
rect 11651 17035 11717 17036
rect 17171 17100 17237 17101
rect 17171 17036 17172 17100
rect 17236 17036 17237 17100
rect 17171 17035 17237 17036
rect 11467 16692 11533 16693
rect 11467 16628 11468 16692
rect 11532 16628 11533 16692
rect 11467 16627 11533 16628
rect 10731 14516 10797 14517
rect 10731 14452 10732 14516
rect 10796 14452 10797 14516
rect 10731 14451 10797 14452
rect 10547 11116 10613 11117
rect 10547 11052 10548 11116
rect 10612 11052 10613 11116
rect 10547 11051 10613 11052
rect 10363 8940 10429 8941
rect 10363 8876 10364 8940
rect 10428 8876 10429 8940
rect 10363 8875 10429 8876
rect 8339 7036 8405 7037
rect 8339 6972 8340 7036
rect 8404 6972 8405 7036
rect 8339 6971 8405 6972
rect 5395 6764 5461 6765
rect 5395 6700 5396 6764
rect 5460 6700 5461 6764
rect 5395 6699 5461 6700
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 10550 3909 10610 11051
rect 10734 8261 10794 14451
rect 11099 13156 11165 13157
rect 11099 13092 11100 13156
rect 11164 13092 11165 13156
rect 11099 13091 11165 13092
rect 10915 10164 10981 10165
rect 10915 10100 10916 10164
rect 10980 10100 10981 10164
rect 10915 10099 10981 10100
rect 10731 8260 10797 8261
rect 10731 8196 10732 8260
rect 10796 8196 10797 8260
rect 10731 8195 10797 8196
rect 10918 4861 10978 10099
rect 11102 9757 11162 13091
rect 11283 12340 11349 12341
rect 11283 12276 11284 12340
rect 11348 12276 11349 12340
rect 11283 12275 11349 12276
rect 11099 9756 11165 9757
rect 11099 9692 11100 9756
rect 11164 9692 11165 9756
rect 11099 9691 11165 9692
rect 11099 8940 11165 8941
rect 11099 8876 11100 8940
rect 11164 8876 11165 8940
rect 11099 8875 11165 8876
rect 11102 5813 11162 8875
rect 11286 8397 11346 12275
rect 11470 9213 11530 16627
rect 11654 14245 11714 17035
rect 15883 16556 15949 16557
rect 15883 16492 15884 16556
rect 15948 16492 15949 16556
rect 15883 16491 15949 16492
rect 15886 14789 15946 16491
rect 16803 15876 16869 15877
rect 16803 15812 16804 15876
rect 16868 15812 16869 15876
rect 16803 15811 16869 15812
rect 15883 14788 15949 14789
rect 15883 14724 15884 14788
rect 15948 14724 15949 14788
rect 15883 14723 15949 14724
rect 11651 14244 11717 14245
rect 11651 14180 11652 14244
rect 11716 14180 11717 14244
rect 11651 14179 11717 14180
rect 14963 13836 15029 13837
rect 14963 13772 14964 13836
rect 15028 13772 15029 13836
rect 14963 13771 15029 13772
rect 11651 13564 11717 13565
rect 11651 13500 11652 13564
rect 11716 13500 11717 13564
rect 11651 13499 11717 13500
rect 11654 10437 11714 13499
rect 13859 12884 13925 12885
rect 13859 12820 13860 12884
rect 13924 12820 13925 12884
rect 13859 12819 13925 12820
rect 12387 12476 12453 12477
rect 12387 12412 12388 12476
rect 12452 12450 12453 12476
rect 12452 12412 12634 12450
rect 12387 12411 12634 12412
rect 12390 12390 12634 12411
rect 11651 10436 11717 10437
rect 11651 10372 11652 10436
rect 11716 10372 11717 10436
rect 11651 10371 11717 10372
rect 11467 9212 11533 9213
rect 11467 9148 11468 9212
rect 11532 9148 11533 9212
rect 11467 9147 11533 9148
rect 11283 8396 11349 8397
rect 11283 8332 11284 8396
rect 11348 8332 11349 8396
rect 11283 8331 11349 8332
rect 11654 6901 11714 10371
rect 12574 8125 12634 12390
rect 13675 9484 13741 9485
rect 13675 9420 13676 9484
rect 13740 9420 13741 9484
rect 13675 9419 13741 9420
rect 12571 8124 12637 8125
rect 12571 8060 12572 8124
rect 12636 8060 12637 8124
rect 12571 8059 12637 8060
rect 11651 6900 11717 6901
rect 11651 6836 11652 6900
rect 11716 6836 11717 6900
rect 11651 6835 11717 6836
rect 13678 6357 13738 9419
rect 13675 6356 13741 6357
rect 13675 6292 13676 6356
rect 13740 6292 13741 6356
rect 13675 6291 13741 6292
rect 11099 5812 11165 5813
rect 11099 5748 11100 5812
rect 11164 5748 11165 5812
rect 11099 5747 11165 5748
rect 10915 4860 10981 4861
rect 10915 4796 10916 4860
rect 10980 4796 10981 4860
rect 10915 4795 10981 4796
rect 13862 4045 13922 12819
rect 14966 6901 15026 13771
rect 15886 11661 15946 14723
rect 15883 11660 15949 11661
rect 15883 11596 15884 11660
rect 15948 11596 15949 11660
rect 15883 11595 15949 11596
rect 16067 11388 16133 11389
rect 16067 11324 16068 11388
rect 16132 11324 16133 11388
rect 16067 11323 16133 11324
rect 15147 10164 15213 10165
rect 15147 10100 15148 10164
rect 15212 10100 15213 10164
rect 15147 10099 15213 10100
rect 14963 6900 15029 6901
rect 14963 6836 14964 6900
rect 15028 6836 15029 6900
rect 14963 6835 15029 6836
rect 15150 4725 15210 10099
rect 16070 8533 16130 11323
rect 16067 8532 16133 8533
rect 16067 8468 16068 8532
rect 16132 8468 16133 8532
rect 16067 8467 16133 8468
rect 16070 6357 16130 8467
rect 16806 8261 16866 15811
rect 17174 9621 17234 17035
rect 17539 12748 17605 12749
rect 17539 12684 17540 12748
rect 17604 12684 17605 12748
rect 17539 12683 17605 12684
rect 17542 9621 17602 12683
rect 17171 9620 17237 9621
rect 17171 9556 17172 9620
rect 17236 9556 17237 9620
rect 17171 9555 17237 9556
rect 17539 9620 17605 9621
rect 17539 9556 17540 9620
rect 17604 9556 17605 9620
rect 17539 9555 17605 9556
rect 16803 8260 16869 8261
rect 16803 8196 16804 8260
rect 16868 8196 16869 8260
rect 16803 8195 16869 8196
rect 16067 6356 16133 6357
rect 16067 6292 16068 6356
rect 16132 6292 16133 6356
rect 16067 6291 16133 6292
rect 15147 4724 15213 4725
rect 15147 4660 15148 4724
rect 15212 4660 15213 4724
rect 15147 4659 15213 4660
rect 13859 4044 13925 4045
rect 13859 3980 13860 4044
rect 13924 3980 13925 4044
rect 13859 3979 13925 3980
rect 10547 3908 10613 3909
rect 10547 3844 10548 3908
rect 10612 3844 10613 3908
rect 10547 3843 10613 3844
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _387_
timestamp 0
transform 1 0 15640 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 0
transform -1 0 13984 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 0
transform -1 0 16468 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 0
transform 1 0 4324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp 0
transform -1 0 16468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 0
transform 1 0 10948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 0
transform -1 0 2392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 0
transform 1 0 17756 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _395_
timestamp 0
transform 1 0 15548 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__and2b_2  _396_
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _397_
timestamp 0
transform -1 0 4968 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _398_
timestamp 0
transform -1 0 13248 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_2  _399_
timestamp 0
transform -1 0 17480 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _400_
timestamp 0
transform -1 0 8464 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _401_
timestamp 0
transform -1 0 9016 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_2  _402_
timestamp 0
transform -1 0 13064 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _403_
timestamp 0
transform 1 0 3864 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _404_
timestamp 0
transform 1 0 15732 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _405_
timestamp 0
transform 1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _406_
timestamp 0
transform -1 0 15272 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _407_
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _408_
timestamp 0
transform -1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _409_
timestamp 0
transform -1 0 14536 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _410_
timestamp 0
transform 1 0 3956 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _411_
timestamp 0
transform 1 0 16836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _412_
timestamp 0
transform 1 0 15640 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _413_
timestamp 0
transform -1 0 3680 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _414_
timestamp 0
transform -1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _415_
timestamp 0
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _416_
timestamp 0
transform 1 0 4232 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _417_
timestamp 0
transform -1 0 12052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _418_
timestamp 0
transform 1 0 3220 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _419_
timestamp 0
transform 1 0 12052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _420_
timestamp 0
transform 1 0 12144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _421_
timestamp 0
transform -1 0 15640 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _422_
timestamp 0
transform -1 0 5888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _423_
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _424_
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_2  _425_
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _426_
timestamp 0
transform 1 0 13064 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _427_
timestamp 0
transform 1 0 8740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _428_
timestamp 0
transform 1 0 12696 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _429_
timestamp 0
transform 1 0 14536 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _430_
timestamp 0
transform -1 0 3680 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _431_
timestamp 0
transform -1 0 12880 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _432_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 0
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _434_
timestamp 0
transform -1 0 6164 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _435_
timestamp 0
transform 1 0 2668 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _436_
timestamp 0
transform -1 0 13892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _437_
timestamp 0
transform -1 0 17480 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _438_
timestamp 0
transform 1 0 6256 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _439_
timestamp 0
transform 1 0 15364 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _440_
timestamp 0
transform -1 0 7820 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _441_
timestamp 0
transform -1 0 17664 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_1  _442_
timestamp 0
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _443_
timestamp 0
transform -1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _444_
timestamp 0
transform -1 0 13616 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _446_
timestamp 0
transform -1 0 13800 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _447_
timestamp 0
transform 1 0 3496 0 -1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _448_
timestamp 0
transform -1 0 12788 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _449_
timestamp 0
transform -1 0 13248 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _450_
timestamp 0
transform 1 0 4876 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_2  _451_
timestamp 0
transform 1 0 14536 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _452_
timestamp 0
transform 1 0 4968 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _453_
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _454_
timestamp 0
transform 1 0 7544 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _455_
timestamp 0
transform 1 0 8096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _456_
timestamp 0
transform -1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _457_
timestamp 0
transform -1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _458_
timestamp 0
transform -1 0 4232 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _459_
timestamp 0
transform -1 0 3680 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_2  _460_
timestamp 0
transform -1 0 9660 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_2  _461_
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _462_
timestamp 0
transform -1 0 8832 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _463_
timestamp 0
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _464_
timestamp 0
transform -1 0 17296 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _465_
timestamp 0
transform -1 0 17664 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _466_
timestamp 0
transform -1 0 14996 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _467_
timestamp 0
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _468_
timestamp 0
transform -1 0 13524 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _469_
timestamp 0
transform -1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _470_
timestamp 0
transform 1 0 14352 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _471_
timestamp 0
transform 1 0 4784 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _472_
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _473_
timestamp 0
transform 1 0 7820 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _474_
timestamp 0
transform 1 0 17296 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _475_
timestamp 0
transform -1 0 4416 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _476_
timestamp 0
transform 1 0 6808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32oi_1  _477_
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _478_
timestamp 0
transform -1 0 8924 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _479_
timestamp 0
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _480_
timestamp 0
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _481_
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _482_
timestamp 0
transform 1 0 4968 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _483_
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _484_
timestamp 0
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _485_
timestamp 0
transform 1 0 4508 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _486_
timestamp 0
transform 1 0 15916 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _487_
timestamp 0
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _488_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _489_
timestamp 0
transform 1 0 5428 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _490_
timestamp 0
transform 1 0 7912 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _491_
timestamp 0
transform 1 0 10396 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _492_
timestamp 0
transform -1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _493_
timestamp 0
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _494_
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _495_
timestamp 0
transform -1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _496_
timestamp 0
transform 1 0 10396 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _497_
timestamp 0
transform -1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _498_
timestamp 0
transform -1 0 10120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _499_
timestamp 0
transform -1 0 9752 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _500_
timestamp 0
transform -1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _501_
timestamp 0
transform -1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _502_
timestamp 0
transform 1 0 7176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _503_
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _504_
timestamp 0
transform 1 0 6440 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _505_
timestamp 0
transform 1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _506_
timestamp 0
transform -1 0 10672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _507_
timestamp 0
transform 1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _508_
timestamp 0
transform 1 0 3864 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _509_
timestamp 0
transform 1 0 6624 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _510_
timestamp 0
transform -1 0 7176 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _511_
timestamp 0
transform -1 0 8832 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _512_
timestamp 0
transform -1 0 9292 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _513_
timestamp 0
transform 1 0 9108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _514_
timestamp 0
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _515_
timestamp 0
transform -1 0 16008 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _516_
timestamp 0
transform 1 0 13616 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _517_
timestamp 0
transform 1 0 13984 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _518_
timestamp 0
transform -1 0 7728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _519_
timestamp 0
transform -1 0 10304 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _520_
timestamp 0
transform -1 0 14168 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _521_
timestamp 0
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _522_
timestamp 0
transform 1 0 15640 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _523_
timestamp 0
transform -1 0 15456 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _524_
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _525_
timestamp 0
transform -1 0 9108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _526_
timestamp 0
transform -1 0 11960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _527_
timestamp 0
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _528_
timestamp 0
transform 1 0 12420 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _529_
timestamp 0
transform -1 0 17480 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _530_
timestamp 0
transform 1 0 7176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _531_
timestamp 0
transform 1 0 17296 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _532_
timestamp 0
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _533_
timestamp 0
transform -1 0 17112 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _534_
timestamp 0
transform -1 0 17296 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _535_
timestamp 0
transform -1 0 14904 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _536_
timestamp 0
transform -1 0 15916 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _537_
timestamp 0
transform -1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _538_
timestamp 0
transform -1 0 15456 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _539_
timestamp 0
transform 1 0 14904 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _540_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _541_
timestamp 0
transform -1 0 8832 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _542_
timestamp 0
transform 1 0 11868 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _543_
timestamp 0
transform 1 0 11316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _544_
timestamp 0
transform -1 0 15088 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _545_
timestamp 0
transform -1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _546_
timestamp 0
transform -1 0 5152 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _547_
timestamp 0
transform 1 0 6716 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _548_
timestamp 0
transform -1 0 7636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _549_
timestamp 0
transform 1 0 14168 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _550_
timestamp 0
transform -1 0 12788 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _551_
timestamp 0
transform 1 0 12788 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _552_
timestamp 0
transform 1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _553_
timestamp 0
transform 1 0 7176 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _554_
timestamp 0
transform 1 0 11960 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _555_
timestamp 0
transform -1 0 12328 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _556_
timestamp 0
transform 1 0 13892 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _557_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _558_
timestamp 0
transform 1 0 15916 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _559_
timestamp 0
transform 1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _560_
timestamp 0
transform -1 0 13984 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _561_
timestamp 0
transform 1 0 12512 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _562_
timestamp 0
transform 1 0 13248 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _563_
timestamp 0
transform -1 0 7820 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _564_
timestamp 0
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _565_
timestamp 0
transform 1 0 6900 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _566_
timestamp 0
transform -1 0 10856 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _567_
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _568_
timestamp 0
transform -1 0 15364 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _569_
timestamp 0
transform -1 0 13340 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _570_
timestamp 0
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _571_
timestamp 0
transform 1 0 12052 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _572_
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _573_
timestamp 0
transform 1 0 7176 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _574_
timestamp 0
transform -1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _575_
timestamp 0
transform -1 0 12696 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _576_
timestamp 0
transform -1 0 10120 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _577_
timestamp 0
transform -1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _578_
timestamp 0
transform 1 0 10028 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _579_
timestamp 0
transform -1 0 5244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _580_
timestamp 0
transform 1 0 6532 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _581_
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _582_
timestamp 0
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _583_
timestamp 0
transform -1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _584_
timestamp 0
transform 1 0 12788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _585_
timestamp 0
transform -1 0 12328 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _586_
timestamp 0
transform 1 0 10120 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _587_
timestamp 0
transform 1 0 11040 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _588_
timestamp 0
transform -1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _589_
timestamp 0
transform 1 0 5612 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _590_
timestamp 0
transform -1 0 9752 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _591_
timestamp 0
transform 1 0 9016 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _592_
timestamp 0
transform -1 0 7452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _593_
timestamp 0
transform 1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _594_
timestamp 0
transform -1 0 9752 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _595_
timestamp 0
transform 1 0 11500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _596_
timestamp 0
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _597_
timestamp 0
transform -1 0 4140 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _598_
timestamp 0
transform 1 0 9292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _599_
timestamp 0
transform -1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _600_
timestamp 0
transform -1 0 9844 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _601_
timestamp 0
transform 1 0 9476 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _602_
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _603_
timestamp 0
transform 1 0 11316 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _604_
timestamp 0
transform 1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _605_
timestamp 0
transform -1 0 7728 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _606_
timestamp 0
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _607_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _608_
timestamp 0
transform 1 0 6164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _609_
timestamp 0
transform -1 0 7268 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _610_
timestamp 0
transform 1 0 5704 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _611_
timestamp 0
transform -1 0 4048 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_4  _612_
timestamp 0
transform -1 0 5612 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__a2bb2o_1  _613_
timestamp 0
transform 1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _614_
timestamp 0
transform 1 0 2392 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _615_
timestamp 0
transform -1 0 4784 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _616_
timestamp 0
transform 1 0 4600 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _617_
timestamp 0
transform 1 0 6348 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _618_
timestamp 0
transform 1 0 5888 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _619_
timestamp 0
transform -1 0 4140 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _620_
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _621_
timestamp 0
transform 1 0 3036 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _622_
timestamp 0
transform 1 0 2760 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _623_
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _624_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _625_
timestamp 0
transform 1 0 2392 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _626_
timestamp 0
transform 1 0 2024 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _627_
timestamp 0
transform -1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _628_
timestamp 0
transform 1 0 7176 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _629_
timestamp 0
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _630_
timestamp 0
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _631_
timestamp 0
transform -1 0 15640 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _632_
timestamp 0
transform -1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _633_
timestamp 0
transform -1 0 2944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _634_
timestamp 0
transform 1 0 6900 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _635_
timestamp 0
transform -1 0 8740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _636_
timestamp 0
transform 1 0 9476 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _637_
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _638_
timestamp 0
transform -1 0 8832 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _639_
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _640_
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _641_
timestamp 0
transform -1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _642_
timestamp 0
transform 1 0 9384 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _643_
timestamp 0
transform 1 0 8280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _644_
timestamp 0
transform 1 0 8096 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _645_
timestamp 0
transform 1 0 7636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _646_
timestamp 0
transform 1 0 9752 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _647_
timestamp 0
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _648_
timestamp 0
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _649_
timestamp 0
transform -1 0 8096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _650_
timestamp 0
transform -1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _651_
timestamp 0
transform -1 0 4876 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _652_
timestamp 0
transform 1 0 5060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _653_
timestamp 0
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _654_
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _655_
timestamp 0
transform 1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _656_
timestamp 0
transform -1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _657_
timestamp 0
transform 1 0 11592 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _658_
timestamp 0
transform -1 0 9476 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _659_
timestamp 0
transform -1 0 4600 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _660_
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _661_
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _662_
timestamp 0
transform 1 0 14168 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _663_
timestamp 0
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _664_
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _665_
timestamp 0
transform 1 0 2300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _666_
timestamp 0
transform -1 0 2852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _667_
timestamp 0
transform -1 0 2484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _668_
timestamp 0
transform 1 0 2116 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _669_
timestamp 0
transform -1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _670_
timestamp 0
transform 1 0 1472 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _671_
timestamp 0
transform 1 0 13340 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _672_
timestamp 0
transform 1 0 10948 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _673_
timestamp 0
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _674_
timestamp 0
transform -1 0 10764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _675_
timestamp 0
transform -1 0 10764 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _676_
timestamp 0
transform 1 0 10304 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _677_
timestamp 0
transform 1 0 7452 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _678_
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _679_
timestamp 0
transform -1 0 6072 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _680_
timestamp 0
transform 1 0 6532 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _681_
timestamp 0
transform -1 0 6440 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _682_
timestamp 0
transform -1 0 7084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _683_
timestamp 0
transform 1 0 5612 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _684_
timestamp 0
transform -1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _685_
timestamp 0
transform -1 0 2116 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _686_
timestamp 0
transform 1 0 1472 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _687_
timestamp 0
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _688_
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _689_
timestamp 0
transform 1 0 7176 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _690_
timestamp 0
transform 1 0 8188 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _691_
timestamp 0
transform -1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _692_
timestamp 0
transform 1 0 7084 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _693_
timestamp 0
transform 1 0 7636 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _694_
timestamp 0
transform -1 0 8096 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _695_
timestamp 0
transform -1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _696_
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _697_
timestamp 0
transform -1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _698_
timestamp 0
transform -1 0 10488 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _699_
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _700_
timestamp 0
transform 1 0 11040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _701_
timestamp 0
transform -1 0 11040 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _702_
timestamp 0
transform 1 0 10028 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _703_
timestamp 0
transform 1 0 9384 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _704_
timestamp 0
transform 1 0 3312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _705_
timestamp 0
transform -1 0 4600 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _706_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _707_
timestamp 0
transform 1 0 5244 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _708_
timestamp 0
transform 1 0 4416 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _709_
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _710_
timestamp 0
transform 1 0 2392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _711_
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _712_
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _713_
timestamp 0
transform 1 0 5152 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _714_
timestamp 0
transform 1 0 4416 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _715_
timestamp 0
transform -1 0 3404 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _716_
timestamp 0
transform 1 0 1472 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _717_
timestamp 0
transform 1 0 16008 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _718_
timestamp 0
transform -1 0 15272 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _719_
timestamp 0
transform 1 0 15088 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _720_
timestamp 0
transform 1 0 14536 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _721_
timestamp 0
transform 1 0 9568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _722_
timestamp 0
transform 1 0 15272 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _723_
timestamp 0
transform 1 0 11040 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _724_
timestamp 0
transform -1 0 14444 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _725_
timestamp 0
transform 1 0 13248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _726_
timestamp 0
transform 1 0 13156 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _727_
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _728_
timestamp 0
transform -1 0 17940 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _729_
timestamp 0
transform -1 0 12328 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _730_
timestamp 0
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _731_
timestamp 0
transform 1 0 13432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _732_
timestamp 0
transform -1 0 13064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _733_
timestamp 0
transform -1 0 13340 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _734_
timestamp 0
transform 1 0 12880 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _735_
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _736_
timestamp 0
transform -1 0 12052 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _737_
timestamp 0
transform 1 0 10396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _738_
timestamp 0
transform 1 0 10856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _739_
timestamp 0
transform -1 0 10856 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _740_
timestamp 0
transform 1 0 9660 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _741_
timestamp 0
transform 1 0 9752 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _742_
timestamp 0
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _743_
timestamp 0
transform 1 0 10120 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _744_
timestamp 0
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _745_
timestamp 0
transform 1 0 17388 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _746_
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _747_
timestamp 0
transform 1 0 9752 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _748_
timestamp 0
transform 1 0 9476 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _749_
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _750_
timestamp 0
transform 1 0 1472 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _751_
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _752_
timestamp 0
transform 1 0 2392 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _753_
timestamp 0
transform 1 0 2852 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _754_
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _755_
timestamp 0
transform 1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _756_
timestamp 0
transform 1 0 2392 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _757_
timestamp 0
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _758_
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _759_
timestamp 0
transform 1 0 2576 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _760_
timestamp 0
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _761_
timestamp 0
transform 1 0 1472 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _762_
timestamp 0
transform -1 0 6716 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _763_
timestamp 0
transform 1 0 4600 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _764_
timestamp 0
transform -1 0 5336 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _765_
timestamp 0
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _766_
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _767_
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _768_
timestamp 0
transform 1 0 1656 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _769_
timestamp 0
transform 1 0 1472 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _770_
timestamp 0
transform 1 0 3036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _771_
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _772_
timestamp 0
transform 1 0 1472 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _773_
timestamp 0
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _774_
timestamp 0
transform -1 0 16284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _775_
timestamp 0
transform -1 0 14536 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _776_
timestamp 0
transform 1 0 14904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _777_
timestamp 0
transform 1 0 14352 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _778_
timestamp 0
transform 1 0 15088 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _779_
timestamp 0
transform 1 0 12604 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _780_
timestamp 0
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _781_
timestamp 0
transform -1 0 13248 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _782_
timestamp 0
transform 1 0 12328 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _783_
timestamp 0
transform 1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _784_
timestamp 0
transform 1 0 17848 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _785_
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _786_
timestamp 0
transform -1 0 17572 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _787_
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _788_
timestamp 0
transform 1 0 14628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _789_
timestamp 0
transform -1 0 13984 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _790_
timestamp 0
transform 1 0 15916 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _791_
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _792_
timestamp 0
transform 1 0 16376 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _793_
timestamp 0
transform 1 0 16008 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _794_
timestamp 0
transform 1 0 15456 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _795_
timestamp 0
transform 1 0 15916 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _796_
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _797_
timestamp 0
transform -1 0 15088 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 17112 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform 1 0 16376 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform -1 0 16560 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 0
transform -1 0 5612 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 0
transform -1 0 2760 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 0
transform -1 0 8648 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 0
transform 1 0 9108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 0
transform -1 0 16744 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 0
transform -1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 0
transform -1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 0
transform -1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 0
transform -1 0 15824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 0
transform -1 0 15088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout29
timestamp 0
transform -1 0 4692 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout30
timestamp 0
transform -1 0 6256 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 0
transform -1 0 5888 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout32
timestamp 0
transform -1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp 0
transform -1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 0
transform 1 0 15640 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 0
transform -1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout36
timestamp 0
transform 1 0 11776 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 0
transform -1 0 3864 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 0
transform -1 0 9108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 0
transform 1 0 14536 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout40
timestamp 0
transform -1 0 16008 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 0
transform -1 0 9752 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp 0
transform -1 0 9476 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 0
transform 1 0 17572 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 0
transform -1 0 10396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 0
transform -1 0 5244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 0
transform 1 0 10396 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 0
transform -1 0 9936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 0
transform -1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 0
transform -1 0 14720 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout50
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 0
transform -1 0 6348 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 0
transform 1 0 7084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout53
timestamp 0
transform -1 0 5612 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout54
timestamp 0
transform 1 0 10120 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout55
timestamp 0
transform -1 0 11132 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 0
transform 1 0 16468 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp 0
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 0
transform -1 0 16008 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout59
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout60
timestamp 0
transform -1 0 17848 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_8  fanout61
timestamp 0
transform -1 0 8280 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 0
transform -1 0 8648 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout63
timestamp 0
transform -1 0 6808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout64
timestamp 0
transform -1 0 8096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp 0
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout66
timestamp 0
transform 1 0 16836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout67
timestamp 0
transform 1 0 15456 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout68
timestamp 0
transform -1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout69
timestamp 0
transform -1 0 18032 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout70
timestamp 0
transform -1 0 7912 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout71
timestamp 0
transform -1 0 8004 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 0
transform -1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 0
transform -1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp 0
transform 1 0 16008 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout75
timestamp 0
transform -1 0 7176 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout76
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp 0
transform 1 0 16928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 0
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout79
timestamp 0
transform -1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91
timestamp 0
transform 1 0 9476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 0
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 0
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 0
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 0
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 0
transform 1 0 18124 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 0
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 0
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 0
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_185
timestamp 0
transform 1 0 18124 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_23
timestamp 0
transform 1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_48
timestamp 0
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_79
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 0
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 0
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 0
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_119
timestamp 0
transform 1 0 12052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_130
timestamp 0
transform 1 0 13064 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 0
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_143
timestamp 0
transform 1 0 14260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_147
timestamp 0
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 0
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_163
timestamp 0
transform 1 0 16100 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_174
timestamp 0
transform 1 0 17112 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp 0
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 0
transform 1 0 6532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_78
timestamp 0
transform 1 0 8280 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_122
timestamp 0
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 0
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 0
transform 1 0 14352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_156
timestamp 0
transform 1 0 15456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_178
timestamp 0
transform 1 0 17480 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 0
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_65
timestamp 0
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp 0
transform 1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp 0
transform 1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 0
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_130
timestamp 0
transform 1 0 13064 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 0
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_178
timestamp 0
transform 1 0 17480 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 0
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_20
timestamp 0
transform 1 0 2944 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_36
timestamp 0
transform 1 0 4416 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_47
timestamp 0
transform 1 0 5428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_54
timestamp 0
transform 1 0 6072 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_66
timestamp 0
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_78
timestamp 0
transform 1 0 8280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_91
timestamp 0
transform 1 0 9476 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_99
timestamp 0
transform 1 0 10212 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_110
timestamp 0
transform 1 0 11224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_118
timestamp 0
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 0
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp 0
transform 1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 0
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_178
timestamp 0
transform 1 0 17480 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 0
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_33
timestamp 0
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_45
timestamp 0
transform 1 0 5244 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_95
timestamp 0
transform 1 0 9844 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 0
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_118
timestamp 0
transform 1 0 11960 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_140
timestamp 0
transform 1 0 13984 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_152
timestamp 0
transform 1 0 15088 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_183
timestamp 0
transform 1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_7
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_18
timestamp 0
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 0
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 0
transform 1 0 5796 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_59
timestamp 0
transform 1 0 6532 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 0
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 0
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_115
timestamp 0
transform 1 0 11684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_127
timestamp 0
transform 1 0 12788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_147
timestamp 0
transform 1 0 14628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_162
timestamp 0
transform 1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_166
timestamp 0
transform 1 0 16376 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_174
timestamp 0
transform 1 0 17112 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_13
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_25
timestamp 0
transform 1 0 3404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_29
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 0
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_131
timestamp 0
transform 1 0 13156 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_143
timestamp 0
transform 1 0 14260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_152
timestamp 0
transform 1 0 15088 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_156
timestamp 0
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 0
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 0
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 0
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_40
timestamp 0
transform 1 0 4784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 0
transform 1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_72
timestamp 0
transform 1 0 7728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 0
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_100
timestamp 0
transform 1 0 10304 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_108
timestamp 0
transform 1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_161
timestamp 0
transform 1 0 15916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_169
timestamp 0
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_179
timestamp 0
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_11
timestamp 0
transform 1 0 2116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_23
timestamp 0
transform 1 0 3220 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 0
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 0
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_80
timestamp 0
transform 1 0 8464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_104
timestamp 0
transform 1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_121
timestamp 0
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_129
timestamp 0
transform 1 0 12972 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 0
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_145
timestamp 0
transform 1 0 14444 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_158
timestamp 0
transform 1 0 15640 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_185
timestamp 0
transform 1 0 18124 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_36
timestamp 0
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 0
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 0
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 0
transform 1 0 9200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 0
transform 1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_118
timestamp 0
transform 1 0 11960 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_130
timestamp 0
transform 1 0 13064 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 0
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 0
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_183
timestamp 0
transform 1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_32
timestamp 0
transform 1 0 4048 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_49
timestamp 0
transform 1 0 5612 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_64
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_76
timestamp 0
transform 1 0 8096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_100
timestamp 0
transform 1 0 10304 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_121
timestamp 0
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_145
timestamp 0
transform 1 0 14444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_157
timestamp 0
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 0
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 0
transform 1 0 18032 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_7
timestamp 0
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 0
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_36
timestamp 0
transform 1 0 4416 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_44
timestamp 0
transform 1 0 5152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_73
timestamp 0
transform 1 0 7820 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 0
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_89
timestamp 0
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_108
timestamp 0
transform 1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_114
timestamp 0
transform 1 0 11592 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_160
timestamp 0
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_184
timestamp 0
transform 1 0 18032 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_23
timestamp 0
transform 1 0 3220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_38
timestamp 0
transform 1 0 4600 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 0
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_65
timestamp 0
transform 1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_85
timestamp 0
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_97
timestamp 0
transform 1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 0
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_122
timestamp 0
transform 1 0 12328 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_134
timestamp 0
transform 1 0 13432 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_138
timestamp 0
transform 1 0 13800 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 0
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 0
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 0
transform 1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 0
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_35
timestamp 0
transform 1 0 4324 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_61
timestamp 0
transform 1 0 6716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_75
timestamp 0
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 0
transform 1 0 9568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_96
timestamp 0
transform 1 0 9936 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_104
timestamp 0
transform 1 0 10672 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_116
timestamp 0
transform 1 0 11776 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 0
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 0
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_160
timestamp 0
transform 1 0 15824 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_21
timestamp 0
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_29
timestamp 0
transform 1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 0
transform 1 0 4600 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_61
timestamp 0
transform 1 0 6716 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_71
timestamp 0
transform 1 0 7636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_83
timestamp 0
transform 1 0 8740 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_91
timestamp 0
transform 1 0 9476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 0
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 0
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_117
timestamp 0
transform 1 0 11868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_138
timestamp 0
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_150
timestamp 0
transform 1 0 14904 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 0
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 0
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_182
timestamp 0
transform 1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_17
timestamp 0
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 0
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_44
timestamp 0
transform 1 0 5152 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_52
timestamp 0
transform 1 0 5888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 0
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_98
timestamp 0
transform 1 0 10120 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_106
timestamp 0
transform 1 0 10856 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 0
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_185
timestamp 0
transform 1 0 18124 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_25
timestamp 0
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 0
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 0
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_80
timestamp 0
transform 1 0 8464 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_89
timestamp 0
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 0
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_136
timestamp 0
transform 1 0 13616 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_141
timestamp 0
transform 1 0 14076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 0
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_180
timestamp 0
transform 1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_7
timestamp 0
transform 1 0 1748 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_13
timestamp 0
transform 1 0 2300 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 0
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_38
timestamp 0
transform 1 0 4600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_50
timestamp 0
transform 1 0 5704 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_62
timestamp 0
transform 1 0 6808 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_74
timestamp 0
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_90
timestamp 0
transform 1 0 9384 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_128
timestamp 0
transform 1 0 12880 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_132
timestamp 0
transform 1 0 13248 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_149
timestamp 0
transform 1 0 14812 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_161
timestamp 0
transform 1 0 15916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_165
timestamp 0
transform 1 0 16284 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_13
timestamp 0
transform 1 0 2300 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_26
timestamp 0
transform 1 0 3496 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_33
timestamp 0
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_44
timestamp 0
transform 1 0 5152 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_70
timestamp 0
transform 1 0 7544 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_78
timestamp 0
transform 1 0 8280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_87
timestamp 0
transform 1 0 9108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 0
transform 1 0 9752 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 0
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_130
timestamp 0
transform 1 0 13064 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 0
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_145
timestamp 0
transform 1 0 14444 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 0
transform 1 0 15180 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 0
transform 1 0 15548 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_44
timestamp 0
transform 1 0 5152 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_59
timestamp 0
transform 1 0 6532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_91
timestamp 0
transform 1 0 9476 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_108
timestamp 0
transform 1 0 11040 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_116
timestamp 0
transform 1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_129
timestamp 0
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 0
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 0
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_174
timestamp 0
transform 1 0 17112 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_180
timestamp 0
transform 1 0 17664 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 0
transform 1 0 18032 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_7
timestamp 0
transform 1 0 1748 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_20
timestamp 0
transform 1 0 2944 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_29
timestamp 0
transform 1 0 3772 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 0
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_67
timestamp 0
transform 1 0 7268 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_86
timestamp 0
transform 1 0 9016 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_95
timestamp 0
transform 1 0 9844 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 0
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 0
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_140
timestamp 0
transform 1 0 13984 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_177
timestamp 0
transform 1 0 17388 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_185
timestamp 0
transform 1 0 18124 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 0
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_13
timestamp 0
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 0
transform 1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_36
timestamp 0
transform 1 0 4416 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 0
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_95
timestamp 0
transform 1 0 9844 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 0
transform 1 0 10488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_110
timestamp 0
transform 1 0 11224 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_127
timestamp 0
transform 1 0 12788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_135
timestamp 0
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 0
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_185
timestamp 0
transform 1 0 18124 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 0
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_22
timestamp 0
transform 1 0 3128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_38
timestamp 0
transform 1 0 4600 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 0
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_71
timestamp 0
transform 1 0 7636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 0
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_126
timestamp 0
transform 1 0 12696 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 0
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_182
timestamp 0
transform 1 0 17848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_13
timestamp 0
transform 1 0 2300 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 0
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_102
timestamp 0
transform 1 0 10488 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_110
timestamp 0
transform 1 0 11224 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 0
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_179
timestamp 0
transform 1 0 17572 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_185
timestamp 0
transform 1 0 18124 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_18
timestamp 0
transform 1 0 2760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_29
timestamp 0
transform 1 0 3772 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_37
timestamp 0
transform 1 0 4508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_43
timestamp 0
transform 1 0 5060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 0
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_75
timestamp 0
transform 1 0 8004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 0
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_122
timestamp 0
transform 1 0 12328 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_134
timestamp 0
transform 1 0 13432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_185
timestamp 0
transform 1 0 18124 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 0
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_19
timestamp 0
transform 1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_34
timestamp 0
transform 1 0 4232 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_40
timestamp 0
transform 1 0 4784 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_45
timestamp 0
transform 1 0 5244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_57
timestamp 0
transform 1 0 6348 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_94
timestamp 0
transform 1 0 9752 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_103
timestamp 0
transform 1 0 10580 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_123
timestamp 0
transform 1 0 12420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_134
timestamp 0
transform 1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 0
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_185
timestamp 0
transform 1 0 18124 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_14
timestamp 0
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_30
timestamp 0
transform 1 0 3864 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_42
timestamp 0
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 0
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_87
timestamp 0
transform 1 0 9108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 0
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 0
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_163
timestamp 0
transform 1 0 16100 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_172
timestamp 0
transform 1 0 16928 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 0
transform 1 0 18032 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 0
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_57
timestamp 0
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_69
timestamp 0
transform 1 0 7452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 0
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 0
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_100
timestamp 0
transform 1 0 10304 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_113
timestamp 0
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_119
timestamp 0
transform 1 0 12052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 0
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_150
timestamp 0
transform 1 0 14904 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_162
timestamp 0
transform 1 0 16008 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_169
timestamp 0
transform 1 0 16652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 0
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_185
timestamp 0
transform 1 0 18124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 0
transform -1 0 18216 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 0
transform 1 0 17848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 0
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 0
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 0
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 0
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 0
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 0
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 17848 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 8280 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform 1 0 9936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 0
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 18492 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 18492 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 18492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 18492 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 18492 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 18492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 18492 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 18492 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 18492 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 18492 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 18492 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 18492 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 18492 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 18492 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 18492 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_68
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_69
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_70
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_71
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_72
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_73
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_74
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_75
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_78
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_79
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_87
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_92
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_93
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_96
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_97
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_102
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_103
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_105
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_106
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_108
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_109
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_111
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_112
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_113
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_114
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_115
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_116
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_117
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_118
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_119
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_120
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_121
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_122
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_123
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_124
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_125
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_126
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_127
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_128
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_129
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_130
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_131
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_132
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_133
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_134
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_135
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_136
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_137
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_138
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_139
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_140
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_141
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_142
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_143
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_144
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_145
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_146
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_147
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_148
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_151
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_152
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_153
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_155
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_156
timestamp 0
transform 1 0 6256 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_157
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_158
timestamp 0
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_159
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_160
timestamp 0
transform 1 0 16560 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire19
timestamp 0
transform -1 0 13616 0 -1 15232
box -38 -48 314 592
<< labels >>
rlabel metal1 s 9798 18496 9798 18496 4 VGND
rlabel metal1 s 9798 19040 9798 19040 4 VPWR
rlabel metal1 s 16008 14042 16008 14042 4 _000_
rlabel metal1 s 13064 15470 13064 15470 4 _001_
rlabel metal1 s 16560 10234 16560 10234 4 _002_
rlabel metal2 s 15870 12002 15870 12002 4 _003_
rlabel metal1 s 15308 16762 15308 16762 4 _004_
rlabel metal2 s 16238 17918 16238 17918 4 _005_
rlabel metal2 s 14398 17884 14398 17884 4 _006_
rlabel metal1 s 12926 18156 12926 18156 4 _007_
rlabel metal2 s 17894 14994 17894 14994 4 _008_
rlabel metal1 s 15042 14586 15042 14586 4 _009_
rlabel metal1 s 17901 11118 17901 11118 4 _010_
rlabel metal2 s 16790 12376 16790 12376 4 _011_
rlabel metal1 s 17211 16490 17211 16490 4 _012_
rlabel metal2 s 16790 17816 16790 17816 4 _013_
rlabel metal1 s 15088 18598 15088 18598 4 _014_
rlabel metal1 s 13800 17850 13800 17850 4 _015_
rlabel metal1 s 14766 12614 14766 12614 4 _016_
rlabel metal1 s 13340 11662 13340 11662 4 _017_
rlabel metal1 s 5888 4046 5888 4046 4 _018_
rlabel metal2 s 12742 8670 12742 8670 4 _019_
rlabel metal2 s 12742 12002 12742 12002 4 _020_
rlabel metal1 s 2346 14382 2346 14382 4 _021_
rlabel metal2 s 14858 9061 14858 9061 4 _022_
rlabel metal4 s 11155 13124 11155 13124 4 _023_
rlabel metal2 s 14398 4998 14398 4998 4 _024_
rlabel metal2 s 7958 11798 7958 11798 4 _025_
rlabel metal2 s 9062 12495 9062 12495 4 _026_
rlabel metal1 s 11868 12138 11868 12138 4 _027_
rlabel metal1 s 14306 13974 14306 13974 4 _028_
rlabel metal2 s 4094 17561 4094 17561 4 _029_
rlabel metal1 s 3496 17510 3496 17510 4 _030_
rlabel metal1 s 9798 9690 9798 9690 4 _031_
rlabel metal2 s 16698 14807 16698 14807 4 _032_
rlabel metal1 s 13018 11084 13018 11084 4 _033_
rlabel metal1 s 13432 11186 13432 11186 4 _034_
rlabel metal3 s 16698 15861 16698 15861 4 _035_
rlabel metal1 s 15088 10642 15088 10642 4 _036_
rlabel metal1 s 14720 10778 14720 10778 4 _037_
rlabel metal2 s 2346 8993 2346 8993 4 _038_
rlabel metal1 s 12972 11322 12972 11322 4 _039_
rlabel metal1 s 13754 12206 13754 12206 4 _040_
rlabel metal1 s 5152 8942 5152 8942 4 _041_
rlabel metal1 s 8648 4590 8648 4590 4 _042_
rlabel metal1 s 8602 10540 8602 10540 4 _043_
rlabel metal1 s 16928 6766 16928 6766 4 _044_
rlabel metal1 s 6026 9588 6026 9588 4 _045_
rlabel metal1 s 7038 15368 7038 15368 4 _046_
rlabel metal1 s 8970 10574 8970 10574 4 _047_
rlabel metal2 s 8418 10234 8418 10234 4 _048_
rlabel metal1 s 5704 9146 5704 9146 4 _049_
rlabel metal1 s 4554 8330 4554 8330 4 _050_
rlabel metal1 s 4186 13226 4186 13226 4 _051_
rlabel metal1 s 8004 16150 8004 16150 4 _052_
rlabel metal1 s 6187 10030 6187 10030 4 _053_
rlabel metal2 s 6486 7548 6486 7548 4 _054_
rlabel metal1 s 11316 6842 11316 6842 4 _055_
rlabel metal1 s 16790 8500 16790 8500 4 _056_
rlabel metal2 s 11914 9010 11914 9010 4 _057_
rlabel metal1 s 6072 9690 6072 9690 4 _058_
rlabel metal1 s 8142 10064 8142 10064 4 _059_
rlabel metal2 s 8533 6358 8533 6358 4 _060_
rlabel metal1 s 10212 9554 10212 9554 4 _061_
rlabel metal2 s 8142 8874 8142 8874 4 _062_
rlabel metal1 s 9890 9588 9890 9588 4 _063_
rlabel metal1 s 9614 6970 9614 6970 4 _064_
rlabel metal2 s 15226 5406 15226 5406 4 _065_
rlabel metal1 s 10120 5338 10120 5338 4 _066_
rlabel metal1 s 10120 6970 10120 6970 4 _067_
rlabel metal1 s 9652 6630 9652 6630 4 _068_
rlabel metal1 s 9430 5780 9430 5780 4 _069_
rlabel metal1 s 7544 4794 7544 4794 4 _070_
rlabel metal2 s 8970 5032 8970 5032 4 _071_
rlabel metal2 s 7866 5474 7866 5474 4 _072_
rlabel metal2 s 8970 6052 8970 6052 4 _073_
rlabel metal1 s 8050 8058 8050 8058 4 _074_
rlabel metal2 s 9062 8653 9062 8653 4 _075_
rlabel metal1 s 11316 8942 11316 8942 4 _076_
rlabel metal2 s 8602 7106 8602 7106 4 _077_
rlabel metal1 s 5888 6290 5888 6290 4 _078_
rlabel metal1 s 7038 6970 7038 6970 4 _079_
rlabel metal1 s 8096 5814 8096 5814 4 _080_
rlabel metal1 s 9062 5168 9062 5168 4 _081_
rlabel metal1 s 9384 5338 9384 5338 4 _082_
rlabel metal1 s 8970 5746 8970 5746 4 _083_
rlabel metal1 s 8740 5882 8740 5882 4 _084_
rlabel metal1 s 15042 6664 15042 6664 4 _085_
rlabel metal2 s 14030 14892 14030 14892 4 _086_
rlabel metal3 s 14651 13804 14651 13804 4 _087_
rlabel metal2 s 5198 7786 5198 7786 4 _088_
rlabel metal1 s 10212 8058 10212 8058 4 _089_
rlabel metal1 s 14214 5338 14214 5338 4 _090_
rlabel metal1 s 16284 6222 16284 6222 4 _091_
rlabel metal1 s 15410 6426 15410 6426 4 _092_
rlabel metal2 s 14582 6188 14582 6188 4 _093_
rlabel metal2 s 14122 5967 14122 5967 4 _094_
rlabel metal1 s 11592 9078 11592 9078 4 _095_
rlabel metal1 s 11822 8330 11822 8330 4 _096_
rlabel metal2 s 12926 8194 12926 8194 4 _097_
rlabel metal2 s 17342 7378 17342 7378 4 _098_
rlabel metal1 s 5474 7922 5474 7922 4 _099_
rlabel metal1 s 16974 8568 16974 8568 4 _100_
rlabel metal2 s 17618 6460 17618 6460 4 _101_
rlabel metal2 s 17158 8551 17158 8551 4 _102_
rlabel metal1 s 16238 7922 16238 7922 4 _103_
rlabel metal1 s 15364 5066 15364 5066 4 _104_
rlabel metal1 s 14398 7412 14398 7412 4 _105_
rlabel metal1 s 14996 3978 14996 3978 4 _106_
rlabel metal2 s 15318 5508 15318 5508 4 _107_
rlabel metal1 s 14858 5338 14858 5338 4 _108_
rlabel metal2 s 11523 8058 11523 8058 4 _109_
rlabel metal1 s 9164 7922 9164 7922 4 _110_
rlabel metal1 s 11822 7888 11822 7888 4 _111_
rlabel metal1 s 14628 7242 14628 7242 4 _112_
rlabel metal1 s 14950 7514 14950 7514 4 _113_
rlabel metal1 s 14858 11186 14858 11186 4 _114_
rlabel metal1 s 4048 14450 4048 14450 4 _115_
rlabel metal1 s 7344 12138 7344 12138 4 _116_
rlabel metal1 s 7935 11526 7935 11526 4 _117_
rlabel metal2 s 14122 10710 14122 10710 4 _118_
rlabel metal1 s 12190 14042 12190 14042 4 _119_
rlabel metal1 s 12328 13294 12328 13294 4 _120_
rlabel metal1 s 11796 10608 11796 10608 4 _121_
rlabel metal2 s 6302 11237 6302 11237 4 _122_
rlabel metal2 s 12098 10438 12098 10438 4 _123_
rlabel metal1 s 13110 10642 13110 10642 4 _124_
rlabel metal2 s 15042 9180 15042 9180 4 _125_
rlabel metal3 s 13570 7803 13570 7803 4 _126_
rlabel metal1 s 14950 8466 14950 8466 4 _127_
rlabel metal2 s 13754 7140 13754 7140 4 _128_
rlabel metal1 s 14490 7888 14490 7888 4 _129_
rlabel metal1 s 13294 7412 13294 7412 4 _130_
rlabel metal2 s 13662 7650 13662 7650 4 _131_
rlabel metal1 s 7820 9554 7820 9554 4 _132_
rlabel metal1 s 10350 8976 10350 8976 4 _133_
rlabel metal1 s 7958 17136 7958 17136 4 _134_
rlabel metal1 s 12834 8024 12834 8024 4 _135_
rlabel metal1 s 15134 7956 15134 7956 4 _136_
rlabel metal1 s 13570 15028 13570 15028 4 _137_
rlabel metal1 s 12558 14518 12558 14518 4 _138_
rlabel metal2 s 12098 15300 12098 15300 4 _139_
rlabel metal2 s 11776 15470 11776 15470 4 _140_
rlabel metal1 s 10442 16014 10442 16014 4 _141_
rlabel metal2 s 12190 15776 12190 15776 4 _142_
rlabel metal1 s 11487 15878 11487 15878 4 _143_
rlabel metal1 s 10350 14348 10350 14348 4 _144_
rlabel metal1 s 11040 16014 11040 16014 4 _145_
rlabel metal1 s 10166 15674 10166 15674 4 _146_
rlabel metal2 s 5198 12376 5198 12376 4 _147_
rlabel metal1 s 7498 12954 7498 12954 4 _148_
rlabel metal1 s 10672 15674 10672 15674 4 _149_
rlabel metal2 s 11362 16864 11362 16864 4 _150_
rlabel metal3 s 12098 17187 12098 17187 4 _151_
rlabel metal2 s 12834 16932 12834 16932 4 _152_
rlabel metal2 s 12282 17408 12282 17408 4 _153_
rlabel metal2 s 10810 16966 10810 16966 4 _154_
rlabel metal1 s 11868 17646 11868 17646 4 _155_
rlabel metal1 s 12006 17748 12006 17748 4 _156_
rlabel metal1 s 9844 14994 9844 14994 4 _157_
rlabel metal2 s 9338 16966 9338 16966 4 _158_
rlabel metal1 s 9522 17306 9522 17306 4 _159_
rlabel metal2 s 7406 16966 7406 16966 4 _160_
rlabel metal1 s 8188 17238 8188 17238 4 _161_
rlabel metal1 s 10672 17578 10672 17578 4 _162_
rlabel metal2 s 11730 16218 11730 16218 4 _163_
rlabel metal2 s 9893 16422 9893 16422 4 _164_
rlabel metal1 s 3404 14586 3404 14586 4 _165_
rlabel metal2 s 9568 15538 9568 15538 4 _166_
rlabel metal2 s 9706 15300 9706 15300 4 _167_
rlabel metal1 s 9660 15674 9660 15674 4 _168_
rlabel metal1 s 12052 16082 12052 16082 4 _169_
rlabel metal2 s 11546 16932 11546 16932 4 _170_
rlabel metal1 s 5336 13838 5336 13838 4 _171_
rlabel metal1 s 6614 12240 6614 12240 4 _172_
rlabel metal1 s 6072 12206 6072 12206 4 _173_
rlabel metal1 s 6302 11594 6302 11594 4 _174_
rlabel metal1 s 2806 8908 2806 8908 4 _175_
rlabel metal2 s 7222 14620 7222 14620 4 _176_
rlabel metal2 s 3174 10387 3174 10387 4 _177_
rlabel metal1 s 3542 9452 3542 9452 4 _178_
rlabel metal1 s 3542 9622 3542 9622 4 _179_
rlabel metal2 s 2898 9146 2898 9146 4 _180_
rlabel metal2 s 2346 7548 2346 7548 4 _181_
rlabel metal3 s 5106 7395 5106 7395 4 _182_
rlabel metal2 s 3910 6630 3910 6630 4 _183_
rlabel metal1 s 6440 4454 6440 4454 4 _184_
rlabel metal1 s 5842 4794 5842 4794 4 _185_
rlabel metal1 s 2438 6324 2438 6324 4 _186_
rlabel metal1 s 3496 6358 3496 6358 4 _187_
rlabel metal1 s 3174 5882 3174 5882 4 _188_
rlabel metal1 s 1978 6222 1978 6222 4 _189_
rlabel metal2 s 1702 5882 1702 5882 4 _190_
rlabel metal1 s 2898 5712 2898 5712 4 _191_
rlabel metal1 s 2484 5882 2484 5882 4 _192_
rlabel metal2 s 1978 5882 1978 5882 4 _193_
rlabel metal1 s 8050 17510 8050 17510 4 _194_
rlabel metal1 s 8878 9146 8878 9146 4 _195_
rlabel metal1 s 8234 17680 8234 17680 4 _196_
rlabel metal3 s 15042 10693 15042 10693 4 _197_
rlabel metal2 s 11638 14280 11638 14280 4 _198_
rlabel metal1 s 2806 14416 2806 14416 4 _199_
rlabel metal1 s 8418 14484 8418 14484 4 _200_
rlabel metal1 s 8418 17646 8418 17646 4 _201_
rlabel metal1 s 9292 13498 9292 13498 4 _202_
rlabel metal2 s 8602 13124 8602 13124 4 _203_
rlabel metal2 s 8786 13702 8786 13702 4 _204_
rlabel metal1 s 8050 17646 8050 17646 4 _205_
rlabel metal1 s 10166 16592 10166 16592 4 _206_
rlabel metal3 s 8602 9979 8602 9979 4 _207_
rlabel metal3 s 9085 16660 9085 16660 4 _208_
rlabel metal2 s 8326 17748 8326 17748 4 _209_
rlabel metal1 s 7820 18122 7820 18122 4 _210_
rlabel metal1 s 7774 17850 7774 17850 4 _211_
rlabel metal2 s 9154 17119 9154 17119 4 _212_
rlabel metal2 s 7130 18054 7130 18054 4 _213_
rlabel metal1 s 7314 18190 7314 18190 4 _214_
rlabel metal2 s 4508 11118 4508 11118 4 _215_
rlabel metal1 s 4554 11322 4554 11322 4 _216_
rlabel metal1 s 5290 9146 5290 9146 4 _217_
rlabel metal1 s 4784 10778 4784 10778 4 _218_
rlabel metal1 s 4830 12172 4830 12172 4 _219_
rlabel metal1 s 4738 12138 4738 12138 4 _220_
rlabel metal1 s 4370 11730 4370 11730 4 _221_
rlabel metal1 s 13018 6324 13018 6324 4 _222_
rlabel metal3 s 4186 11747 4186 11747 4 _223_
rlabel metal2 s 2438 11458 2438 11458 4 _224_
rlabel metal1 s 13938 13498 13938 13498 4 _225_
rlabel metal2 s 13938 13056 13938 13056 4 _226_
rlabel metal1 s 14122 12818 14122 12818 4 _227_
rlabel metal1 s 3174 12648 3174 12648 4 _228_
rlabel metal1 s 2990 12206 2990 12206 4 _229_
rlabel metal2 s 2346 10370 2346 10370 4 _230_
rlabel metal1 s 2070 11220 2070 11220 4 _231_
rlabel metal1 s 1932 11322 1932 11322 4 _232_
rlabel metal2 s 2714 11934 2714 11934 4 _233_
rlabel metal1 s 2162 11866 2162 11866 4 _234_
rlabel metal2 s 12926 6494 12926 6494 4 _235_
rlabel metal2 s 10994 7072 10994 7072 4 _236_
rlabel metal1 s 6210 7820 6210 7820 4 _237_
rlabel metal2 s 10718 7106 10718 7106 4 _238_
rlabel metal1 s 10120 8942 10120 8942 4 _239_
rlabel metal1 s 8269 7446 8269 7446 4 _240_
rlabel metal1 s 7314 4726 7314 4726 4 _241_
rlabel metal1 s 6118 5338 6118 5338 4 _242_
rlabel metal1 s 5796 5746 5796 5746 4 _243_
rlabel metal2 s 6762 14382 6762 14382 4 _244_
rlabel metal1 s 6670 13498 6670 13498 4 _245_
rlabel metal3 s 6279 13804 6279 13804 4 _246_
rlabel metal1 s 2162 7956 2162 7956 4 _247_
rlabel metal1 s 1932 14382 1932 14382 4 _248_
rlabel metal1 s 1794 9146 1794 9146 4 _249_
rlabel metal1 s 10948 14042 10948 14042 4 _250_
rlabel metal1 s 10304 18258 10304 18258 4 _251_
rlabel metal2 s 7820 9894 7820 9894 4 _252_
rlabel metal1 s 8142 14790 8142 14790 4 _253_
rlabel metal1 s 7728 15130 7728 15130 4 _254_
rlabel metal1 s 7820 14042 7820 14042 4 _255_
rlabel metal1 s 7590 14586 7590 14586 4 _256_
rlabel metal2 s 10350 18496 10350 18496 4 _257_
rlabel metal1 s 9706 18088 9706 18088 4 _258_
rlabel metal1 s 11684 11866 11684 11866 4 _259_
rlabel metal1 s 10580 17646 10580 17646 4 _260_
rlabel metal2 s 10442 17204 10442 17204 4 _261_
rlabel metal1 s 9936 17850 9936 17850 4 _262_
rlabel metal3 s 11201 16660 11201 16660 4 _263_
rlabel metal1 s 10534 17850 10534 17850 4 _264_
rlabel metal1 s 9982 18258 9982 18258 4 _265_
rlabel metal2 s 4002 10234 4002 10234 4 _266_
rlabel metal1 s 4278 10064 4278 10064 4 _267_
rlabel metal2 s 3082 8636 3082 8636 4 _268_
rlabel metal1 s 4370 7344 4370 7344 4 _269_
rlabel metal1 s 4002 8262 4002 8262 4 _270_
rlabel metal1 s 2990 7412 2990 7412 4 _271_
rlabel metal2 s 2530 6970 2530 6970 4 _272_
rlabel metal2 s 3174 7106 3174 7106 4 _273_
rlabel metal1 s 5060 6766 5060 6766 4 _274_
rlabel metal1 s 5060 6834 5060 6834 4 _275_
rlabel metal1 s 3910 6970 3910 6970 4 _276_
rlabel metal1 s 2162 7276 2162 7276 4 _277_
rlabel metal1 s 15410 9010 15410 9010 4 _278_
rlabel metal1 s 15640 8602 15640 8602 4 _279_
rlabel metal1 s 14398 8602 14398 8602 4 _280_
rlabel metal1 s 11270 9112 11270 9112 4 _281_
rlabel metal1 s 13386 8908 13386 8908 4 _282_
rlabel metal1 s 10718 11662 10718 11662 4 _283_
rlabel metal1 s 13754 9520 13754 9520 4 _284_
rlabel metal2 s 13662 9180 13662 9180 4 _285_
rlabel metal1 s 13156 5678 13156 5678 4 _286_
rlabel metal1 s 17710 6324 17710 6324 4 _287_
rlabel metal2 s 13662 5848 13662 5848 4 _288_
rlabel metal1 s 12374 5168 12374 5168 4 _289_
rlabel metal2 s 12466 5406 12466 5406 4 _290_
rlabel metal1 s 12834 5712 12834 5712 4 _291_
rlabel metal2 s 12834 5355 12834 5355 4 _292_
rlabel metal2 s 13294 6086 13294 6086 4 _293_
rlabel metal1 s 12466 5644 12466 5644 4 _294_
rlabel metal1 s 11362 4794 11362 4794 4 _295_
rlabel metal2 s 10350 4794 10350 4794 4 _296_
rlabel metal1 s 10856 4590 10856 4590 4 _297_
rlabel metal2 s 10258 4352 10258 4352 4 _298_
rlabel metal1 s 9660 3910 9660 3910 4 _299_
rlabel metal2 s 9706 4522 9706 4522 4 _300_
rlabel metal1 s 9890 4114 9890 4114 4 _301_
rlabel metal3 s 10534 3893 10534 3893 4 _302_
rlabel metal2 s 17066 10438 17066 10438 4 _303_
rlabel metal1 s 17158 10574 17158 10574 4 _304_
rlabel metal1 s 16652 10778 16652 10778 4 _305_
rlabel metal1 s 9752 11866 9752 11866 4 _306_
rlabel metal2 s 10258 11594 10258 11594 4 _307_
rlabel metal3 s 4462 9996 4462 9996 4 _308_
rlabel metal1 s 3036 13294 3036 13294 4 _309_
rlabel metal2 s 2438 13736 2438 13736 4 _310_
rlabel metal1 s 2691 13702 2691 13702 4 _311_
rlabel metal1 s 3588 12410 3588 12410 4 _312_
rlabel metal1 s 3036 12682 3036 12682 4 _313_
rlabel metal1 s 2990 14042 2990 14042 4 _314_
rlabel metal1 s 4232 14382 4232 14382 4 _315_
rlabel metal1 s 3266 14348 3266 14348 4 _316_
rlabel metal1 s 2392 13838 2392 13838 4 _317_
rlabel metal2 s 1978 14280 1978 14280 4 _318_
rlabel metal1 s 2714 16150 2714 16150 4 _319_
rlabel metal2 s 5124 16558 5124 16558 4 _320_
rlabel metal1 s 2990 16524 2990 16524 4 _321_
rlabel metal1 s 3726 15674 3726 15674 4 _322_
rlabel metal1 s 3174 16592 3174 16592 4 _323_
rlabel metal2 s 2162 16218 2162 16218 4 _324_
rlabel metal2 s 1886 16762 1886 16762 4 _325_
rlabel metal1 s 3036 16082 3036 16082 4 _326_
rlabel metal2 s 2530 16422 2530 16422 4 _327_
rlabel metal1 s 15778 12920 15778 12920 4 _328_
rlabel metal1 s 13386 17680 13386 17680 4 _329_
rlabel metal1 s 14858 16694 14858 16694 4 _330_
rlabel metal2 s 13018 18054 13018 18054 4 _331_
rlabel metal2 s 13202 18054 13202 18054 4 _332_
rlabel metal1 s 16008 18258 16008 18258 4 _333_
rlabel metal2 s 17710 10523 17710 10523 4 _334_
rlabel metal2 s 16330 4930 16330 4930 4 _335_
rlabel metal1 s 6854 8330 6854 8330 4 _336_
rlabel metal2 s 2254 14433 2254 14433 4 _337_
rlabel metal1 s 15640 4794 15640 4794 4 _338_
rlabel metal2 s 5198 14943 5198 14943 4 _339_
rlabel metal1 s 8510 12818 8510 12818 4 _340_
rlabel metal1 s 12972 9350 12972 9350 4 _341_
rlabel metal2 s 15226 4318 15226 4318 4 _342_
rlabel metal2 s 8326 11900 8326 11900 4 _343_
rlabel metal1 s 8740 5202 8740 5202 4 _344_
rlabel metal1 s 7130 4624 7130 4624 4 _345_
rlabel metal2 s 3358 6052 3358 6052 4 _346_
rlabel metal1 s 15870 11730 15870 11730 4 _347_
rlabel metal2 s 7038 16830 7038 16830 4 _348_
rlabel metal1 s 8878 12886 8878 12886 4 _349_
rlabel metal1 s 8372 4182 8372 4182 4 _350_
rlabel metal2 s 15226 8024 15226 8024 4 _351_
rlabel metal1 s 14168 17170 14168 17170 4 _352_
rlabel metal1 s 15870 6732 15870 6732 4 _353_
rlabel metal1 s 16192 9962 16192 9962 4 _354_
rlabel metal1 s 15226 11118 15226 11118 4 _355_
rlabel metal1 s 2668 9554 2668 9554 4 _356_
rlabel metal1 s 11684 10234 11684 10234 4 _357_
rlabel metal1 s 14904 12886 14904 12886 4 _358_
rlabel metal1 s 6762 8942 6762 8942 4 _359_
rlabel metal2 s 11270 4420 11270 4420 4 _360_
rlabel metal1 s 6762 7888 6762 7888 4 _361_
rlabel metal2 s 12282 6732 12282 6732 4 _362_
rlabel metal2 s 14950 12138 14950 12138 4 _363_
rlabel metal1 s 15410 12410 15410 12410 4 _364_
rlabel metal1 s 5520 10778 5520 10778 4 _365_
rlabel metal1 s 4094 11322 4094 11322 4 _366_
rlabel metal1 s 16698 5678 16698 5678 4 _367_
rlabel metal2 s 6854 15810 6854 15810 4 _368_
rlabel metal1 s 13202 16218 13202 16218 4 _369_
rlabel metal1 s 8418 15028 8418 15028 4 _370_
rlabel metal1 s 13386 12852 13386 12852 4 _371_
rlabel metal2 s 14398 7650 14398 7650 4 _372_
rlabel metal2 s 3450 16456 3450 16456 4 _373_
rlabel metal1 s 12466 13192 12466 13192 4 _374_
rlabel metal2 s 7498 6460 7498 6460 4 _375_
rlabel metal1 s 5474 13226 5474 13226 4 _376_
rlabel metal1 s 14076 12886 14076 12886 4 _377_
rlabel metal1 s 13616 4250 13616 4250 4 _378_
rlabel metal1 s 13570 6324 13570 6324 4 _379_
rlabel metal2 s 7038 15470 7038 15470 4 _380_
rlabel metal1 s 15134 10778 15134 10778 4 _381_
rlabel metal1 s 7820 4794 7820 4794 4 _382_
rlabel metal2 s 14490 13498 14490 13498 4 _383_
rlabel metal1 s 9154 7820 9154 7820 4 _384_
rlabel metal2 s 13110 12597 13110 12597 4 _385_
rlabel metal1 s 14444 12682 14444 12682 4 _386_
rlabel metal1 s 17526 14314 17526 14314 4 clk
rlabel metal1 s 16146 14586 16146 14586 4 clknet_0_clk
rlabel metal1 s 16790 13158 16790 13158 4 clknet_1_0__leaf_clk
rlabel metal2 s 14122 16558 14122 16558 4 clknet_1_1__leaf_clk
rlabel metal2 s 13938 18190 13938 18190 4 net1
rlabel metal1 s 16790 7854 16790 7854 4 net10
rlabel metal1 s 11546 17850 11546 17850 4 net11
rlabel metal2 s 2070 7174 2070 7174 4 net12
rlabel metal2 s 8050 18564 8050 18564 4 net13
rlabel metal2 s 1702 11322 1702 11322 4 net14
rlabel metal1 s 1610 8058 1610 8058 4 net15
rlabel metal2 s 9430 18564 9430 18564 4 net16
rlabel metal2 s 1702 6970 1702 6970 4 net17
rlabel metal1 s 5290 8976 5290 8976 4 net18
rlabel metal2 s 12650 14586 12650 14586 4 net19
rlabel metal1 s 16698 12750 16698 12750 4 net2
rlabel metal1 s 2300 14450 2300 14450 4 net20
rlabel metal1 s 10166 15096 10166 15096 4 net21
rlabel metal1 s 9246 6120 9246 6120 4 net22
rlabel metal2 s 9154 4930 9154 4930 4 net23
rlabel metal1 s 5842 10642 5842 10642 4 net24
rlabel metal1 s 2208 9554 2208 9554 4 net25
rlabel metal1 s 8004 4998 8004 4998 4 net26
rlabel metal1 s 11638 8466 11638 8466 4 net27
rlabel metal1 s 14674 5882 14674 5882 4 net28
rlabel metal1 s 8878 4148 8878 4148 4 net29
rlabel metal2 s 12052 5202 12052 5202 4 net3
rlabel metal1 s 8786 13974 8786 13974 4 net30
rlabel metal2 s 6210 16762 6210 16762 4 net31
rlabel metal1 s 14490 14994 14490 14994 4 net32
rlabel metal1 s 7728 15470 7728 15470 4 net33
rlabel metal1 s 15318 7854 15318 7854 4 net34
rlabel metal1 s 1978 8908 1978 8908 4 net35
rlabel metal1 s 12604 5678 12604 5678 4 net36
rlabel metal1 s 3726 8942 3726 8942 4 net37
rlabel metal1 s 3542 17136 3542 17136 4 net38
rlabel metal1 s 13846 12818 13846 12818 4 net39
rlabel metal1 s 1610 9690 1610 9690 4 net4
rlabel metal1 s 8970 18156 8970 18156 4 net40
rlabel metal1 s 2714 8976 2714 8976 4 net41
rlabel metal1 s 2691 13294 2691 13294 4 net42
rlabel metal1 s 9384 13906 9384 13906 4 net43
rlabel metal2 s 5566 7769 5566 7769 4 net44
rlabel metal2 s 5106 13532 5106 13532 4 net45
rlabel metal1 s 6946 11764 6946 11764 4 net46
rlabel metal1 s 8142 9554 8142 9554 4 net47
rlabel metal1 s 10028 5202 10028 5202 4 net48
rlabel metal2 s 14214 12988 14214 12988 4 net49
rlabel metal2 s 1702 13498 1702 13498 4 net5
rlabel metal1 s 16606 8908 16606 8908 4 net50
rlabel metal1 s 3772 4590 3772 4590 4 net51
rlabel metal1 s 7268 12614 7268 12614 4 net52
rlabel metal2 s 6210 15810 6210 15810 4 net53
rlabel metal1 s 9890 13362 9890 13362 4 net54
rlabel metal1 s 9476 7854 9476 7854 4 net55
rlabel metal2 s 15962 7038 15962 7038 4 net56
rlabel metal2 s 11868 5134 11868 5134 4 net57
rlabel metal1 s 12328 15470 12328 15470 4 net58
rlabel metal2 s 16957 14994 16957 14994 4 net59
rlabel metal2 s 1702 15674 1702 15674 4 net6
rlabel metal1 s 13570 13328 13570 13328 4 net60
rlabel metal1 s 4094 9044 4094 9044 4 net61
rlabel metal1 s 8694 4012 8694 4012 4 net62
rlabel metal2 s 6302 16354 6302 16354 4 net63
rlabel metal1 s 7038 16116 7038 16116 4 net64
rlabel metal1 s 12374 4114 12374 4114 4 net65
rlabel metal2 s 15778 5100 15778 5100 4 net66
rlabel metal1 s 15410 10064 15410 10064 4 net67
rlabel metal1 s 15916 14314 15916 14314 4 net68
rlabel metal1 s 17296 9622 17296 9622 4 net69
rlabel metal1 s 1610 16762 1610 16762 4 net7
rlabel metal1 s 7061 7854 7061 7854 4 net70
rlabel metal1 s 4232 12818 4232 12818 4 net71
rlabel metal2 s 7866 16031 7866 16031 4 net72
rlabel metal1 s 13478 4012 13478 4012 4 net73
rlabel metal1 s 14306 14960 14306 14960 4 net74
rlabel metal2 s 4140 6766 4140 6766 4 net75
rlabel metal1 s 9108 4114 9108 4114 4 net76
rlabel metal2 s 16790 13430 16790 13430 4 net77
rlabel metal1 s 12834 3978 12834 3978 4 net78
rlabel metal3 s 15042 14331 15042 14331 4 net79
rlabel metal2 s 1610 14790 1610 14790 4 net8
rlabel metal1 s 9108 2414 9108 2414 4 net9
rlabel metal2 s 18078 14161 18078 14161 4 rst
rlabel metal3 s 18454 12308 18454 12308 4 sine_out[0]
rlabel metal2 s 11638 1520 11638 1520 4 sine_out[10]
rlabel metal3 s 1096 9588 1096 9588 4 sine_out[11]
rlabel metal1 s 1426 13498 1426 13498 4 sine_out[12]
rlabel metal1 s 1426 15674 1426 15674 4 sine_out[13]
rlabel metal3 s 1096 16388 1096 16388 4 sine_out[14]
rlabel metal3 s 0 14288 800 14408 4 sine_out[15]
port 11 nsew
rlabel metal2 s 9062 1520 9062 1520 4 sine_out[1]
rlabel metal2 s 18078 7633 18078 7633 4 sine_out[2]
rlabel metal1 s 11776 18938 11776 18938 4 sine_out[3]
rlabel metal3 s 1280 7548 1280 7548 4 sine_out[4]
rlabel metal1 s 8142 18938 8142 18938 4 sine_out[5]
rlabel metal1 s 1334 11322 1334 11322 4 sine_out[6]
rlabel metal3 s 1096 8228 1096 8228 4 sine_out[7]
rlabel metal1 s 9936 18938 9936 18938 4 sine_out[8]
rlabel metal3 s 0 6808 800 6928 4 sine_out[9]
port 20 nsew
rlabel metal1 s 17618 12886 17618 12886 4 tcout\[0\]
rlabel metal2 s 13110 15147 13110 15147 4 tcout\[1\]
rlabel metal1 s 18032 9622 18032 9622 4 tcout\[2\]
rlabel metal2 s 17802 11900 17802 11900 4 tcout\[3\]
rlabel metal2 s 16698 17918 16698 17918 4 tcout\[4\]
rlabel metal2 s 17710 17119 17710 17119 4 tcout\[5\]
rlabel metal2 s 15962 16796 15962 16796 4 tcout\[6\]
rlabel metal1 s 12857 18394 12857 18394 4 tcout\[7\]
flabel metal4 s 4868 2128 5188 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4208 2128 4528 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 18812 13608 19612 13728 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 18812 14288 19612 14408 0 FreeSans 600 0 0 0 rst
port 4 nsew
flabel metal3 s 18812 12248 19612 12368 0 FreeSans 600 0 0 0 sine_out[0]
port 5 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 sine_out[10]
port 6 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 sine_out[11]
port 7 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 sine_out[12]
port 8 nsew
flabel metal3 s 0 15648 800 15768 0 FreeSans 600 0 0 0 sine_out[13]
port 9 nsew
flabel metal3 s 0 16328 800 16448 0 FreeSans 600 0 0 0 sine_out[14]
port 10 nsew
flabel metal3 s 400 14348 400 14348 0 FreeSans 600 0 0 0 sine_out[15]
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 sine_out[1]
port 12 nsew
flabel metal3 s 18812 7488 19612 7608 0 FreeSans 600 0 0 0 sine_out[2]
port 13 nsew
flabel metal2 s 11610 20956 11666 21756 0 FreeSans 280 90 0 0 sine_out[3]
port 14 nsew
flabel metal3 s 0 7488 800 7608 0 FreeSans 600 0 0 0 sine_out[4]
port 15 nsew
flabel metal2 s 7746 20956 7802 21756 0 FreeSans 280 90 0 0 sine_out[5]
port 16 nsew
flabel metal3 s 0 11568 800 11688 0 FreeSans 600 0 0 0 sine_out[6]
port 17 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 sine_out[7]
port 18 nsew
flabel metal2 s 9678 20956 9734 21756 0 FreeSans 280 90 0 0 sine_out[8]
port 19 nsew
flabel metal3 s 400 6868 400 6868 0 FreeSans 600 0 0 0 sine_out[9]
<< properties >>
string FIXED_BBOX 0 0 19612 21756
<< end >>
