module counter (clk,
    csb00,
    csb01,
    rst,
    addr00,
    addr01,
    denum,
    din00,
    din01,
    num,
    sine_out);
 input clk;
 input csb00;
 input csb01;
 input rst;
 input [7:0] addr00;
 input [7:0] addr01;
 input [3:0] denum;
 input [15:0] din00;
 input [15:0] din01;
 input [3:0] num;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire net115;
 wire clknet_0_clk;
 wire \sine_out_reg0[0] ;
 wire \sine_out_reg0[10] ;
 wire \sine_out_reg0[11] ;
 wire \sine_out_reg0[12] ;
 wire \sine_out_reg0[13] ;
 wire \sine_out_reg0[14] ;
 wire \sine_out_reg0[15] ;
 wire \sine_out_reg0[1] ;
 wire \sine_out_reg0[2] ;
 wire \sine_out_reg0[3] ;
 wire \sine_out_reg0[4] ;
 wire \sine_out_reg0[5] ;
 wire \sine_out_reg0[6] ;
 wire \sine_out_reg0[7] ;
 wire \sine_out_reg0[8] ;
 wire \sine_out_reg0[9] ;
 wire \sine_out_reg1[0] ;
 wire \sine_out_reg1[10] ;
 wire \sine_out_reg1[11] ;
 wire \sine_out_reg1[12] ;
 wire \sine_out_reg1[13] ;
 wire \sine_out_reg1[14] ;
 wire \sine_out_reg1[15] ;
 wire \sine_out_reg1[1] ;
 wire \sine_out_reg1[2] ;
 wire \sine_out_reg1[3] ;
 wire \sine_out_reg1[4] ;
 wire \sine_out_reg1[5] ;
 wire \sine_out_reg1[6] ;
 wire \sine_out_reg1[7] ;
 wire \sine_out_reg1[8] ;
 wire \sine_out_reg1[9] ;
 wire \sine_out_temp0[0] ;
 wire \sine_out_temp0[10] ;
 wire \sine_out_temp0[11] ;
 wire \sine_out_temp0[12] ;
 wire \sine_out_temp0[13] ;
 wire \sine_out_temp0[14] ;
 wire \sine_out_temp0[15] ;
 wire \sine_out_temp0[1] ;
 wire \sine_out_temp0[2] ;
 wire \sine_out_temp0[3] ;
 wire \sine_out_temp0[4] ;
 wire \sine_out_temp0[5] ;
 wire \sine_out_temp0[6] ;
 wire \sine_out_temp0[7] ;
 wire \sine_out_temp0[8] ;
 wire \sine_out_temp0[9] ;
 wire \sine_out_temp1[0] ;
 wire \sine_out_temp1[10] ;
 wire \sine_out_temp1[11] ;
 wire \sine_out_temp1[12] ;
 wire \sine_out_temp1[13] ;
 wire \sine_out_temp1[14] ;
 wire \sine_out_temp1[15] ;
 wire \sine_out_temp1[1] ;
 wire \sine_out_temp1[2] ;
 wire \sine_out_temp1[3] ;
 wire \sine_out_temp1[4] ;
 wire \sine_out_temp1[5] ;
 wire \sine_out_temp1[6] ;
 wire \sine_out_temp1[7] ;
 wire \sine_out_temp1[8] ;
 wire \sine_out_temp1[9] ;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;
 wire \tcout[8] ;
 wire \tcout_delay[0] ;
 wire \tcout_delay[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sky130_fd_sc_hd__inv_2 _293_ (.A(net22),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _294_ (.A(net21),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _295_ (.A(net19),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _296_ (.A(net113),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _297_ (.A(net107),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _298_ (.A(net111),
    .Y(_055_));
 sky130_fd_sc_hd__clkinv_4 _299_ (.A(net110),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _300_ (.A(net105),
    .Y(_025_));
 sky130_fd_sc_hd__or2_1 _301_ (.A(net106),
    .B(net109),
    .X(_057_));
 sky130_fd_sc_hd__or4b_1 _302_ (.A(net108),
    .B(net111),
    .C(net109),
    .D_N(net113),
    .X(_058_));
 sky130_fd_sc_hd__or3b_1 _303_ (.A(_050_),
    .B(net111),
    .C_N(_058_),
    .X(_059_));
 sky130_fd_sc_hd__nand2_1 _304_ (.A(_050_),
    .B(net111),
    .Y(_060_));
 sky130_fd_sc_hd__nand2_1 _305_ (.A(_051_),
    .B(net113),
    .Y(_061_));
 sky130_fd_sc_hd__and3_1 _306_ (.A(_059_),
    .B(_060_),
    .C(_061_),
    .X(_062_));
 sky130_fd_sc_hd__a221o_1 _307_ (.A1(_051_),
    .A2(net113),
    .B1(net111),
    .B2(_050_),
    .C1(_057_),
    .X(_063_));
 sky130_fd_sc_hd__a21boi_1 _308_ (.A1(net22),
    .A2(_058_),
    .B1_N(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__a21oi_1 _309_ (.A1(_059_),
    .A2(_060_),
    .B1(_061_),
    .Y(_065_));
 sky130_fd_sc_hd__o21ba_1 _310_ (.A1(_062_),
    .A2(_065_),
    .B1_N(_063_),
    .X(_066_));
 sky130_fd_sc_hd__nand2_1 _311_ (.A(_050_),
    .B(net108),
    .Y(_067_));
 sky130_fd_sc_hd__a2111o_1 _312_ (.A1(_050_),
    .A2(net111),
    .B1(_057_),
    .C1(_051_),
    .D1(_053_),
    .X(_068_));
 sky130_fd_sc_hd__nand2_1 _313_ (.A(net21),
    .B(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__and3_1 _314_ (.A(net21),
    .B(_055_),
    .C(_068_),
    .X(_070_));
 sky130_fd_sc_hd__a21o_1 _315_ (.A1(net21),
    .A2(_068_),
    .B1(_055_),
    .X(_071_));
 sky130_fd_sc_hd__and2b_1 _316_ (.A_N(_070_),
    .B(_071_),
    .X(_072_));
 sky130_fd_sc_hd__or2_1 _317_ (.A(net20),
    .B(_053_),
    .X(_073_));
 sky130_fd_sc_hd__a21oi_1 _318_ (.A1(_071_),
    .A2(_073_),
    .B1(_070_),
    .Y(_074_));
 sky130_fd_sc_hd__nand2_1 _319_ (.A(net109),
    .B(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__or2_1 _320_ (.A(net109),
    .B(_074_),
    .X(_076_));
 sky130_fd_sc_hd__a311o_1 _321_ (.A1(_054_),
    .A2(_075_),
    .A3(_076_),
    .B1(_064_),
    .C1(_066_),
    .X(_077_));
 sky130_fd_sc_hd__nor2_1 _322_ (.A(net108),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__o31a_1 _323_ (.A1(net109),
    .A2(_064_),
    .A3(_066_),
    .B1(_074_),
    .X(_079_));
 sky130_fd_sc_hd__a21o_1 _324_ (.A1(_050_),
    .A2(net110),
    .B1(net108),
    .X(_080_));
 sky130_fd_sc_hd__nor2_1 _325_ (.A(_079_),
    .B(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__xnor2_1 _326_ (.A(_072_),
    .B(_073_),
    .Y(_082_));
 sky130_fd_sc_hd__mux2_1 _327_ (.A0(_069_),
    .A1(_082_),
    .S(_081_),
    .X(_083_));
 sky130_fd_sc_hd__nor2_1 _328_ (.A(net110),
    .B(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__xnor2_1 _329_ (.A(_056_),
    .B(_083_),
    .Y(_085_));
 sky130_fd_sc_hd__o31ai_1 _330_ (.A1(_053_),
    .A2(_079_),
    .A3(_080_),
    .B1(net20),
    .Y(_086_));
 sky130_fd_sc_hd__or4_1 _331_ (.A(net20),
    .B(_053_),
    .C(_079_),
    .D(_080_),
    .X(_087_));
 sky130_fd_sc_hd__and2_1 _332_ (.A(net86),
    .B(_087_),
    .X(_088_));
 sky130_fd_sc_hd__a21o_1 _333_ (.A1(net85),
    .A2(_087_),
    .B1(net111),
    .X(_089_));
 sky130_fd_sc_hd__nand3_1 _334_ (.A(net112),
    .B(_086_),
    .C(_087_),
    .Y(_090_));
 sky130_fd_sc_hd__nand2_1 _335_ (.A(_052_),
    .B(net113),
    .Y(_091_));
 sky130_fd_sc_hd__and3_1 _336_ (.A(_089_),
    .B(_090_),
    .C(_091_),
    .X(_092_));
 sky130_fd_sc_hd__a21bo_1 _337_ (.A1(_090_),
    .A2(_091_),
    .B1_N(_089_),
    .X(_093_));
 sky130_fd_sc_hd__a211o_1 _338_ (.A1(_085_),
    .A2(_093_),
    .B1(_078_),
    .C1(_084_),
    .X(_094_));
 sky130_fd_sc_hd__and2_1 _339_ (.A(_067_),
    .B(_094_),
    .X(_095_));
 sky130_fd_sc_hd__inv_2 _340_ (.A(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__xnor2_1 _341_ (.A(_085_),
    .B(_093_),
    .Y(_097_));
 sky130_fd_sc_hd__mux2_1 _342_ (.A0(_083_),
    .A1(_097_),
    .S(_095_),
    .X(_098_));
 sky130_fd_sc_hd__xnor2_1 _343_ (.A(net107),
    .B(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_1 _344_ (.A1(_089_),
    .A2(_090_),
    .B1(_091_),
    .Y(_100_));
 sky130_fd_sc_hd__or2_1 _345_ (.A(_092_),
    .B(_100_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _346_ (.A0(_088_),
    .A1(_101_),
    .S(_095_),
    .X(_102_));
 sky130_fd_sc_hd__or2_1 _347_ (.A(net110),
    .B(_102_),
    .X(_103_));
 sky130_fd_sc_hd__and2_1 _348_ (.A(net110),
    .B(_102_),
    .X(_104_));
 sky130_fd_sc_hd__a31o_1 _349_ (.A1(net113),
    .A2(_067_),
    .A3(_094_),
    .B1(_052_),
    .X(_105_));
 sky130_fd_sc_hd__nand3b_1 _350_ (.A_N(_091_),
    .B(_094_),
    .C(_067_),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_1 _351_ (.A(_105_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__a21oi_1 _352_ (.A1(_105_),
    .A2(_106_),
    .B1(net112),
    .Y(_108_));
 sky130_fd_sc_hd__and3_1 _353_ (.A(net112),
    .B(_105_),
    .C(_106_),
    .X(_109_));
 sky130_fd_sc_hd__or2_1 _354_ (.A(_108_),
    .B(_109_),
    .X(_110_));
 sky130_fd_sc_hd__o21ba_1 _355_ (.A1(net113),
    .A2(_109_),
    .B1_N(_108_),
    .X(_111_));
 sky130_fd_sc_hd__a21o_1 _356_ (.A1(_103_),
    .A2(_111_),
    .B1(_104_),
    .X(_112_));
 sky130_fd_sc_hd__a211o_2 _357_ (.A1(_103_),
    .A2(_111_),
    .B1(_104_),
    .C1(_099_),
    .X(_113_));
 sky130_fd_sc_hd__or3_1 _358_ (.A(_062_),
    .B(_063_),
    .C(_065_),
    .X(_114_));
 sky130_fd_sc_hd__o221a_2 _359_ (.A1(_077_),
    .A2(_095_),
    .B1(_098_),
    .B2(net107),
    .C1(_114_),
    .X(_115_));
 sky130_fd_sc_hd__and2_1 _360_ (.A(_113_),
    .B(_115_),
    .X(_116_));
 sky130_fd_sc_hd__nand2_2 _361_ (.A(_113_),
    .B(_115_),
    .Y(_117_));
 sky130_fd_sc_hd__a21bo_1 _362_ (.A1(_098_),
    .A2(_115_),
    .B1_N(_113_),
    .X(_118_));
 sky130_fd_sc_hd__a21oi_2 _363_ (.A1(_099_),
    .A2(_112_),
    .B1(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__xnor2_1 _364_ (.A(_056_),
    .B(_102_),
    .Y(_120_));
 sky130_fd_sc_hd__nand2_1 _365_ (.A(_111_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__or2_1 _366_ (.A(_111_),
    .B(_120_),
    .X(_122_));
 sky130_fd_sc_hd__nand3b_1 _367_ (.A_N(_102_),
    .B(_113_),
    .C(_115_),
    .Y(_123_));
 sky130_fd_sc_hd__a22o_1 _368_ (.A1(_113_),
    .A2(_115_),
    .B1(_121_),
    .B2(_122_),
    .X(_124_));
 sky130_fd_sc_hd__and2_1 _369_ (.A(_123_),
    .B(_124_),
    .X(_125_));
 sky130_fd_sc_hd__a21oi_1 _370_ (.A1(_123_),
    .A2(_124_),
    .B1(net107),
    .Y(_126_));
 sky130_fd_sc_hd__nand2_1 _371_ (.A(net107),
    .B(_125_),
    .Y(_127_));
 sky130_fd_sc_hd__and3_1 _372_ (.A(_107_),
    .B(_113_),
    .C(_115_),
    .X(_128_));
 sky130_fd_sc_hd__xnor2_1 _373_ (.A(_053_),
    .B(_110_),
    .Y(_129_));
 sky130_fd_sc_hd__a21o_1 _374_ (.A1(_113_),
    .A2(_115_),
    .B1(_129_),
    .X(_130_));
 sky130_fd_sc_hd__o21a_1 _375_ (.A1(_107_),
    .A2(_117_),
    .B1(_130_),
    .X(_131_));
 sky130_fd_sc_hd__inv_2 _376_ (.A(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__o211a_1 _377_ (.A1(_107_),
    .A2(_117_),
    .B1(_130_),
    .C1(_056_),
    .X(_133_));
 sky130_fd_sc_hd__a211o_1 _378_ (.A1(_117_),
    .A2(_129_),
    .B1(_128_),
    .C1(_056_),
    .X(_134_));
 sky130_fd_sc_hd__and2b_1 _379_ (.A_N(_133_),
    .B(_134_),
    .X(_135_));
 sky130_fd_sc_hd__a21oi_2 _380_ (.A1(net113),
    .A2(_116_),
    .B1(net112),
    .Y(_136_));
 sky130_fd_sc_hd__a21oi_1 _381_ (.A1(_134_),
    .A2(_136_),
    .B1(_133_),
    .Y(_137_));
 sky130_fd_sc_hd__a211o_1 _382_ (.A1(_134_),
    .A2(_136_),
    .B1(_126_),
    .C1(_133_),
    .X(_138_));
 sky130_fd_sc_hd__a21oi_1 _383_ (.A1(_127_),
    .A2(_138_),
    .B1(_119_),
    .Y(_139_));
 sky130_fd_sc_hd__inv_2 _384_ (.A(net84),
    .Y(_140_));
 sky130_fd_sc_hd__xnor2_1 _385_ (.A(_135_),
    .B(_136_),
    .Y(_141_));
 sky130_fd_sc_hd__mux2_1 _386_ (.A0(_141_),
    .A1(_132_),
    .S(_139_),
    .X(_142_));
 sky130_fd_sc_hd__nand2_2 _387_ (.A(net107),
    .B(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__a211oi_1 _388_ (.A1(_127_),
    .A2(_138_),
    .B1(_053_),
    .C1(_119_),
    .Y(_144_));
 sky130_fd_sc_hd__and3_1 _389_ (.A(net113),
    .B(net112),
    .C(_116_),
    .X(_145_));
 sky130_fd_sc_hd__or2_1 _390_ (.A(_136_),
    .B(_145_),
    .X(_146_));
 sky130_fd_sc_hd__o2bb2a_1 _391_ (.A1_N(_117_),
    .A2_N(net81),
    .B1(_146_),
    .B2(net84),
    .X(_147_));
 sky130_fd_sc_hd__nand2_1 _392_ (.A(net110),
    .B(_147_),
    .Y(_148_));
 sky130_fd_sc_hd__nor2_1 _393_ (.A(net112),
    .B(net81),
    .Y(_149_));
 sky130_fd_sc_hd__o21bai_2 _394_ (.A1(net110),
    .A2(_147_),
    .B1_N(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__and2_1 _395_ (.A(_148_),
    .B(_150_),
    .X(_151_));
 sky130_fd_sc_hd__nand2_1 _396_ (.A(_143_),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__or2_1 _397_ (.A(net107),
    .B(_142_),
    .X(_153_));
 sky130_fd_sc_hd__xnor2_1 _398_ (.A(_054_),
    .B(_137_),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_1 _399_ (.A(_119_),
    .B(_125_),
    .Y(_155_));
 sky130_fd_sc_hd__mux2_1 _400_ (.A0(_125_),
    .A1(_155_),
    .S(_154_),
    .X(_156_));
 sky130_fd_sc_hd__o21ai_2 _401_ (.A1(net107),
    .A2(_142_),
    .B1(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__a31oi_4 _402_ (.A1(_143_),
    .A2(_148_),
    .A3(_150_),
    .B1(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(_143_),
    .B(_153_),
    .Y(_159_));
 sky130_fd_sc_hd__xor2_1 _404_ (.A(_151_),
    .B(_159_),
    .X(_160_));
 sky130_fd_sc_hd__mux2_1 _405_ (.A0(_160_),
    .A1(_142_),
    .S(_158_),
    .X(_161_));
 sky130_fd_sc_hd__a21o_1 _406_ (.A1(_152_),
    .A2(_153_),
    .B1(_156_),
    .X(_162_));
 sky130_fd_sc_hd__nand3_1 _407_ (.A(_119_),
    .B(_127_),
    .C(_138_),
    .Y(_163_));
 sky130_fd_sc_hd__nand4_1 _408_ (.A(_114_),
    .B(_161_),
    .C(_162_),
    .D(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__xnor2_1 _409_ (.A(_056_),
    .B(_147_),
    .Y(_165_));
 sky130_fd_sc_hd__xnor2_1 _410_ (.A(_149_),
    .B(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__mux2_1 _411_ (.A0(_166_),
    .A1(_147_),
    .S(_158_),
    .X(_167_));
 sky130_fd_sc_hd__nor2_1 _412_ (.A(net107),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__nand2_1 _413_ (.A(net107),
    .B(_167_),
    .Y(_169_));
 sky130_fd_sc_hd__a311oi_2 _414_ (.A1(_143_),
    .A2(_148_),
    .A3(_150_),
    .B1(_157_),
    .C1(_053_),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_1 _415_ (.A(net112),
    .B(net82),
    .Y(_171_));
 sky130_fd_sc_hd__nand2b_1 _416_ (.A_N(_149_),
    .B(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__o2bb2a_1 _417_ (.A1_N(_140_),
    .A2_N(_170_),
    .B1(_172_),
    .B2(_158_),
    .X(_173_));
 sky130_fd_sc_hd__nor2_1 _418_ (.A(net110),
    .B(_173_),
    .Y(_174_));
 sky130_fd_sc_hd__xnor2_1 _419_ (.A(_056_),
    .B(_173_),
    .Y(_175_));
 sky130_fd_sc_hd__nor2_1 _420_ (.A(net112),
    .B(_170_),
    .Y(_176_));
 sky130_fd_sc_hd__a21o_1 _421_ (.A1(net79),
    .A2(net80),
    .B1(_174_),
    .X(_177_));
 sky130_fd_sc_hd__a211o_1 _422_ (.A1(_175_),
    .A2(net80),
    .B1(_168_),
    .C1(_174_),
    .X(_178_));
 sky130_fd_sc_hd__a21o_1 _423_ (.A1(_169_),
    .A2(_178_),
    .B1(_164_),
    .X(_179_));
 sky130_fd_sc_hd__xnor2_1 _424_ (.A(net79),
    .B(net80),
    .Y(_180_));
 sky130_fd_sc_hd__mux2_1 _425_ (.A0(_173_),
    .A1(_180_),
    .S(_179_),
    .X(_181_));
 sky130_fd_sc_hd__inv_2 _426_ (.A(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__or2_1 _427_ (.A(net106),
    .B(_181_),
    .X(_183_));
 sky130_fd_sc_hd__xnor2_1 _428_ (.A(net106),
    .B(_181_),
    .Y(_184_));
 sky130_fd_sc_hd__a211o_1 _429_ (.A1(_169_),
    .A2(_178_),
    .B1(_053_),
    .C1(_164_),
    .X(_185_));
 sky130_fd_sc_hd__and2_1 _430_ (.A(net112),
    .B(_170_),
    .X(_186_));
 sky130_fd_sc_hd__nor2_1 _431_ (.A(_176_),
    .B(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__o2bb2a_1 _432_ (.A1_N(_187_),
    .A2_N(_179_),
    .B1(_158_),
    .B2(_185_),
    .X(_188_));
 sky130_fd_sc_hd__and2_1 _433_ (.A(net109),
    .B(_188_),
    .X(_189_));
 sky130_fd_sc_hd__and2_1 _434_ (.A(_055_),
    .B(_185_),
    .X(_190_));
 sky130_fd_sc_hd__o21ba_1 _435_ (.A1(net109),
    .A2(_188_),
    .B1_N(_190_),
    .X(_191_));
 sky130_fd_sc_hd__or2_1 _436_ (.A(_189_),
    .B(_191_),
    .X(_192_));
 sky130_fd_sc_hd__nand2b_1 _437_ (.A_N(_168_),
    .B(_169_),
    .Y(_193_));
 sky130_fd_sc_hd__xor2_1 _438_ (.A(_177_),
    .B(_193_),
    .X(_194_));
 sky130_fd_sc_hd__mux2_1 _439_ (.A0(_167_),
    .A1(_194_),
    .S(_179_),
    .X(_195_));
 sky130_fd_sc_hd__o311a_1 _440_ (.A1(_184_),
    .A2(_189_),
    .A3(_191_),
    .B1(_195_),
    .C1(_183_),
    .X(_196_));
 sky130_fd_sc_hd__xnor2_1 _441_ (.A(_056_),
    .B(_188_),
    .Y(_197_));
 sky130_fd_sc_hd__xnor2_1 _442_ (.A(_190_),
    .B(_197_),
    .Y(_198_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(_198_),
    .A1(_188_),
    .S(net78),
    .X(_199_));
 sky130_fd_sc_hd__and2_1 _444_ (.A(net106),
    .B(_199_),
    .X(_200_));
 sky130_fd_sc_hd__nand2_1 _445_ (.A(net106),
    .B(_199_),
    .Y(_201_));
 sky130_fd_sc_hd__nand2_1 _446_ (.A(net113),
    .B(_179_),
    .Y(_202_));
 sky130_fd_sc_hd__nor2_1 _447_ (.A(_055_),
    .B(_185_),
    .Y(_203_));
 sky130_fd_sc_hd__or2_1 _448_ (.A(_190_),
    .B(_203_),
    .X(_204_));
 sky130_fd_sc_hd__mux2_1 _449_ (.A0(_204_),
    .A1(_202_),
    .S(net78),
    .X(_205_));
 sky130_fd_sc_hd__nor2_1 _450_ (.A(net110),
    .B(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__xnor2_1 _451_ (.A(_056_),
    .B(_205_),
    .Y(_207_));
 sky130_fd_sc_hd__a21oi_1 _452_ (.A1(net55),
    .A2(net78),
    .B1(net111),
    .Y(_208_));
 sky130_fd_sc_hd__a21o_1 _453_ (.A1(_207_),
    .A2(net77),
    .B1(_206_),
    .X(_209_));
 sky130_fd_sc_hd__nor2_1 _454_ (.A(net106),
    .B(_199_),
    .Y(_210_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(_200_),
    .B(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__a21oi_1 _456_ (.A1(_184_),
    .A2(_192_),
    .B1(net78),
    .Y(_212_));
 sky130_fd_sc_hd__o21a_1 _457_ (.A1(_184_),
    .A2(_192_),
    .B1(_212_),
    .X(_213_));
 sky130_fd_sc_hd__and3_1 _458_ (.A(_164_),
    .B(_169_),
    .C(_178_),
    .X(_214_));
 sky130_fd_sc_hd__a2111o_1 _459_ (.A1(_182_),
    .A2(_196_),
    .B1(_210_),
    .C1(_213_),
    .D1(_214_),
    .X(_215_));
 sky130_fd_sc_hd__a21oi_1 _460_ (.A1(_201_),
    .A2(_209_),
    .B1(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__xnor2_1 _461_ (.A(_207_),
    .B(net77),
    .Y(_217_));
 sky130_fd_sc_hd__mux2_1 _462_ (.A0(_217_),
    .A1(_205_),
    .S(_216_),
    .X(_218_));
 sky130_fd_sc_hd__nand2_1 _463_ (.A(net106),
    .B(_218_),
    .Y(_219_));
 sky130_fd_sc_hd__a211o_1 _464_ (.A1(_201_),
    .A2(_209_),
    .B1(_215_),
    .C1(_053_),
    .X(_220_));
 sky130_fd_sc_hd__and3_1 _465_ (.A(net55),
    .B(net111),
    .C(_196_),
    .X(_221_));
 sky130_fd_sc_hd__o32a_2 _466_ (.A1(_208_),
    .A2(net76),
    .A3(_221_),
    .B1(_220_),
    .B2(_196_),
    .X(_222_));
 sky130_fd_sc_hd__nand2_1 _467_ (.A(net109),
    .B(_222_),
    .Y(_223_));
 sky130_fd_sc_hd__and2_1 _468_ (.A(_055_),
    .B(_220_),
    .X(_224_));
 sky130_fd_sc_hd__o21bai_2 _469_ (.A1(net109),
    .A2(_222_),
    .B1_N(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__xnor2_1 _470_ (.A(_209_),
    .B(_211_),
    .Y(_226_));
 sky130_fd_sc_hd__mux2_1 _471_ (.A0(_226_),
    .A1(_199_),
    .S(_216_),
    .X(_227_));
 sky130_fd_sc_hd__inv_2 _472_ (.A(_227_),
    .Y(_228_));
 sky130_fd_sc_hd__o21ai_2 _473_ (.A1(net106),
    .A2(_218_),
    .B1(_227_),
    .Y(_229_));
 sky130_fd_sc_hd__a31oi_4 _474_ (.A1(_219_),
    .A2(_223_),
    .A3(_225_),
    .B1(_229_),
    .Y(_230_));
 sky130_fd_sc_hd__a311o_1 _475_ (.A1(_219_),
    .A2(_223_),
    .A3(_225_),
    .B1(_229_),
    .C1(_053_),
    .X(_231_));
 sky130_fd_sc_hd__or3b_1 _476_ (.A(net111),
    .B(net109),
    .C_N(_231_),
    .X(_232_));
 sky130_fd_sc_hd__nor2_1 _477_ (.A(_055_),
    .B(_220_),
    .Y(_233_));
 sky130_fd_sc_hd__o32a_1 _478_ (.A1(_224_),
    .A2(_230_),
    .A3(_233_),
    .B1(_231_),
    .B2(net76),
    .X(_234_));
 sky130_fd_sc_hd__xnor2_1 _479_ (.A(_056_),
    .B(_222_),
    .Y(_235_));
 sky130_fd_sc_hd__xnor2_1 _480_ (.A(_224_),
    .B(_235_),
    .Y(_236_));
 sky130_fd_sc_hd__mux2_1 _481_ (.A0(_236_),
    .A1(_222_),
    .S(_230_),
    .X(_237_));
 sky130_fd_sc_hd__a21oi_1 _482_ (.A1(_055_),
    .A2(_231_),
    .B1(_056_),
    .Y(_238_));
 sky130_fd_sc_hd__a221o_1 _483_ (.A1(_232_),
    .A2(_234_),
    .B1(_237_),
    .B2(net106),
    .C1(_238_),
    .X(_239_));
 sky130_fd_sc_hd__a21bo_1 _484_ (.A1(_218_),
    .A2(_227_),
    .B1_N(_230_),
    .X(_240_));
 sky130_fd_sc_hd__a22o_1 _485_ (.A1(_223_),
    .A2(_225_),
    .B1(_228_),
    .B2(_219_),
    .X(_241_));
 sky130_fd_sc_hd__a21oi_1 _486_ (.A1(_229_),
    .A2(_241_),
    .B1(_214_),
    .Y(_242_));
 sky130_fd_sc_hd__o211a_1 _487_ (.A1(net106),
    .A2(_237_),
    .B1(_240_),
    .C1(_242_),
    .X(_243_));
 sky130_fd_sc_hd__and2_1 _488_ (.A(_239_),
    .B(_243_),
    .X(_244_));
 sky130_fd_sc_hd__and4_2 _489_ (.A(net76),
    .B(_230_),
    .C(_239_),
    .D(_243_),
    .X(_245_));
 sky130_fd_sc_hd__nand2_1 _490_ (.A(net78),
    .B(_245_),
    .Y(_246_));
 sky130_fd_sc_hd__and4_1 _491_ (.A(net84),
    .B(_158_),
    .C(net78),
    .D(_245_),
    .X(_247_));
 sky130_fd_sc_hd__nand4_1 _492_ (.A(net84),
    .B(_158_),
    .C(net78),
    .D(_245_),
    .Y(_248_));
 sky130_fd_sc_hd__xnor2_1 _493_ (.A(_117_),
    .B(_247_),
    .Y(_249_));
 sky130_fd_sc_hd__xnor2_1 _494_ (.A(\tcout[7] ),
    .B(_249_),
    .Y(_250_));
 sky130_fd_sc_hd__a31o_1 _495_ (.A1(_158_),
    .A2(net78),
    .A3(_245_),
    .B1(net84),
    .X(_251_));
 sky130_fd_sc_hd__and3_1 _496_ (.A(\tcout[6] ),
    .B(_248_),
    .C(_251_),
    .X(_252_));
 sky130_fd_sc_hd__xnor2_1 _497_ (.A(_158_),
    .B(_246_),
    .Y(_253_));
 sky130_fd_sc_hd__xnor2_1 _498_ (.A(\tcout[5] ),
    .B(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__a21oi_1 _499_ (.A1(_248_),
    .A2(_251_),
    .B1(\tcout[6] ),
    .Y(_255_));
 sky130_fd_sc_hd__xor2_1 _500_ (.A(net78),
    .B(_245_),
    .X(_256_));
 sky130_fd_sc_hd__xnor2_1 _501_ (.A(\tcout[3] ),
    .B(_256_),
    .Y(_257_));
 sky130_fd_sc_hd__a21oi_1 _502_ (.A1(net78),
    .A2(_245_),
    .B1(_179_),
    .Y(_258_));
 sky130_fd_sc_hd__xnor2_1 _503_ (.A(\tcout[4] ),
    .B(_258_),
    .Y(_259_));
 sky130_fd_sc_hd__a31o_1 _504_ (.A1(_230_),
    .A2(_239_),
    .A3(_243_),
    .B1(net76),
    .X(_260_));
 sky130_fd_sc_hd__and2b_1 _505_ (.A_N(_245_),
    .B(_260_),
    .X(_261_));
 sky130_fd_sc_hd__xnor2_1 _506_ (.A(\tcout[1] ),
    .B(_230_),
    .Y(_262_));
 sky130_fd_sc_hd__nand2_1 _507_ (.A(net102),
    .B(_262_),
    .Y(_263_));
 sky130_fd_sc_hd__o21ba_1 _508_ (.A1(net102),
    .A2(_262_),
    .B1_N(_244_),
    .X(_264_));
 sky130_fd_sc_hd__a221o_1 _509_ (.A1(\tcout[8] ),
    .A2(_096_),
    .B1(_244_),
    .B2(_263_),
    .C1(_264_),
    .X(_265_));
 sky130_fd_sc_hd__xnor2_1 _510_ (.A(\tcout[2] ),
    .B(_261_),
    .Y(_266_));
 sky130_fd_sc_hd__or4_1 _511_ (.A(_257_),
    .B(_259_),
    .C(_265_),
    .D(_266_),
    .X(_267_));
 sky130_fd_sc_hd__or2_1 _512_ (.A(\tcout[8] ),
    .B(_096_),
    .X(_268_));
 sky130_fd_sc_hd__and3_1 _513_ (.A(_116_),
    .B(_247_),
    .C(_268_),
    .X(_269_));
 sky130_fd_sc_hd__a21oi_1 _514_ (.A1(_116_),
    .A2(_247_),
    .B1(_268_),
    .Y(_270_));
 sky130_fd_sc_hd__or4_1 _515_ (.A(_252_),
    .B(_255_),
    .C(_269_),
    .D(_270_),
    .X(_271_));
 sky130_fd_sc_hd__or4_4 _516_ (.A(_250_),
    .B(_254_),
    .C(_267_),
    .D(_271_),
    .X(_272_));
 sky130_fd_sc_hd__and2b_1 _517_ (.A_N(net102),
    .B(_272_),
    .X(_016_));
 sky130_fd_sc_hd__or2_1 _518_ (.A(net102),
    .B(\tcout[1] ),
    .X(_273_));
 sky130_fd_sc_hd__nand2_1 _519_ (.A(net102),
    .B(\tcout[1] ),
    .Y(_274_));
 sky130_fd_sc_hd__and3_1 _520_ (.A(_272_),
    .B(_273_),
    .C(_274_),
    .X(_017_));
 sky130_fd_sc_hd__nand3_1 _521_ (.A(net102),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .Y(_275_));
 sky130_fd_sc_hd__a21o_1 _522_ (.A1(net102),
    .A2(\tcout[1] ),
    .B1(\tcout[2] ),
    .X(_276_));
 sky130_fd_sc_hd__and3_1 _523_ (.A(_272_),
    .B(_275_),
    .C(_276_),
    .X(_018_));
 sky130_fd_sc_hd__and4_1 _524_ (.A(net102),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .D(\tcout[3] ),
    .X(_277_));
 sky130_fd_sc_hd__inv_2 _525_ (.A(_277_),
    .Y(_278_));
 sky130_fd_sc_hd__a31o_1 _526_ (.A1(net102),
    .A2(\tcout[1] ),
    .A3(\tcout[2] ),
    .B1(\tcout[3] ),
    .X(_279_));
 sky130_fd_sc_hd__and3_1 _527_ (.A(_272_),
    .B(_278_),
    .C(_279_),
    .X(_019_));
 sky130_fd_sc_hd__nand2_1 _528_ (.A(\tcout[4] ),
    .B(_277_),
    .Y(_280_));
 sky130_fd_sc_hd__or2_1 _529_ (.A(\tcout[4] ),
    .B(_277_),
    .X(_281_));
 sky130_fd_sc_hd__and3_1 _530_ (.A(_272_),
    .B(_280_),
    .C(_281_),
    .X(_020_));
 sky130_fd_sc_hd__and3_1 _531_ (.A(\tcout[4] ),
    .B(\tcout[5] ),
    .C(_277_),
    .X(_282_));
 sky130_fd_sc_hd__inv_2 _532_ (.A(_282_),
    .Y(_283_));
 sky130_fd_sc_hd__a21o_1 _533_ (.A1(\tcout[4] ),
    .A2(_277_),
    .B1(\tcout[5] ),
    .X(_284_));
 sky130_fd_sc_hd__and3_1 _534_ (.A(_272_),
    .B(_283_),
    .C(_284_),
    .X(_021_));
 sky130_fd_sc_hd__and2_1 _535_ (.A(\tcout[6] ),
    .B(_282_),
    .X(_285_));
 sky130_fd_sc_hd__nand2_1 _536_ (.A(\tcout[6] ),
    .B(_282_),
    .Y(_286_));
 sky130_fd_sc_hd__or2_1 _537_ (.A(\tcout[6] ),
    .B(_282_),
    .X(_287_));
 sky130_fd_sc_hd__and3_1 _538_ (.A(_272_),
    .B(_286_),
    .C(_287_),
    .X(_022_));
 sky130_fd_sc_hd__nand2_1 _539_ (.A(\tcout[7] ),
    .B(_285_),
    .Y(_288_));
 sky130_fd_sc_hd__or2_1 _540_ (.A(\tcout[7] ),
    .B(_285_),
    .X(_289_));
 sky130_fd_sc_hd__and3_1 _541_ (.A(_272_),
    .B(_288_),
    .C(_289_),
    .X(_023_));
 sky130_fd_sc_hd__xnor2_1 _542_ (.A(\tcout[8] ),
    .B(_288_),
    .Y(_290_));
 sky130_fd_sc_hd__and2_1 _543_ (.A(_272_),
    .B(_290_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _544_ (.A0(\sine_out_reg0[0] ),
    .A1(\sine_out_reg1[0] ),
    .S(net100),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _545_ (.A0(\sine_out_reg0[1] ),
    .A1(\sine_out_reg1[1] ),
    .S(net100),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _546_ (.A0(\sine_out_reg0[2] ),
    .A1(\sine_out_reg1[2] ),
    .S(net100),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _547_ (.A0(\sine_out_reg0[3] ),
    .A1(\sine_out_reg1[3] ),
    .S(net100),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _548_ (.A0(\sine_out_reg0[4] ),
    .A1(\sine_out_reg1[4] ),
    .S(net100),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _549_ (.A0(\sine_out_reg0[5] ),
    .A1(\sine_out_reg1[5] ),
    .S(net100),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _550_ (.A0(\sine_out_reg0[6] ),
    .A1(\sine_out_reg1[6] ),
    .S(net100),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _551_ (.A0(\sine_out_reg0[7] ),
    .A1(\sine_out_reg1[7] ),
    .S(net100),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _552_ (.A0(\sine_out_reg0[8] ),
    .A1(\sine_out_reg1[8] ),
    .S(net100),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _553_ (.A0(\sine_out_reg0[9] ),
    .A1(\sine_out_reg1[9] ),
    .S(net100),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _554_ (.A0(\sine_out_reg0[10] ),
    .A1(\sine_out_reg1[10] ),
    .S(net101),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _555_ (.A0(\sine_out_reg0[11] ),
    .A1(\sine_out_reg1[11] ),
    .S(net101),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _556_ (.A0(\sine_out_reg0[12] ),
    .A1(\sine_out_reg1[12] ),
    .S(net101),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _557_ (.A0(\sine_out_reg0[13] ),
    .A1(\sine_out_reg1[13] ),
    .S(net101),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _558_ (.A0(\sine_out_reg0[14] ),
    .A1(\sine_out_reg1[14] ),
    .S(net101),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _559_ (.A0(\sine_out_reg0[15] ),
    .A1(\sine_out_reg1[15] ),
    .S(net101),
    .X(_006_));
 sky130_fd_sc_hd__inv_2 _560_ (.A(net105),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _561_ (.A(net105),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _562_ (.A(net105),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _563_ (.A(net105),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _564_ (.A(net105),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _565_ (.A(net105),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _566_ (.A(net104),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _567_ (.A(net104),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _568_ (.A(net103),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _569_ (.A(net103),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _570_ (.A(net103),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _571_ (.A(net103),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _572_ (.A(net103),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _573_ (.A(net104),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _574_ (.A(net104),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _575_ (.A(net104),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _576_ (.A(net104),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _577_ (.A(net103),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _578_ (.A(net103),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _579_ (.A(net103),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _580_ (.A(net103),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _581_ (.A(net103),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _582_ (.A(net104),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _583_ (.A(net104),
    .Y(_049_));
 sky130_fd_sc_hd__dfrtp_1 _584_ (.CLK(clknet_3_4__leaf_clk),
    .D(_000_),
    .RESET_B(_025_),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _585_ (.CLK(clknet_3_4__leaf_clk),
    .D(_007_),
    .RESET_B(_026_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _586_ (.CLK(clknet_3_4__leaf_clk),
    .D(_008_),
    .RESET_B(_027_),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _587_ (.CLK(clknet_3_6__leaf_clk),
    .D(_009_),
    .RESET_B(_028_),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _588_ (.CLK(clknet_3_4__leaf_clk),
    .D(_010_),
    .RESET_B(_029_),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _589_ (.CLK(clknet_3_6__leaf_clk),
    .D(_011_),
    .RESET_B(_030_),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _590_ (.CLK(clknet_3_6__leaf_clk),
    .D(_012_),
    .RESET_B(_031_),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _591_ (.CLK(clknet_3_1__leaf_clk),
    .D(_013_),
    .RESET_B(_032_),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _592_ (.CLK(clknet_3_1__leaf_clk),
    .D(_014_),
    .RESET_B(_033_),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _593_ (.CLK(clknet_3_2__leaf_clk),
    .D(_015_),
    .RESET_B(_034_),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _594_ (.CLK(clknet_3_2__leaf_clk),
    .D(_001_),
    .RESET_B(_035_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _595_ (.CLK(clknet_3_2__leaf_clk),
    .D(_002_),
    .RESET_B(_036_),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _596_ (.CLK(clknet_3_2__leaf_clk),
    .D(_003_),
    .RESET_B(_037_),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _597_ (.CLK(clknet_3_3__leaf_clk),
    .D(_004_),
    .RESET_B(_038_),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _598_ (.CLK(clknet_3_2__leaf_clk),
    .D(_005_),
    .RESET_B(_039_),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_1 _599_ (.CLK(clknet_3_3__leaf_clk),
    .D(_006_),
    .RESET_B(_040_),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_4 _600_ (.CLK(clknet_3_2__leaf_clk),
    .D(_016_),
    .RESET_B(_041_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_4 _601_ (.CLK(clknet_3_2__leaf_clk),
    .D(_017_),
    .RESET_B(_042_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_4 _602_ (.CLK(clknet_3_1__leaf_clk),
    .D(_018_),
    .RESET_B(_043_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_4 _603_ (.CLK(clknet_3_1__leaf_clk),
    .D(_019_),
    .RESET_B(_044_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_4 _604_ (.CLK(clknet_3_2__leaf_clk),
    .D(_020_),
    .RESET_B(_045_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_4 _605_ (.CLK(clknet_3_1__leaf_clk),
    .D(_021_),
    .RESET_B(_046_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_4 _606_ (.CLK(clknet_3_1__leaf_clk),
    .D(_022_),
    .RESET_B(_047_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_4 _607_ (.CLK(clknet_3_1__leaf_clk),
    .D(_023_),
    .RESET_B(_048_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__dfrtp_2 _608_ (.CLK(clknet_3_1__leaf_clk),
    .D(_024_),
    .RESET_B(_049_),
    .Q(\tcout[8] ));
 sky130_fd_sc_hd__dfxtp_1 _609_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sine_out_temp0[0] ),
    .Q(\sine_out_reg0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _610_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sine_out_temp0[1] ),
    .Q(\sine_out_reg0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _611_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sine_out_temp0[2] ),
    .Q(\sine_out_reg0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _612_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sine_out_temp0[3] ),
    .Q(\sine_out_reg0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _613_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sine_out_temp0[4] ),
    .Q(\sine_out_reg0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _614_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sine_out_temp0[5] ),
    .Q(\sine_out_reg0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _615_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sine_out_temp0[6] ),
    .Q(\sine_out_reg0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _616_ (.CLK(clknet_3_7__leaf_clk),
    .D(\sine_out_temp0[7] ),
    .Q(\sine_out_reg0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _617_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sine_out_temp0[8] ),
    .Q(\sine_out_reg0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _618_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sine_out_temp0[9] ),
    .Q(\sine_out_reg0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _619_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sine_out_temp0[10] ),
    .Q(\sine_out_reg0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _620_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sine_out_temp0[11] ),
    .Q(\sine_out_reg0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _621_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sine_out_temp0[12] ),
    .Q(\sine_out_reg0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _622_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sine_out_temp0[13] ),
    .Q(\sine_out_reg0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _623_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sine_out_temp0[14] ),
    .Q(\sine_out_reg0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _624_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sine_out_temp0[15] ),
    .Q(\sine_out_reg0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _625_ (.CLK(clknet_3_5__leaf_clk),
    .D(net99),
    .Q(\sine_out_reg1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _626_ (.CLK(clknet_3_5__leaf_clk),
    .D(net94),
    .Q(\sine_out_reg1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _627_ (.CLK(clknet_3_4__leaf_clk),
    .D(net93),
    .Q(\sine_out_reg1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _628_ (.CLK(clknet_3_7__leaf_clk),
    .D(net92),
    .Q(\sine_out_reg1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _629_ (.CLK(clknet_3_5__leaf_clk),
    .D(\sine_out_temp1[4] ),
    .Q(\sine_out_reg1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _630_ (.CLK(clknet_3_7__leaf_clk),
    .D(net91),
    .Q(\sine_out_reg1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _631_ (.CLK(clknet_3_7__leaf_clk),
    .D(net90),
    .Q(\sine_out_reg1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _632_ (.CLK(clknet_3_7__leaf_clk),
    .D(net89),
    .Q(\sine_out_reg1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _633_ (.CLK(clknet_3_0__leaf_clk),
    .D(net88),
    .Q(\sine_out_reg1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _634_ (.CLK(clknet_3_0__leaf_clk),
    .D(net87),
    .Q(\sine_out_reg1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _635_ (.CLK(clknet_3_0__leaf_clk),
    .D(net98),
    .Q(\sine_out_reg1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _636_ (.CLK(clknet_3_3__leaf_clk),
    .D(\sine_out_temp1[11] ),
    .Q(\sine_out_reg1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _637_ (.CLK(clknet_3_2__leaf_clk),
    .D(net97),
    .Q(\sine_out_reg1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _638_ (.CLK(clknet_3_3__leaf_clk),
    .D(\sine_out_temp1[13] ),
    .Q(\sine_out_reg1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _639_ (.CLK(clknet_3_3__leaf_clk),
    .D(net96),
    .Q(\sine_out_reg1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _640_ (.CLK(clknet_3_3__leaf_clk),
    .D(net95),
    .Q(\sine_out_reg1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _641_ (.CLK(clknet_3_0__leaf_clk),
    .D(\tcout_delay[1] ),
    .Q(\tcout_delay[0] ));
 sky130_fd_sc_hd__dfxtp_1 _642_ (.CLK(clknet_3_1__leaf_clk),
    .D(\tcout[8] ),
    .Q(\tcout_delay[1] ));
 sky130_fd_sc_hd__conb_1 mem_i1_115 (.LO(net115));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 ram256x16 mem_i0 (.csb0(net17),
    .csb1(net114),
    .clk0(clknet_3_4__leaf_clk),
    .clk1(clknet_3_1__leaf_clk),
    .addr0({net8,
    net7,
    net6,
    net5,
    net4,
    net3,
    net2,
    net1}),
    .addr1({\tcout[7] ,
    \tcout[6] ,
    \tcout[5] ,
    \tcout[4] ,
    \tcout[3] ,
    \tcout[2] ,
    \tcout[1] ,
    net102}),
    .din0({net29,
    net28,
    net27,
    net26,
    net25,
    net24,
    net38,
    net37,
    net36,
    net35,
    net34,
    net33,
    net32,
    net31,
    net30,
    net23}),
    .dout1({\sine_out_temp0[15] ,
    \sine_out_temp0[14] ,
    \sine_out_temp0[13] ,
    \sine_out_temp0[12] ,
    \sine_out_temp0[11] ,
    \sine_out_temp0[10] ,
    \sine_out_temp0[9] ,
    \sine_out_temp0[8] ,
    \sine_out_temp0[7] ,
    \sine_out_temp0[6] ,
    \sine_out_temp0[5] ,
    \sine_out_temp0[4] ,
    \sine_out_temp0[3] ,
    \sine_out_temp0[2] ,
    \sine_out_temp0[1] ,
    \sine_out_temp0[0] }));
 ram256x16 mem_i1 (.csb0(net18),
    .csb1(net115),
    .clk0(clknet_3_5__leaf_clk),
    .clk1(clknet_3_3__leaf_clk),
    .addr0({net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net10,
    net9}),
    .addr1({\tcout[7] ,
    \tcout[6] ,
    \tcout[5] ,
    \tcout[4] ,
    \tcout[3] ,
    \tcout[2] ,
    \tcout[1] ,
    \tcout[0] }),
    .din0({net45,
    net44,
    net43,
    net42,
    net41,
    net40,
    net54,
    net53,
    net52,
    net51,
    net50,
    net49,
    net48,
    net47,
    net46,
    net39}),
    .dout1({\sine_out_temp1[15] ,
    \sine_out_temp1[14] ,
    \sine_out_temp1[13] ,
    \sine_out_temp1[12] ,
    \sine_out_temp1[11] ,
    \sine_out_temp1[10] ,
    \sine_out_temp1[9] ,
    \sine_out_temp1[8] ,
    \sine_out_temp1[7] ,
    \sine_out_temp1[6] ,
    \sine_out_temp1[5] ,
    \sine_out_temp1[4] ,
    \sine_out_temp1[3] ,
    \sine_out_temp1[2] ,
    \sine_out_temp1[1] ,
    \sine_out_temp1[0] }));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_246_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_247_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_248_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_249_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_250_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_251_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_252_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_253_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_254_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_255_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_256_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_257_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_258_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_259_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_260_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_261_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_262_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_263_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_264_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_265_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_266_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_2_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_2_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_2_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_2_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_2_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_2_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_2_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_2_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_2_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_2_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_2_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_2_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_2_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_2_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_2_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_2_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_2_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_2_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_2_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_2_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_2_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_2_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_2_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_2_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_2_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_2_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_2_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_2_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_2_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_2_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_2_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_2_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_2_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_2_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_2_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_2_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_2_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_2_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_2_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_2_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_2_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_2_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_2_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_2_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_2_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_2_Right_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_2_Right_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_2_Right_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_2_Right_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_2_Right_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_2_Right_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_2_Right_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_2_Right_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_2_Right_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_2_Right_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_2_Right_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_2_Right_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_2_Right_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_2_Right_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_2_Right_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_2_Right_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_2_Right_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_2_Right_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_2_Right_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_2_Right_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_2_Right_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_2_Right_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_2_Right_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_2_Right_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_2_Right_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_2_Right_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_2_Right_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_2_Right_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_2_Right_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_2_Right_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_2_Right_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_2_Right_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_2_Right_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_2_Right_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_2_Right_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_2_Right_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_2_Right_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_2_Right_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_2_Right_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_2_Right_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_2_Right_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_2_Right_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_2_Right_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_2_Right_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_2_Right_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_1_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_1_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_1_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_1_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_1_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_1_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_1_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_1_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_1_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_1_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_1_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_1_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_1_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_1_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_1_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_1_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_1_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_1_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_1_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_1_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_1_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_1_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_1_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_1_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_1_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_1_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_1_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_1_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_1_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_1_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_1_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_1_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_1_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_1_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_1_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_1_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_1_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_1_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_1_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_1_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_1_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_1_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_1_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_1_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_1_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_1_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_1_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_1_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_1_Left_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_1_Left_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_1_Left_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_1_Left_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_1_Left_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_1_Left_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_1_Left_459 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_1_Left_460 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_1_Left_461 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_1_Left_462 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_1_Left_463 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_1_Left_464 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_1_Left_465 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_1_Left_466 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_1_Left_467 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_1_Left_468 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_1_Left_469 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_1_Left_470 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_1_Left_471 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_1_Left_472 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_1_Left_473 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_1_Left_474 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_1_Left_475 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_1_Left_476 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_1_Left_477 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_1_Left_478 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_1_Left_479 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_1_Left_480 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_1_Left_481 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_1_Left_482 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_1_Left_483 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_1_Left_484 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_1_Left_485 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_1_Left_486 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_1_Left_487 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_1_Left_488 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_1_Left_489 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_1_Left_490 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_1_Left_491 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_1_Left_492 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_1_Left_493 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_1_Left_494 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_1_Left_495 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_1_Left_496 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_1_Left_497 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_1_Left_498 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_1_Left_499 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_1_Left_500 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_1_Left_501 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_1_Left_502 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_1_Left_503 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_1_Left_504 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_1_Left_505 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_1_Left_506 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_1_Left_507 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_1_Left_508 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_1_Left_509 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_1_Left_510 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_1_Left_511 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_246_Left_512 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_247_Left_513 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_248_Left_514 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_249_Left_515 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_250_Left_516 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_251_Left_517 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_252_Left_518 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_253_Left_519 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_254_Left_520 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_255_Left_521 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_256_Left_522 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_257_Left_523 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_258_Left_524 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_259_Left_525 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_260_Left_526 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_261_Left_527 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_262_Left_528 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_263_Left_529 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_264_Left_530 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_265_Left_531 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_266_Left_532 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_533 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_534 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_535 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_536 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_537 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_538 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_539 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_540 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_541 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_542 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_543 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_544 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_545 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_546 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_547 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_548 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_549 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_550 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_551 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_552 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_553 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_554 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_555 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_556 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_557 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_558 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_559 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_560 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_561 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_562 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_563 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_564 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_565 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_566 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_567 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_568 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_569 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_570 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_571 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_572 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_573 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_574 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_575 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_576 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_577 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_578 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_579 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_580 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_581 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_582 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_583 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_584 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_585 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_586 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_587 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_588 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_589 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_590 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_591 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_592 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_593 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_594 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_595 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_596 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_597 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_598 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_599 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_600 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_601 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_602 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_603 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_604 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_605 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_606 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_607 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_608 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_609 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_610 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_611 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_612 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_613 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_614 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_615 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_616 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_617 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_618 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_619 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Left_620 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Left_621 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Left_622 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Left_623 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Left_624 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Left_625 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Left_626 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Left_627 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Left_628 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Left_629 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Left_630 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Left_631 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Left_632 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Left_633 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Left_634 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Left_635 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Left_636 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Left_637 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Left_638 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Left_639 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Left_640 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_641 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_642 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_643 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_644 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_645 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_646 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_647 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_648 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_649 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_650 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_651 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_652 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_653 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_654 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_655 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_656 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_657 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_658 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_659 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_660 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_661 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_662 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_663 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_664 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_665 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_666 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_667 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_668 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_669 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_670 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_671 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_672 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_673 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_674 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_675 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_676 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_677 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_678 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_679 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_680 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_681 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_682 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_683 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_684 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_685 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_686 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_687 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_688 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_689 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_690 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_691 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_692 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_693 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_694 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_695 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_696 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_697 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_698 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_699 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Right_700 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Right_701 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Right_702 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Right_703 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Right_704 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Right_705 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Right_706 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Right_707 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Right_708 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Right_709 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Right_710 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Right_711 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Right_712 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Right_713 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Right_714 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Right_715 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Right_716 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Right_717 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Right_718 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Right_719 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Right_720 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Right_721 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Right_722 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Right_723 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Right_724 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Right_725 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Right_726 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Right_727 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Right_728 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Right_729 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Right_730 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Right_731 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Right_732 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Right_733 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Right_734 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Right_735 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Right_736 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Right_737 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Right_738 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Right_739 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Right_740 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Right_741 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Right_742 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Right_743 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Right_744 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Right_745 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Right_746 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_747 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Left_748 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Left_749 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Left_750 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Left_751 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Left_752 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Left_753 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Left_754 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Left_755 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Left_756 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Left_757 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Left_758 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Left_759 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Left_760 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Left_761 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Left_762 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Left_763 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Left_764 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_2_Left_765 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_2_Left_766 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_2_Left_767 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_2_Left_768 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_2_Left_769 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_2_Left_770 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_2_Left_771 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_2_Left_772 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_2_Left_773 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_2_Left_774 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_2_Left_775 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_2_Left_776 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_2_Left_777 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_2_Left_778 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_2_Left_779 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_2_Left_780 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_2_Left_781 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_2_Left_782 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_2_Left_783 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_2_Left_784 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_2_Left_785 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_2_Left_786 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_2_Left_787 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_2_Left_788 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_2_Left_789 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_2_Left_790 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_2_Left_791 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_2_Left_792 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_2_Left_793 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_2_Left_794 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_2_Left_795 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_2_Left_796 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_2_Left_797 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_2_Left_798 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_2_Left_799 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_2_Left_800 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_2_Left_801 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_2_Left_802 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_2_Left_803 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_2_Left_804 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_2_Left_805 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_2_Left_806 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_2_Left_807 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_2_Left_808 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_2_Left_809 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_2_Left_810 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_2_Left_811 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_2_Left_812 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_2_Left_813 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_2_Left_814 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_2_Left_815 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_2_Left_816 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_2_Left_817 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_2_Left_818 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_2_Left_819 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_2_Left_820 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_2_Left_821 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_2_Left_822 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_2_Left_823 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_2_Left_824 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_2_Left_825 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_2_Left_826 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_2_Left_827 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_2_Left_828 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_2_Left_829 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_2_Left_830 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_2_Left_831 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_2_Left_832 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_2_Left_833 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_2_Left_834 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_2_Left_835 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_2_Left_836 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_2_Left_837 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_2_Left_838 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_2_Left_839 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_2_Left_840 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_2_Left_841 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_2_Left_842 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_2_Left_843 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_2_Left_844 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_2_Left_845 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_2_Left_846 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_2_Left_847 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_2_Left_848 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_2_Left_849 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_2_Left_850 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_2_Left_851 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_2_Left_852 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_2_Left_853 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_2_Left_854 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_1_Right_855 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_1_Right_856 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_1_Right_857 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_1_Right_858 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_1_Right_859 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_1_Right_860 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_1_Right_861 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_1_Right_862 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_1_Right_863 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_1_Right_864 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_1_Right_865 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_1_Right_866 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_1_Right_867 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_1_Right_868 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_1_Right_869 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_1_Right_870 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_1_Right_871 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_1_Right_872 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_1_Right_873 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_1_Right_874 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_1_Right_875 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_1_Right_876 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_1_Right_877 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_1_Right_878 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_1_Right_879 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_1_Right_880 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_1_Right_881 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_1_Right_882 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_1_Right_883 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_1_Right_884 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_1_Right_885 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_1_Right_886 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_1_Right_887 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_1_Right_888 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_1_Right_889 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_1_Right_890 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_1_Right_891 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_1_Right_892 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_1_Right_893 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_1_Right_894 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_1_Right_895 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_1_Right_896 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_1_Right_897 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_1_Right_898 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_1_Right_899 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_1_Right_900 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_1_Right_901 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_1_Right_902 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_1_Right_903 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_1_Right_904 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_1_Right_905 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_1_Right_906 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_1_Right_907 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_1_Right_908 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_1_Right_909 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_1_Right_910 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_1_Right_911 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_1_Right_912 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_1_Right_913 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_1_Right_914 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_1_Right_915 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_1_Right_916 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_1_Right_917 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_1_Right_918 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_1_Right_919 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_1_Right_920 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_1_Right_921 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_1_Right_922 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_1_Right_923 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_1_Right_924 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_1_Right_925 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_1_Right_926 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_1_Right_927 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_1_Right_928 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_1_Right_929 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_1_Right_930 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_1_Right_931 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_1_Right_932 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_1_Right_933 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_1_Right_934 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_1_Right_935 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_1_Right_936 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_1_Right_937 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_1_Right_938 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_1_Right_939 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_1_Right_940 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_1_Right_941 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_1_Right_942 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_1_Right_943 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_1_Right_944 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_1_Right_945 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_230_1_Right_946 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_231_1_Right_947 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_232_1_Right_948 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_233_1_Right_949 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_234_1_Right_950 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_235_1_Right_951 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_236_1_Right_952 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_237_1_Right_953 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_238_1_Right_954 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_239_1_Right_955 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_240_1_Right_956 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_241_1_Right_957 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_242_1_Right_958 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_243_1_Right_959 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_244_1_Right_960 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_245_1_Right_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_1_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_1_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_1_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_1_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_1_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_1_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_1_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_1_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_1_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_1_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_1_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_1_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_1_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_1_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_1_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_1_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_253_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_254_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_255_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_256_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_257_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_258_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_259_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_260_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_261_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_262_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_263_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_264_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_265_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_266_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_2_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_2_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_2_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_2_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_2_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_2_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_2_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_2_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_2_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_2_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_2_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_2_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_2_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_2_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_2_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_2_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_2_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_2_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_2_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_2_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_2_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_2_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_2_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_2_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_2_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_2_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_2_2491 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(addr00[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(addr00[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(addr00[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(addr00[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(addr00[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(addr00[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(addr00[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(addr00[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(addr01[0]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(addr01[1]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(addr01[2]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(addr01[3]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(addr01[4]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(addr01[5]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(addr01[6]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(addr01[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(csb00),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(csb01),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(denum[0]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(denum[1]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(denum[2]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(denum[3]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(din00[0]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(din00[10]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(din00[11]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(din00[12]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(din00[13]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(din00[14]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(din00[15]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(din00[1]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(din00[2]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(din00[3]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(din00[4]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(din00[5]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(din00[6]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(din00[7]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(din00[8]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(din00[9]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(din01[0]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(din01[10]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(din01[11]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(din01[12]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(din01[13]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(din01[14]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(din01[15]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(din01[1]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(din01[2]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(din01[3]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(din01[4]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(din01[5]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(din01[6]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(din01[7]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(din01[8]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(din01[9]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(num[0]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(num[1]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(num[2]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(num[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(rst),
    .X(net59));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(sine_out[0]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(sine_out[10]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(sine_out[11]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(sine_out[12]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(sine_out[13]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(sine_out[14]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(sine_out[15]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(sine_out[1]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(sine_out[2]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(sine_out[3]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(sine_out[4]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(sine_out[5]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(sine_out[6]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(sine_out[7]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(sine_out[8]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(sine_out[9]));
 sky130_fd_sc_hd__clkbuf_2 max_cap76 (.A(_216_),
    .X(net76));
 sky130_fd_sc_hd__buf_1 max_cap77 (.A(_208_),
    .X(net77));
 sky130_fd_sc_hd__buf_2 fanout78 (.A(_196_),
    .X(net78));
 sky130_fd_sc_hd__buf_1 max_cap79 (.A(_175_),
    .X(net79));
 sky130_fd_sc_hd__buf_1 max_cap80 (.A(_176_),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 wire81 (.A(net83),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 max_cap82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 wire83 (.A(_144_),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 max_cap84 (.A(_139_),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 max_cap85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 max_cap86 (.A(_086_),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 wire87 (.A(\sine_out_temp1[9] ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 wire88 (.A(\sine_out_temp1[8] ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 wire89 (.A(\sine_out_temp1[7] ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 wire90 (.A(\sine_out_temp1[6] ),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 wire91 (.A(\sine_out_temp1[5] ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 wire92 (.A(\sine_out_temp1[3] ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 wire93 (.A(\sine_out_temp1[2] ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 wire94 (.A(\sine_out_temp1[1] ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 wire95 (.A(\sine_out_temp1[15] ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 wire96 (.A(\sine_out_temp1[14] ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 wire97 (.A(\sine_out_temp1[12] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 wire98 (.A(\sine_out_temp1[10] ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 wire99 (.A(\sine_out_temp1[0] ),
    .X(net99));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(\tcout_delay[0] ),
    .X(net100));
 sky130_fd_sc_hd__buf_2 fanout101 (.A(\tcout_delay[0] ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(\tcout[0] ),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_4 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(net59),
    .X(net105));
 sky130_fd_sc_hd__buf_2 fanout106 (.A(net108),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(net58),
    .X(net107));
 sky130_fd_sc_hd__buf_1 fanout108 (.A(net58),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net57),
    .X(net110));
 sky130_fd_sc_hd__buf_2 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_2 fanout112 (.A(net56),
    .X(net112));
 sky130_fd_sc_hd__buf_2 fanout113 (.A(net55),
    .X(net113));
 sky130_fd_sc_hd__conb_1 mem_i0_114 (.LO(net114));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_3_7__leaf_clk));
endmodule
