magic
tech sky130A
magscale 1 2
timestamp 1741712758
<< viali >>
rect 55597 97257 55631 97291
rect 57989 97257 58023 97291
rect 58817 97257 58851 97291
rect 60105 97257 60139 97291
rect 60749 97257 60783 97291
rect 62681 97257 62715 97291
rect 63325 97257 63359 97291
rect 64613 97257 64647 97291
rect 65257 97257 65291 97291
rect 67189 97189 67223 97223
rect 67833 97189 67867 97223
rect 70501 97189 70535 97223
rect 71697 97189 71731 97223
rect 72341 97189 72375 97223
rect 74365 97189 74399 97223
rect 107485 97189 107519 97223
rect 55781 97053 55815 97087
rect 58173 97053 58207 97087
rect 59001 97053 59035 97087
rect 60289 97053 60323 97087
rect 60933 97053 60967 97087
rect 62865 97053 62899 97087
rect 63509 97053 63543 97087
rect 64797 97053 64831 97087
rect 65441 97053 65475 97087
rect 67373 97053 67407 97087
rect 68017 97053 68051 97087
rect 69949 97053 69983 97087
rect 70317 97053 70351 97087
rect 71881 97053 71915 97087
rect 72525 97053 72559 97087
rect 74181 97053 74215 97087
rect 107669 97053 107703 97087
rect 57621 96985 57655 97019
rect 58265 96985 58299 97019
rect 68201 96985 68235 97019
rect 56149 96917 56183 96951
rect 67649 96917 67683 96951
rect 107853 96917 107887 96951
rect 108037 96917 108071 96951
rect 56241 96645 56275 96679
rect 69305 96577 69339 96611
rect 69121 96441 69155 96475
rect 58541 96169 58575 96203
rect 67833 96169 67867 96203
rect 73445 96169 73479 96203
rect 56793 96033 56827 96067
rect 66085 96033 66119 96067
rect 71697 95965 71731 95999
rect 57069 95897 57103 95931
rect 66361 95897 66395 95931
rect 71973 95897 72007 95931
rect 57437 95625 57471 95659
rect 61025 95625 61059 95659
rect 62865 95625 62899 95659
rect 64981 95625 65015 95659
rect 66821 95625 66855 95659
rect 71789 95625 71823 95659
rect 55965 95557 55999 95591
rect 59553 95557 59587 95591
rect 68201 95489 68235 95523
rect 70041 95489 70075 95523
rect 55689 95421 55723 95455
rect 59277 95421 59311 95455
rect 61117 95421 61151 95455
rect 61393 95421 61427 95455
rect 63233 95421 63267 95455
rect 63509 95421 63543 95455
rect 65073 95421 65107 95455
rect 65349 95421 65383 95455
rect 68477 95421 68511 95455
rect 70317 95421 70351 95455
rect 69949 95353 69983 95387
rect 59645 95081 59679 95115
rect 63785 95081 63819 95115
rect 67373 95081 67407 95115
rect 69213 95081 69247 95115
rect 72525 95081 72559 95115
rect 56057 94945 56091 94979
rect 57897 94945 57931 94979
rect 62037 94945 62071 94979
rect 65625 94945 65659 94979
rect 67465 94945 67499 94979
rect 70777 94877 70811 94911
rect 56241 94809 56275 94843
rect 58173 94809 58207 94843
rect 62313 94809 62347 94843
rect 65901 94809 65935 94843
rect 67741 94809 67775 94843
rect 71053 94809 71087 94843
rect 56333 94741 56367 94775
rect 56701 94741 56735 94775
rect 55321 94537 55355 94571
rect 58357 94537 58391 94571
rect 61301 94537 61335 94571
rect 61761 94537 61795 94571
rect 65349 94537 65383 94571
rect 59369 94469 59403 94503
rect 54953 94401 54987 94435
rect 55597 94401 55631 94435
rect 55864 94401 55898 94435
rect 58449 94401 58483 94435
rect 59461 94401 59495 94435
rect 59553 94401 59587 94435
rect 61853 94401 61887 94435
rect 64153 94401 64187 94435
rect 65441 94401 65475 94435
rect 54677 94333 54711 94367
rect 54861 94333 54895 94367
rect 58173 94333 58207 94367
rect 59829 94333 59863 94367
rect 58817 94265 58851 94299
rect 64429 94265 64463 94299
rect 55505 94197 55539 94231
rect 56977 94197 57011 94231
rect 63877 94197 63911 94231
rect 57805 93993 57839 94027
rect 60013 93993 60047 94027
rect 64153 93993 64187 94027
rect 66361 93993 66395 94027
rect 69949 93993 69983 94027
rect 55597 93925 55631 93959
rect 59461 93857 59495 93891
rect 60565 93857 60599 93891
rect 61577 93857 61611 93891
rect 62405 93857 62439 93891
rect 63601 93857 63635 93891
rect 64521 93857 64555 93891
rect 65717 93857 65751 93891
rect 57161 93789 57195 93823
rect 59185 93789 59219 93823
rect 59645 93789 59679 93823
rect 60289 93789 60323 93823
rect 60749 93789 60783 93823
rect 62589 93789 62623 93823
rect 63141 93789 63175 93823
rect 63233 93789 63267 93823
rect 63785 93789 63819 93823
rect 64613 93789 64647 93823
rect 65257 93789 65291 93823
rect 65349 93789 65383 93823
rect 65901 93789 65935 93823
rect 66637 93789 66671 93823
rect 67097 93789 67131 93823
rect 67189 93789 67223 93823
rect 68385 93789 68419 93823
rect 68661 93789 68695 93823
rect 68753 93789 68787 93823
rect 69121 93789 69155 93823
rect 69213 93789 69247 93823
rect 70041 93789 70075 93823
rect 70961 93789 70995 93823
rect 56916 93721 56950 93755
rect 58940 93721 58974 93755
rect 60197 93721 60231 93755
rect 60841 93721 60875 93755
rect 70317 93721 70351 93755
rect 70501 93721 70535 93755
rect 54677 93653 54711 93687
rect 55781 93653 55815 93687
rect 59553 93653 59587 93687
rect 61209 93653 61243 93687
rect 61669 93653 61703 93687
rect 61761 93653 61795 93687
rect 62129 93653 62163 93687
rect 62497 93653 62531 93687
rect 62957 93653 62991 93687
rect 63693 93653 63727 93687
rect 64705 93653 64739 93687
rect 65073 93653 65107 93687
rect 65993 93653 66027 93687
rect 66545 93653 66579 93687
rect 68845 93653 68879 93687
rect 70869 93653 70903 93687
rect 71145 93653 71179 93687
rect 72249 93653 72283 93687
rect 54493 93449 54527 93483
rect 57713 93449 57747 93483
rect 60013 93449 60047 93483
rect 61485 93449 61519 93483
rect 63417 93449 63451 93483
rect 66637 93449 66671 93483
rect 72709 93449 72743 93483
rect 72985 93449 73019 93483
rect 74733 93449 74767 93483
rect 54033 93381 54067 93415
rect 70225 93381 70259 93415
rect 72249 93381 72283 93415
rect 72433 93381 72467 93415
rect 46121 93313 46155 93347
rect 49781 93313 49815 93347
rect 54125 93313 54159 93347
rect 54677 93313 54711 93347
rect 56609 93313 56643 93347
rect 57345 93313 57379 93347
rect 59665 93313 59699 93347
rect 59921 93313 59955 93347
rect 61137 93313 61171 93347
rect 61393 93313 61427 93347
rect 62609 93313 62643 93347
rect 62865 93313 62899 93347
rect 63233 93313 63267 93347
rect 63325 93313 63359 93347
rect 64541 93313 64575 93347
rect 64797 93313 64831 93347
rect 66013 93313 66047 93347
rect 66269 93313 66303 93347
rect 66729 93313 66763 93347
rect 68569 93313 68603 93347
rect 69397 93313 69431 93347
rect 70317 93313 70351 93347
rect 71901 93313 71935 93347
rect 72617 93313 72651 93347
rect 73077 93313 73111 93347
rect 73445 93313 73479 93347
rect 73629 93313 73663 93347
rect 73905 93313 73939 93347
rect 74457 93313 74491 93347
rect 74825 93313 74859 93347
rect 46305 93245 46339 93279
rect 46949 93245 46983 93279
rect 47133 93245 47167 93279
rect 49249 93245 49283 93279
rect 49525 93245 49559 93279
rect 53849 93245 53883 93279
rect 56425 93245 56459 93279
rect 57069 93245 57103 93279
rect 57253 93245 57287 93279
rect 66453 93245 66487 93279
rect 68385 93245 68419 93279
rect 68477 93245 68511 93279
rect 69121 93245 69155 93279
rect 69305 93245 69339 93279
rect 70133 93245 70167 93279
rect 72157 93245 72191 93279
rect 75193 93245 75227 93279
rect 49341 93177 49375 93211
rect 50905 93177 50939 93211
rect 58541 93177 58575 93211
rect 67097 93177 67131 93211
rect 70777 93177 70811 93211
rect 75009 93177 75043 93211
rect 64889 93109 64923 93143
rect 68937 93109 68971 93143
rect 69765 93109 69799 93143
rect 70685 93109 70719 93143
rect 75377 93109 75411 93143
rect 46949 92905 46983 92939
rect 48421 92905 48455 92939
rect 52193 92905 52227 92939
rect 53665 92905 53699 92939
rect 55137 92905 55171 92939
rect 56517 92905 56551 92939
rect 59553 92905 59587 92939
rect 63509 92905 63543 92939
rect 65625 92905 65659 92939
rect 67097 92905 67131 92939
rect 70777 92905 70811 92939
rect 72249 92905 72283 92939
rect 68569 92837 68603 92871
rect 47041 92769 47075 92803
rect 50629 92769 50663 92803
rect 57989 92769 58023 92803
rect 63601 92769 63635 92803
rect 45569 92701 45603 92735
rect 50813 92701 50847 92735
rect 52285 92701 52319 92735
rect 53757 92701 53791 92735
rect 55505 92701 55539 92735
rect 57897 92701 57931 92735
rect 58173 92701 58207 92735
rect 61945 92701 61979 92735
rect 67005 92701 67039 92735
rect 68477 92701 68511 92735
rect 69949 92701 69983 92735
rect 72157 92701 72191 92735
rect 73629 92701 73663 92735
rect 45385 92633 45419 92667
rect 45814 92633 45848 92667
rect 47286 92633 47320 92667
rect 48513 92633 48547 92667
rect 51058 92633 51092 92667
rect 52552 92633 52586 92667
rect 54024 92633 54058 92667
rect 57652 92633 57686 92667
rect 58440 92633 58474 92667
rect 61761 92633 61795 92667
rect 62190 92633 62224 92667
rect 63846 92633 63880 92667
rect 66760 92633 66794 92667
rect 68232 92633 68266 92667
rect 69704 92633 69738 92667
rect 71912 92633 71946 92667
rect 73384 92633 73418 92667
rect 77401 92633 77435 92667
rect 77493 92633 77527 92667
rect 79241 92633 79275 92667
rect 55321 92565 55355 92599
rect 63325 92565 63359 92599
rect 64981 92565 65015 92599
rect 73813 92565 73847 92599
rect 79425 92565 79459 92599
rect 45661 92361 45695 92395
rect 47133 92361 47167 92395
rect 54769 92361 54803 92395
rect 60289 92361 60323 92395
rect 63509 92361 63543 92395
rect 65073 92361 65107 92395
rect 65349 92361 65383 92395
rect 72985 92361 73019 92395
rect 47317 92293 47351 92327
rect 47961 92293 47995 92327
rect 56578 92293 56612 92327
rect 64981 92293 65015 92327
rect 69428 92293 69462 92327
rect 70961 92293 70995 92327
rect 72801 92293 72835 92327
rect 46949 92225 46983 92259
rect 48237 92225 48271 92259
rect 48493 92225 48527 92259
rect 49985 92225 50019 92259
rect 50445 92225 50479 92259
rect 50701 92225 50735 92259
rect 53389 92225 53423 92259
rect 53645 92225 53679 92259
rect 56149 92225 56183 92259
rect 56333 92225 56367 92259
rect 58909 92225 58943 92259
rect 59165 92225 59199 92259
rect 60749 92225 60783 92259
rect 61005 92225 61039 92259
rect 69673 92225 69707 92259
rect 70317 92225 70351 92259
rect 74477 92225 74511 92259
rect 74733 92225 74767 92259
rect 74917 92225 74951 92259
rect 77677 92225 77711 92259
rect 50261 92089 50295 92123
rect 51825 92089 51859 92123
rect 58725 92089 58759 92123
rect 60565 92089 60599 92123
rect 62129 92089 62163 92123
rect 68293 92089 68327 92123
rect 71329 92089 71363 92123
rect 73353 92089 73387 92123
rect 100125 92089 100159 92123
rect 48053 92021 48087 92055
rect 49617 92021 49651 92055
rect 53205 92021 53239 92055
rect 57713 92021 57747 92055
rect 77953 92021 77987 92055
rect 89453 92021 89487 92055
rect 108313 86581 108347 86615
rect 108405 67337 108439 67371
rect 109877 67337 109911 67371
rect 109529 67201 109563 67235
rect 109785 67133 109819 67167
rect 110061 66997 110095 67031
rect 108313 57885 108347 57919
rect 109969 57885 110003 57919
rect 108580 57817 108614 57851
rect 109785 57817 109819 57851
rect 109693 57749 109727 57783
rect 108589 54825 108623 54859
rect 108313 54621 108347 54655
rect 108405 54553 108439 54587
rect 108313 54281 108347 54315
rect 108313 53533 108347 53567
rect 110061 53465 110095 53499
rect 110245 53397 110279 53431
rect 109049 53193 109083 53227
rect 108773 53057 108807 53091
rect 108313 52513 108347 52547
rect 110521 52445 110555 52479
rect 108589 52377 108623 52411
rect 110337 52377 110371 52411
rect 108313 52105 108347 52139
rect 109325 52037 109359 52071
rect 109601 52037 109635 52071
rect 109049 51969 109083 52003
rect 108313 51357 108347 51391
rect 109601 51221 109635 51255
rect 108773 50949 108807 50983
rect 108865 50881 108899 50915
rect 109141 50881 109175 50915
rect 108957 50677 108991 50711
rect 108681 50473 108715 50507
rect 108313 50269 108347 50303
rect 108405 50201 108439 50235
rect 108957 49385 108991 49419
rect 108681 49317 108715 49351
rect 109141 49317 109175 49351
rect 108313 49181 108347 49215
rect 108405 49113 108439 49147
rect 109417 49113 109451 49147
rect 110337 48161 110371 48195
rect 110061 48025 110095 48059
rect 108589 47957 108623 47991
rect 108681 47209 108715 47243
rect 110705 47209 110739 47243
rect 110429 47073 110463 47107
rect 110153 46937 110187 46971
rect 109233 46529 109267 46563
rect 109693 46325 109727 46359
rect 110429 45985 110463 46019
rect 108313 45917 108347 45951
rect 110153 45849 110187 45883
rect 108405 45781 108439 45815
rect 108681 45781 108715 45815
rect 108313 45577 108347 45611
rect 109217 45509 109251 45543
rect 109417 45509 109451 45543
rect 110613 45509 110647 45543
rect 108773 45441 108807 45475
rect 110337 45441 110371 45475
rect 110429 45441 110463 45475
rect 109049 45305 109083 45339
rect 110797 45305 110831 45339
rect 108957 45237 108991 45271
rect 109233 45237 109267 45271
rect 109785 45237 109819 45271
rect 109509 45033 109543 45067
rect 109417 44829 109451 44863
rect 109601 44829 109635 44863
rect 1409 44353 1443 44387
rect 1685 44353 1719 44387
rect 108313 44353 108347 44387
rect 108589 44353 108623 44387
rect 1593 44217 1627 44251
rect 108405 44217 108439 44251
rect 108589 43945 108623 43979
rect 109601 43945 109635 43979
rect 110245 43945 110279 43979
rect 110429 43945 110463 43979
rect 109969 43809 110003 43843
rect 108313 43741 108347 43775
rect 109785 43741 109819 43775
rect 108405 43673 108439 43707
rect 110061 43673 110095 43707
rect 110261 43605 110295 43639
rect 109601 43401 109635 43435
rect 109509 43333 109543 43367
rect 1409 43265 1443 43299
rect 1685 43265 1719 43299
rect 109325 43265 109359 43299
rect 109601 43265 109635 43299
rect 109693 43265 109727 43299
rect 109969 43265 110003 43299
rect 110429 43265 110463 43299
rect 1593 43129 1627 43163
rect 110245 43129 110279 43163
rect 109877 43061 109911 43095
rect 110153 43061 110187 43095
rect 108681 42857 108715 42891
rect 109877 42857 109911 42891
rect 108405 42653 108439 42687
rect 109417 42653 109451 42687
rect 109509 42653 109543 42687
rect 109693 42653 109727 42687
rect 108497 42517 108531 42551
rect 110337 42177 110371 42211
rect 110061 42109 110095 42143
rect 108589 41973 108623 42007
rect 108589 41769 108623 41803
rect 109969 41769 110003 41803
rect 109601 41633 109635 41667
rect 108313 41565 108347 41599
rect 109417 41565 109451 41599
rect 109693 41565 109727 41599
rect 110705 41565 110739 41599
rect 110889 41565 110923 41599
rect 108405 41429 108439 41463
rect 110797 41429 110831 41463
rect 1409 41089 1443 41123
rect 1685 41089 1719 41123
rect 109969 41089 110003 41123
rect 110429 41089 110463 41123
rect 110613 41089 110647 41123
rect 110889 41089 110923 41123
rect 1593 40953 1627 40987
rect 110153 40885 110187 40919
rect 111073 40885 111107 40919
rect 110153 40681 110187 40715
rect 110337 40681 110371 40715
rect 110705 40613 110739 40647
rect 108313 40545 108347 40579
rect 110981 40545 111015 40579
rect 1409 40477 1443 40511
rect 1685 40477 1719 40511
rect 111073 40477 111107 40511
rect 108589 40409 108623 40443
rect 110521 40409 110555 40443
rect 1593 40341 1627 40375
rect 110061 40341 110095 40375
rect 110311 40341 110345 40375
rect 109969 40137 110003 40171
rect 110429 40137 110463 40171
rect 110889 40069 110923 40103
rect 109509 40001 109543 40035
rect 109601 40001 109635 40035
rect 109693 40001 109727 40035
rect 109785 40001 109819 40035
rect 110061 40001 110095 40035
rect 110613 40001 110647 40035
rect 110761 40001 110795 40035
rect 110981 40001 111015 40035
rect 111119 40001 111153 40035
rect 110245 39797 110279 39831
rect 111257 39797 111291 39831
rect 110705 39593 110739 39627
rect 110245 39457 110279 39491
rect 110521 39389 110555 39423
rect 109969 39321 110003 39355
rect 108497 39253 108531 39287
rect 110337 39253 110371 39287
rect 109509 39049 109543 39083
rect 110337 39049 110371 39083
rect 110613 39049 110647 39083
rect 109693 38981 109727 39015
rect 109877 38981 109911 39015
rect 110981 38981 111015 39015
rect 109601 38913 109635 38947
rect 109969 38913 110003 38947
rect 110245 38913 110279 38947
rect 111165 38913 111199 38947
rect 109325 38777 109359 38811
rect 110153 38709 110187 38743
rect 110797 38709 110831 38743
rect 111717 38505 111751 38539
rect 110337 38369 110371 38403
rect 1409 38301 1443 38335
rect 1685 38301 1719 38335
rect 111901 38301 111935 38335
rect 112085 38301 112119 38335
rect 110061 38233 110095 38267
rect 1593 38165 1627 38199
rect 108589 38165 108623 38199
rect 109141 37961 109175 37995
rect 109785 37961 109819 37995
rect 109309 37893 109343 37927
rect 109509 37893 109543 37927
rect 1409 37825 1443 37859
rect 1685 37825 1719 37859
rect 110429 37825 110463 37859
rect 110705 37825 110739 37859
rect 112545 37825 112579 37859
rect 113465 37825 113499 37859
rect 113925 37825 113959 37859
rect 114569 37825 114603 37859
rect 110061 37757 110095 37791
rect 110797 37757 110831 37791
rect 112269 37757 112303 37791
rect 112361 37757 112395 37791
rect 112453 37757 112487 37791
rect 113833 37757 113867 37791
rect 1593 37689 1627 37723
rect 111073 37689 111107 37723
rect 109325 37621 109359 37655
rect 110153 37621 110187 37655
rect 110291 37621 110325 37655
rect 112085 37621 112119 37655
rect 114109 37621 114143 37655
rect 114477 37621 114511 37655
rect 109325 37417 109359 37451
rect 109509 37417 109543 37451
rect 111073 37417 111107 37451
rect 111257 37349 111291 37383
rect 112821 37349 112855 37383
rect 113281 37349 113315 37383
rect 109693 37281 109727 37315
rect 116409 37281 116443 37315
rect 109877 37213 109911 37247
rect 112637 37213 112671 37247
rect 113557 37213 113591 37247
rect 113925 37213 113959 37247
rect 114293 37213 114327 37247
rect 114385 37213 114419 37247
rect 115121 37213 115155 37247
rect 115305 37213 115339 37247
rect 109141 37145 109175 37179
rect 111533 37145 111567 37179
rect 112269 37145 112303 37179
rect 114753 37145 114787 37179
rect 114845 37145 114879 37179
rect 109341 37077 109375 37111
rect 112453 37077 112487 37111
rect 112545 37077 112579 37111
rect 115857 37077 115891 37111
rect 116225 37077 116259 37111
rect 116317 37077 116351 37111
rect 110245 36873 110279 36907
rect 113281 36873 113315 36907
rect 114569 36873 114603 36907
rect 114753 36873 114787 36907
rect 116225 36873 116259 36907
rect 111165 36805 111199 36839
rect 112361 36805 112395 36839
rect 114201 36805 114235 36839
rect 115121 36805 115155 36839
rect 115489 36805 115523 36839
rect 110061 36737 110095 36771
rect 112453 36737 112487 36771
rect 113557 36737 113591 36771
rect 113649 36737 113683 36771
rect 113741 36737 113775 36771
rect 113925 36737 113959 36771
rect 114017 36737 114051 36771
rect 114293 36737 114327 36771
rect 114385 36737 114419 36771
rect 114661 36737 114695 36771
rect 114937 36737 114971 36771
rect 115029 36737 115063 36771
rect 115213 36737 115247 36771
rect 115882 36737 115916 36771
rect 116317 36737 116351 36771
rect 116501 36737 116535 36771
rect 116685 36737 116719 36771
rect 116777 36737 116811 36771
rect 116961 36737 116995 36771
rect 109785 36669 109819 36703
rect 110797 36669 110831 36703
rect 111018 36669 111052 36703
rect 112269 36669 112303 36703
rect 115765 36669 115799 36703
rect 116961 36601 116995 36635
rect 108313 36533 108347 36567
rect 110705 36533 110739 36567
rect 110889 36533 110923 36567
rect 112821 36533 112855 36567
rect 114937 36533 114971 36567
rect 115397 36533 115431 36567
rect 109325 36329 109359 36363
rect 109509 36329 109543 36363
rect 110797 36329 110831 36363
rect 111809 36329 111843 36363
rect 114477 36329 114511 36363
rect 115581 36329 115615 36363
rect 116593 36329 116627 36363
rect 116961 36329 116995 36363
rect 113005 36261 113039 36295
rect 116409 36261 116443 36295
rect 110981 36193 111015 36227
rect 113373 36193 113407 36227
rect 113649 36193 113683 36227
rect 113741 36193 113775 36227
rect 115029 36193 115063 36227
rect 116501 36193 116535 36227
rect 110153 36125 110187 36159
rect 110337 36125 110371 36159
rect 111073 36125 111107 36159
rect 111988 36125 112022 36159
rect 112360 36125 112394 36159
rect 112453 36125 112487 36159
rect 112545 36125 112579 36159
rect 112913 36125 112947 36159
rect 113189 36125 113223 36159
rect 113557 36125 113591 36159
rect 113833 36125 113867 36159
rect 114017 36125 114051 36159
rect 115305 36125 115339 36159
rect 115857 36125 115891 36159
rect 116041 36125 116075 36159
rect 116869 36125 116903 36159
rect 116961 36125 116995 36159
rect 117145 36125 117179 36159
rect 109141 36057 109175 36091
rect 112085 36057 112119 36091
rect 112177 36057 112211 36091
rect 115581 36057 115615 36091
rect 116133 36057 116167 36091
rect 109341 35989 109375 36023
rect 114845 35989 114879 36023
rect 114937 35989 114971 36023
rect 115397 35989 115431 36023
rect 115857 35989 115891 36023
rect 116777 35989 116811 36023
rect 1593 35785 1627 35819
rect 108773 35785 108807 35819
rect 109233 35785 109267 35819
rect 109325 35785 109359 35819
rect 111901 35785 111935 35819
rect 113373 35785 113407 35819
rect 114753 35785 114787 35819
rect 116961 35785 116995 35819
rect 117145 35785 117179 35819
rect 117421 35785 117455 35819
rect 108865 35717 108899 35751
rect 109065 35717 109099 35751
rect 113005 35717 113039 35751
rect 113649 35717 113683 35751
rect 117973 35717 118007 35751
rect 1409 35649 1443 35683
rect 1685 35649 1719 35683
rect 108589 35649 108623 35683
rect 108773 35649 108807 35683
rect 109509 35649 109543 35683
rect 109693 35649 109727 35683
rect 109969 35649 110003 35683
rect 110429 35649 110463 35683
rect 111073 35649 111107 35683
rect 111533 35649 111567 35683
rect 112913 35649 112947 35683
rect 113097 35649 113131 35683
rect 113557 35649 113591 35683
rect 113741 35649 113775 35683
rect 113925 35649 113959 35683
rect 114017 35649 114051 35683
rect 114385 35649 114419 35683
rect 115213 35649 115247 35683
rect 115305 35649 115339 35683
rect 115489 35649 115523 35683
rect 115581 35649 115615 35683
rect 116593 35649 116627 35683
rect 117329 35649 117363 35683
rect 117605 35649 117639 35683
rect 118157 35649 118191 35683
rect 118249 35649 118283 35683
rect 110521 35581 110555 35615
rect 110797 35581 110831 35615
rect 111625 35581 111659 35615
rect 114477 35581 114511 35615
rect 116409 35581 116443 35615
rect 116501 35581 116535 35615
rect 117881 35581 117915 35615
rect 110889 35513 110923 35547
rect 117973 35513 118007 35547
rect 109049 35445 109083 35479
rect 109785 35445 109819 35479
rect 115029 35445 115063 35479
rect 117789 35445 117823 35479
rect 109233 35241 109267 35275
rect 111625 35241 111659 35275
rect 112269 35241 112303 35275
rect 112821 35241 112855 35275
rect 114109 35241 114143 35275
rect 114937 35241 114971 35275
rect 116501 35241 116535 35275
rect 117329 35241 117363 35275
rect 118525 35241 118559 35275
rect 110337 35173 110371 35207
rect 112637 35173 112671 35207
rect 115029 35173 115063 35207
rect 110061 35105 110095 35139
rect 111441 35105 111475 35139
rect 113741 35105 113775 35139
rect 113833 35105 113867 35139
rect 115581 35105 115615 35139
rect 116133 35105 116167 35139
rect 117605 35105 117639 35139
rect 109325 35037 109359 35071
rect 109969 35037 110003 35071
rect 111349 35037 111383 35071
rect 112545 35037 112579 35071
rect 112913 35037 112947 35071
rect 113189 35037 113223 35071
rect 113557 35037 113591 35071
rect 113649 35037 113683 35071
rect 114017 35037 114051 35071
rect 114109 35037 114143 35071
rect 114293 35037 114327 35071
rect 114477 35037 114511 35071
rect 114753 35037 114787 35071
rect 115213 35037 115247 35071
rect 115305 35037 115339 35071
rect 115489 35037 115523 35071
rect 115673 35037 115707 35071
rect 116225 35037 116259 35071
rect 117421 35037 117455 35071
rect 117697 35037 117731 35071
rect 112269 34969 112303 35003
rect 118157 34969 118191 35003
rect 118341 34969 118375 35003
rect 112453 34901 112487 34935
rect 113373 34901 113407 34935
rect 114569 34901 114603 34935
rect 118065 34901 118099 34935
rect 108589 34697 108623 34731
rect 109233 34697 109267 34731
rect 109417 34697 109451 34731
rect 109693 34697 109727 34731
rect 111986 34697 112020 34731
rect 114109 34697 114143 34731
rect 114385 34697 114419 34731
rect 116041 34697 116075 34731
rect 109969 34629 110003 34663
rect 110705 34629 110739 34663
rect 110965 34629 110999 34663
rect 111165 34629 111199 34663
rect 112269 34629 112303 34663
rect 108497 34561 108531 34595
rect 108681 34561 108715 34595
rect 108865 34561 108899 34595
rect 109049 34561 109083 34595
rect 109325 34561 109359 34595
rect 109509 34561 109543 34595
rect 109601 34561 109635 34595
rect 109877 34561 109911 34595
rect 111809 34561 111843 34595
rect 111901 34561 111935 34595
rect 112085 34561 112119 34595
rect 112361 34561 112395 34595
rect 113741 34561 113775 34595
rect 114201 34565 114235 34599
rect 115029 34561 115063 34595
rect 115673 34561 115707 34595
rect 117237 34561 117271 34595
rect 117513 34561 117547 34595
rect 117697 34561 117731 34595
rect 110337 34493 110371 34527
rect 113833 34493 113867 34527
rect 115121 34493 115155 34527
rect 115305 34493 115339 34527
rect 115581 34493 115615 34527
rect 117329 34493 117363 34527
rect 110540 34425 110574 34459
rect 114661 34425 114695 34459
rect 117421 34425 117455 34459
rect 109877 34357 109911 34391
rect 110429 34357 110463 34391
rect 110797 34357 110831 34391
rect 110981 34357 111015 34391
rect 117053 34357 117087 34391
rect 108865 34153 108899 34187
rect 109969 34153 110003 34187
rect 110429 34153 110463 34187
rect 113557 34153 113591 34187
rect 113741 34153 113775 34187
rect 114017 34153 114051 34187
rect 115581 34153 115615 34187
rect 117237 34153 117271 34187
rect 118157 34153 118191 34187
rect 111441 34085 111475 34119
rect 110153 34017 110187 34051
rect 115857 34017 115891 34051
rect 117329 34017 117363 34051
rect 117697 34017 117731 34051
rect 108497 33949 108531 33983
rect 108681 33949 108715 33983
rect 109049 33949 109083 33983
rect 109509 33949 109543 33983
rect 109969 33949 110003 33983
rect 110245 33949 110279 33983
rect 110981 33949 111015 33983
rect 111165 33949 111199 33983
rect 111625 33949 111659 33983
rect 114017 33949 114051 33983
rect 114293 33949 114327 33983
rect 114937 33949 114971 33983
rect 115121 33949 115155 33983
rect 115397 33949 115431 33983
rect 116041 33949 116075 33983
rect 116133 33949 116167 33983
rect 116593 33949 116627 33983
rect 116777 33949 116811 33983
rect 117053 33949 117087 33983
rect 117513 33949 117547 33983
rect 117973 33949 118007 33983
rect 111993 33881 112027 33915
rect 113725 33881 113759 33915
rect 113925 33881 113959 33915
rect 115029 33881 115063 33915
rect 115213 33881 115247 33915
rect 117789 33881 117823 33915
rect 109233 33813 109267 33847
rect 109325 33813 109359 33847
rect 110981 33813 111015 33847
rect 111717 33813 111751 33847
rect 111809 33813 111843 33847
rect 114201 33813 114235 33847
rect 108589 33609 108623 33643
rect 109785 33609 109819 33643
rect 110705 33609 110739 33643
rect 110889 33609 110923 33643
rect 113005 33609 113039 33643
rect 113833 33609 113867 33643
rect 114201 33609 114235 33643
rect 114845 33609 114879 33643
rect 115397 33609 115431 33643
rect 115581 33609 115615 33643
rect 117697 33609 117731 33643
rect 109601 33541 109635 33575
rect 110981 33541 111015 33575
rect 115825 33541 115859 33575
rect 116041 33541 116075 33575
rect 108313 33473 108347 33507
rect 108773 33473 108807 33507
rect 108957 33473 108991 33507
rect 109141 33473 109175 33507
rect 109877 33473 109911 33507
rect 111073 33473 111107 33507
rect 111349 33473 111383 33507
rect 111441 33473 111475 33507
rect 111533 33473 111567 33507
rect 111993 33473 112027 33507
rect 112637 33473 112671 33507
rect 113741 33473 113775 33507
rect 114661 33473 114695 33507
rect 114845 33473 114879 33507
rect 115456 33473 115490 33507
rect 116409 33473 116443 33507
rect 116593 33473 116627 33507
rect 117329 33473 117363 33507
rect 110705 33405 110739 33439
rect 111165 33405 111199 33439
rect 111625 33405 111659 33439
rect 112085 33405 112119 33439
rect 112545 33405 112579 33439
rect 113649 33405 113683 33439
rect 114937 33405 114971 33439
rect 115029 33405 115063 33439
rect 117145 33405 117179 33439
rect 117237 33405 117271 33439
rect 109601 33337 109635 33371
rect 112361 33337 112395 33371
rect 108497 33269 108531 33303
rect 109233 33269 109267 33303
rect 109417 33269 109451 33303
rect 115673 33269 115707 33303
rect 115857 33269 115891 33303
rect 116593 33269 116627 33303
rect 108773 33065 108807 33099
rect 109049 33065 109083 33099
rect 109693 33065 109727 33099
rect 109877 33065 109911 33099
rect 115213 33065 115247 33099
rect 116409 33065 116443 33099
rect 116685 33065 116719 33099
rect 117605 33065 117639 33099
rect 117697 33065 117731 33099
rect 110245 32929 110279 32963
rect 117053 32929 117087 32963
rect 118157 32929 118191 32963
rect 108313 32861 108347 32895
rect 108589 32861 108623 32895
rect 109233 32861 109267 32895
rect 110337 32861 110371 32895
rect 112729 32861 112763 32895
rect 112913 32861 112947 32895
rect 113189 32861 113223 32895
rect 115397 32861 115431 32895
rect 115673 32861 115707 32895
rect 115857 32861 115891 32895
rect 115949 32861 115983 32895
rect 116133 32861 116167 32895
rect 116225 32861 116259 32895
rect 116501 32861 116535 32895
rect 118065 32861 118099 32895
rect 108405 32793 108439 32827
rect 109509 32793 109543 32827
rect 109725 32793 109759 32827
rect 109969 32725 110003 32759
rect 112913 32725 112947 32759
rect 113281 32725 113315 32759
rect 115581 32725 115615 32759
rect 117145 32725 117179 32759
rect 117237 32725 117271 32759
rect 108513 32521 108547 32555
rect 108681 32521 108715 32555
rect 109325 32521 109359 32555
rect 114293 32521 114327 32555
rect 115673 32521 115707 32555
rect 116593 32521 116627 32555
rect 117329 32521 117363 32555
rect 117697 32521 117731 32555
rect 118157 32521 118191 32555
rect 108313 32453 108347 32487
rect 108957 32385 108991 32419
rect 109601 32385 109635 32419
rect 109969 32385 110003 32419
rect 110981 32385 111015 32419
rect 111165 32385 111199 32419
rect 111625 32385 111659 32419
rect 111901 32385 111935 32419
rect 112177 32385 112211 32419
rect 112729 32385 112763 32419
rect 112913 32385 112947 32419
rect 113281 32385 113315 32419
rect 113374 32385 113408 32419
rect 114296 32385 114330 32419
rect 114845 32385 114879 32419
rect 115305 32385 115339 32419
rect 115581 32385 115615 32419
rect 115765 32385 115799 32419
rect 115949 32385 115983 32419
rect 116133 32385 116167 32419
rect 116501 32385 116535 32419
rect 116777 32385 116811 32419
rect 116869 32385 116903 32419
rect 117012 32385 117046 32419
rect 117145 32385 117179 32419
rect 117237 32385 117271 32419
rect 117513 32385 117547 32419
rect 117789 32385 117823 32419
rect 117882 32385 117916 32419
rect 109049 32317 109083 32351
rect 113649 32317 113683 32351
rect 113833 32317 113867 32351
rect 109785 32249 109819 32283
rect 112637 32249 112671 32283
rect 114477 32249 114511 32283
rect 116041 32249 116075 32283
rect 108497 32181 108531 32215
rect 109509 32181 109543 32215
rect 110061 32181 110095 32215
rect 111349 32181 111383 32215
rect 111809 32181 111843 32215
rect 112085 32181 112119 32215
rect 113925 32181 113959 32215
rect 114937 32181 114971 32215
rect 115489 32181 115523 32215
rect 116317 32181 116351 32215
rect 109509 31977 109543 32011
rect 111533 31977 111567 32011
rect 115397 31977 115431 32011
rect 115489 31977 115523 32011
rect 116317 31977 116351 32011
rect 117329 31977 117363 32011
rect 109233 31909 109267 31943
rect 110981 31909 111015 31943
rect 112729 31909 112763 31943
rect 116593 31909 116627 31943
rect 117881 31909 117915 31943
rect 108957 31841 108991 31875
rect 109877 31841 109911 31875
rect 110889 31841 110923 31875
rect 111625 31841 111659 31875
rect 112361 31841 112395 31875
rect 114385 31841 114419 31875
rect 115949 31841 115983 31875
rect 117513 31841 117547 31875
rect 108313 31773 108347 31807
rect 108497 31773 108531 31807
rect 108865 31773 108899 31807
rect 109785 31773 109819 31807
rect 111352 31773 111386 31807
rect 111809 31773 111843 31807
rect 112177 31773 112211 31807
rect 112545 31773 112579 31807
rect 113005 31773 113039 31807
rect 113281 31773 113315 31807
rect 113833 31773 113867 31807
rect 114109 31773 114143 31807
rect 114845 31773 114879 31807
rect 115121 31773 115155 31807
rect 115213 31773 115247 31807
rect 115489 31773 115523 31807
rect 115673 31773 115707 31807
rect 116041 31773 116075 31807
rect 116777 31773 116811 31807
rect 116869 31773 116903 31807
rect 117053 31773 117087 31807
rect 117605 31773 117639 31807
rect 118065 31773 118099 31807
rect 118249 31773 118283 31807
rect 118525 31773 118559 31807
rect 114201 31705 114235 31739
rect 111349 31637 111383 31671
rect 111809 31637 111843 31671
rect 118341 31637 118375 31671
rect 111165 31433 111199 31467
rect 111993 31433 112027 31467
rect 112453 31433 112487 31467
rect 114477 31433 114511 31467
rect 115489 31433 115523 31467
rect 116593 31433 116627 31467
rect 118065 31433 118099 31467
rect 108865 31365 108899 31399
rect 111317 31365 111351 31399
rect 111533 31365 111567 31399
rect 116961 31365 116995 31399
rect 117329 31365 117363 31399
rect 117605 31365 117639 31399
rect 110613 31297 110647 31331
rect 111901 31297 111935 31331
rect 112085 31297 112119 31331
rect 112269 31297 112303 31331
rect 112453 31297 112487 31331
rect 112729 31297 112763 31331
rect 113097 31297 113131 31331
rect 113465 31297 113499 31331
rect 113649 31297 113683 31331
rect 113833 31297 113867 31331
rect 114109 31297 114143 31331
rect 114385 31297 114419 31331
rect 114937 31297 114971 31331
rect 115397 31297 115431 31331
rect 116225 31297 116259 31331
rect 116409 31297 116443 31331
rect 116501 31297 116535 31331
rect 116685 31297 116719 31331
rect 117421 31297 117455 31331
rect 118249 31297 118283 31331
rect 118525 31297 118559 31331
rect 110429 31229 110463 31263
rect 110521 31229 110555 31263
rect 112545 31229 112579 31263
rect 113005 31229 113039 31263
rect 115029 31229 115063 31263
rect 115121 31229 115155 31263
rect 109049 31161 109083 31195
rect 110981 31161 111015 31195
rect 108773 31093 108807 31127
rect 109233 31093 109267 31127
rect 111349 31093 111383 31127
rect 114569 31093 114603 31127
rect 116317 31093 116351 31127
rect 117789 31093 117823 31127
rect 109509 30889 109543 30923
rect 109785 30889 109819 30923
rect 111441 30889 111475 30923
rect 112545 30889 112579 30923
rect 114293 30889 114327 30923
rect 116041 30889 116075 30923
rect 117145 30889 117179 30923
rect 117329 30889 117363 30923
rect 110061 30821 110095 30855
rect 112269 30821 112303 30855
rect 117237 30821 117271 30855
rect 109325 30753 109359 30787
rect 111533 30753 111567 30787
rect 114017 30753 114051 30787
rect 114753 30753 114787 30787
rect 116133 30753 116167 30787
rect 118065 30753 118099 30787
rect 109233 30685 109267 30719
rect 109693 30685 109727 30719
rect 110245 30685 110279 30719
rect 110429 30685 110463 30719
rect 111625 30685 111659 30719
rect 111993 30685 112027 30719
rect 112453 30685 112487 30719
rect 112913 30685 112947 30719
rect 113097 30685 113131 30719
rect 113189 30685 113223 30719
rect 113925 30685 113959 30719
rect 114385 30685 114419 30719
rect 114569 30685 114603 30719
rect 114661 30685 114695 30719
rect 114845 30685 114879 30719
rect 115857 30685 115891 30719
rect 116317 30685 116351 30719
rect 116593 30685 116627 30719
rect 116777 30685 116811 30719
rect 116869 30685 116903 30719
rect 117973 30685 118007 30719
rect 118249 30685 118283 30719
rect 111901 30617 111935 30651
rect 112269 30617 112303 30651
rect 113281 30617 113315 30651
rect 113465 30617 113499 30651
rect 114477 30617 114511 30651
rect 116685 30617 116719 30651
rect 111809 30549 111843 30583
rect 112085 30549 112119 30583
rect 113649 30549 113683 30583
rect 116501 30549 116535 30583
rect 116961 30549 116995 30583
rect 117605 30549 117639 30583
rect 117789 30549 117823 30583
rect 109233 30345 109267 30379
rect 112085 30345 112119 30379
rect 113649 30345 113683 30379
rect 111165 30277 111199 30311
rect 111901 30277 111935 30311
rect 113281 30277 113315 30311
rect 113925 30277 113959 30311
rect 114036 30277 114070 30311
rect 115489 30277 115523 30311
rect 115705 30277 115739 30311
rect 116869 30277 116903 30311
rect 118525 30277 118559 30311
rect 109785 30209 109819 30243
rect 109969 30209 110003 30243
rect 110061 30209 110095 30243
rect 110153 30209 110187 30243
rect 110521 30209 110555 30243
rect 110613 30209 110647 30243
rect 110797 30209 110831 30243
rect 110889 30209 110923 30243
rect 111349 30209 111383 30243
rect 111441 30209 111475 30243
rect 111717 30209 111751 30243
rect 111993 30209 112027 30243
rect 112085 30209 112119 30243
rect 112269 30209 112303 30243
rect 113465 30209 113499 30243
rect 113741 30209 113775 30243
rect 113833 30209 113867 30243
rect 115121 30209 115155 30243
rect 115213 30209 115247 30243
rect 115397 30209 115431 30243
rect 116225 30209 116259 30243
rect 116501 30209 116535 30243
rect 116731 30209 116765 30243
rect 116961 30209 116995 30243
rect 117144 30209 117178 30243
rect 117237 30209 117271 30243
rect 117697 30209 117731 30243
rect 117881 30209 117915 30243
rect 117973 30209 118007 30243
rect 118249 30209 118283 30243
rect 109693 30141 109727 30175
rect 110429 30141 110463 30175
rect 111073 30141 111107 30175
rect 114201 30141 114235 30175
rect 109417 30073 109451 30107
rect 111993 30073 112027 30107
rect 114109 30073 114143 30107
rect 115949 30073 115983 30107
rect 118157 30073 118191 30107
rect 111165 30005 111199 30039
rect 115397 30005 115431 30039
rect 115673 30005 115707 30039
rect 115857 30005 115891 30039
rect 116133 30005 116167 30039
rect 116593 30005 116627 30039
rect 117513 30005 117547 30039
rect 109325 29801 109359 29835
rect 110245 29801 110279 29835
rect 115305 29801 115339 29835
rect 115673 29801 115707 29835
rect 117789 29801 117823 29835
rect 118157 29801 118191 29835
rect 111257 29733 111291 29767
rect 113005 29733 113039 29767
rect 112361 29665 112395 29699
rect 113281 29665 113315 29699
rect 115581 29665 115615 29699
rect 109509 29597 109543 29631
rect 109693 29597 109727 29631
rect 109785 29597 109819 29631
rect 109969 29597 110003 29631
rect 110705 29597 110739 29631
rect 110797 29597 110831 29631
rect 110981 29597 111015 29631
rect 111073 29597 111107 29631
rect 111717 29597 111751 29631
rect 111901 29597 111935 29631
rect 113373 29597 113407 29631
rect 114201 29597 114235 29631
rect 114937 29597 114971 29631
rect 115121 29597 115155 29631
rect 115673 29597 115707 29631
rect 115857 29597 115891 29631
rect 116041 29597 116075 29631
rect 116317 29597 116351 29631
rect 116593 29597 116627 29631
rect 117053 29597 117087 29631
rect 117145 29597 117179 29631
rect 118065 29597 118099 29631
rect 118525 29597 118559 29631
rect 110245 29529 110279 29563
rect 112545 29529 112579 29563
rect 114109 29529 114143 29563
rect 116961 29529 116995 29563
rect 117757 29529 117791 29563
rect 117973 29529 118007 29563
rect 110061 29461 110095 29495
rect 111901 29461 111935 29495
rect 112453 29461 112487 29495
rect 112913 29461 112947 29495
rect 114937 29461 114971 29495
rect 116501 29461 116535 29495
rect 116869 29461 116903 29495
rect 117329 29461 117363 29495
rect 117605 29461 117639 29495
rect 118341 29461 118375 29495
rect 109601 29257 109635 29291
rect 109693 29257 109727 29291
rect 110613 29257 110647 29291
rect 117421 29257 117455 29291
rect 110245 29189 110279 29223
rect 110461 29189 110495 29223
rect 115029 29189 115063 29223
rect 115581 29189 115615 29223
rect 117237 29189 117271 29223
rect 117697 29189 117731 29223
rect 109417 29121 109451 29155
rect 109601 29121 109635 29155
rect 109877 29121 109911 29155
rect 110061 29121 110095 29155
rect 110153 29121 110187 29155
rect 111349 29121 111383 29155
rect 113557 29121 113591 29155
rect 113741 29121 113775 29155
rect 113926 29127 113960 29161
rect 114109 29121 114143 29155
rect 114937 29121 114971 29155
rect 115121 29121 115155 29155
rect 115305 29121 115339 29155
rect 115397 29121 115431 29155
rect 115489 29121 115523 29155
rect 115673 29121 115707 29155
rect 115857 29121 115891 29155
rect 115949 29121 115983 29155
rect 116041 29121 116075 29155
rect 116133 29121 116167 29155
rect 116409 29121 116443 29155
rect 116501 29121 116535 29155
rect 116685 29121 116719 29155
rect 116961 29121 116995 29155
rect 117513 29121 117547 29155
rect 111441 29053 111475 29087
rect 113833 29053 113867 29087
rect 110981 28985 111015 29019
rect 113373 28985 113407 29019
rect 114753 28985 114787 29019
rect 117145 28985 117179 29019
rect 117973 28985 118007 29019
rect 118157 28985 118191 29019
rect 118525 28985 118559 29019
rect 110429 28917 110463 28951
rect 116317 28917 116351 28951
rect 116869 28917 116903 28951
rect 117237 28917 117271 28951
rect 110245 28713 110279 28747
rect 111073 28713 111107 28747
rect 111993 28713 112027 28747
rect 113005 28713 113039 28747
rect 114017 28713 114051 28747
rect 115857 28713 115891 28747
rect 118065 28713 118099 28747
rect 112545 28645 112579 28679
rect 113281 28645 113315 28679
rect 110705 28577 110739 28611
rect 114753 28577 114787 28611
rect 114845 28577 114879 28611
rect 117053 28577 117087 28611
rect 109877 28509 109911 28543
rect 109969 28509 110003 28543
rect 110061 28509 110095 28543
rect 110889 28509 110923 28543
rect 112177 28509 112211 28543
rect 112453 28509 112487 28543
rect 112637 28509 112671 28543
rect 113557 28509 113591 28543
rect 114201 28509 114235 28543
rect 114385 28509 114419 28543
rect 114661 28509 114695 28543
rect 114937 28509 114971 28543
rect 115121 28509 115155 28543
rect 115305 28509 115339 28543
rect 116041 28509 116075 28543
rect 116225 28509 116259 28543
rect 117421 28509 117455 28543
rect 117697 28509 117731 28543
rect 117881 28509 117915 28543
rect 118249 28509 118283 28543
rect 118525 28509 118559 28543
rect 112361 28441 112395 28475
rect 113189 28441 113223 28475
rect 113281 28441 113315 28475
rect 113465 28441 113499 28475
rect 117237 28441 117271 28475
rect 112821 28373 112855 28407
rect 112989 28373 113023 28407
rect 114477 28373 114511 28407
rect 115213 28373 115247 28407
rect 117605 28373 117639 28407
rect 117789 28373 117823 28407
rect 118341 28373 118375 28407
rect 109601 28169 109635 28203
rect 113465 28169 113499 28203
rect 114293 28169 114327 28203
rect 117329 28169 117363 28203
rect 118065 28169 118099 28203
rect 118433 28169 118467 28203
rect 113925 28101 113959 28135
rect 115673 28101 115707 28135
rect 109785 28033 109819 28067
rect 109877 28033 109911 28067
rect 109969 28033 110003 28067
rect 110153 28033 110187 28067
rect 111625 28033 111659 28067
rect 111717 28033 111751 28067
rect 112269 28033 112303 28067
rect 112545 28033 112579 28067
rect 112729 28033 112763 28067
rect 113833 28033 113867 28067
rect 114477 28033 114511 28067
rect 114569 28033 114603 28067
rect 114661 28033 114695 28067
rect 114845 28033 114879 28067
rect 115029 28033 115063 28067
rect 115581 28033 115615 28067
rect 115765 28033 115799 28067
rect 116133 28033 116167 28067
rect 116409 28033 116443 28067
rect 116593 28033 116627 28067
rect 116685 28033 116719 28067
rect 116869 28033 116903 28067
rect 117789 28033 117823 28067
rect 118249 28033 118283 28067
rect 111257 27965 111291 27999
rect 114109 27965 114143 27999
rect 116271 27965 116305 27999
rect 117421 27965 117455 27999
rect 117513 27965 117547 27999
rect 117881 27965 117915 27999
rect 116869 27897 116903 27931
rect 111901 27829 111935 27863
rect 112085 27829 112119 27863
rect 115029 27829 115063 27863
rect 116501 27829 116535 27863
rect 116961 27829 116995 27863
rect 110337 27625 110371 27659
rect 114477 27625 114511 27659
rect 116961 27625 116995 27659
rect 118249 27625 118283 27659
rect 111073 27557 111107 27591
rect 113557 27557 113591 27591
rect 116501 27557 116535 27591
rect 117513 27557 117547 27591
rect 118341 27557 118375 27591
rect 109877 27489 109911 27523
rect 111717 27489 111751 27523
rect 113281 27489 113315 27523
rect 114201 27489 114235 27523
rect 115857 27489 115891 27523
rect 116777 27489 116811 27523
rect 117789 27489 117823 27523
rect 109785 27421 109819 27455
rect 110245 27421 110279 27455
rect 110429 27421 110463 27455
rect 110889 27421 110923 27455
rect 111165 27421 111199 27455
rect 111349 27421 111383 27455
rect 111993 27421 112027 27455
rect 112269 27421 112303 27455
rect 113189 27421 113223 27455
rect 114661 27421 114695 27455
rect 114753 27421 114787 27455
rect 114937 27421 114971 27455
rect 115029 27421 115063 27455
rect 115489 27421 115523 27455
rect 116041 27421 116075 27455
rect 116317 27421 116351 27455
rect 116685 27421 116719 27455
rect 116961 27421 116995 27455
rect 117881 27421 117915 27455
rect 118525 27421 118559 27455
rect 110705 27353 110739 27387
rect 111809 27353 111843 27387
rect 112545 27353 112579 27387
rect 112729 27353 112763 27387
rect 114017 27353 114051 27387
rect 116225 27353 116259 27387
rect 110153 27285 110187 27319
rect 111625 27285 111659 27319
rect 112177 27285 112211 27319
rect 112361 27285 112395 27319
rect 113649 27285 113683 27319
rect 114109 27285 114143 27319
rect 115673 27285 115707 27319
rect 110797 27081 110831 27115
rect 113925 27081 113959 27115
rect 115305 27081 115339 27115
rect 115397 27081 115431 27115
rect 118525 27081 118559 27115
rect 115949 27013 115983 27047
rect 116133 27013 116167 27047
rect 110981 26945 111015 26979
rect 111073 26945 111107 26979
rect 111257 26945 111291 26979
rect 111349 26945 111383 26979
rect 112085 26945 112119 26979
rect 113557 26945 113591 26979
rect 114845 26945 114879 26979
rect 115581 26945 115615 26979
rect 115673 26945 115707 26979
rect 115857 26945 115891 26979
rect 112177 26877 112211 26911
rect 113649 26877 113683 26911
rect 114661 26877 114695 26911
rect 114937 26877 114971 26911
rect 111717 26809 111751 26843
rect 115857 26741 115891 26775
rect 111441 26537 111475 26571
rect 114661 26537 114695 26571
rect 115305 26537 115339 26571
rect 115121 26469 115155 26503
rect 111625 26333 111659 26367
rect 111809 26333 111843 26367
rect 114845 26333 114879 26367
rect 115029 26265 115063 26299
rect 115489 26265 115523 26299
rect 115279 26197 115313 26231
rect 115029 25993 115063 26027
rect 114845 25925 114879 25959
rect 115121 25857 115155 25891
rect 114845 25721 114879 25755
rect 7573 17629 7607 17663
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 1593 15929 1627 15963
rect 15945 7497 15979 7531
rect 26985 7497 27019 7531
rect 27905 7497 27939 7531
rect 29561 7497 29595 7531
rect 30205 7497 30239 7531
rect 92857 7497 92891 7531
rect 93041 7497 93075 7531
rect 93225 7497 93259 7531
rect 93409 7497 93443 7531
rect 25881 2601 25915 2635
rect 31677 2601 31711 2635
rect 32965 2601 32999 2635
rect 33793 2601 33827 2635
rect 35081 2601 35115 2635
rect 36185 2601 36219 2635
rect 37473 2601 37507 2635
rect 38301 2601 38335 2635
rect 40049 2601 40083 2635
rect 40877 2601 40911 2635
rect 41981 2601 42015 2635
rect 43269 2601 43303 2635
rect 44557 2601 44591 2635
rect 45845 2601 45879 2635
rect 46673 2601 46707 2635
rect 47777 2601 47811 2635
rect 49065 2601 49099 2635
rect 50353 2601 50387 2635
rect 51641 2601 51675 2635
rect 52469 2601 52503 2635
rect 53573 2601 53607 2635
rect 55045 2601 55079 2635
rect 56149 2601 56183 2635
rect 57437 2601 57471 2635
rect 58265 2601 58299 2635
rect 59553 2601 59587 2635
rect 60841 2601 60875 2635
rect 61945 2601 61979 2635
rect 63233 2601 63267 2635
rect 64061 2601 64095 2635
rect 65349 2601 65383 2635
rect 66637 2601 66671 2635
rect 67741 2601 67775 2635
rect 26065 2397 26099 2431
rect 31861 2397 31895 2431
rect 33149 2397 33183 2431
rect 33609 2397 33643 2431
rect 34897 2397 34931 2431
rect 36369 2397 36403 2431
rect 37657 2397 37691 2431
rect 38117 2397 38151 2431
rect 40233 2397 40267 2431
rect 40693 2397 40727 2431
rect 42165 2397 42199 2431
rect 43453 2397 43487 2431
rect 44741 2397 44775 2431
rect 46029 2397 46063 2431
rect 46489 2397 46523 2431
rect 47961 2397 47995 2431
rect 49249 2397 49283 2431
rect 50537 2397 50571 2431
rect 51825 2397 51859 2431
rect 52285 2397 52319 2431
rect 53757 2397 53791 2431
rect 54861 2397 54895 2431
rect 56333 2397 56367 2431
rect 57621 2397 57655 2431
rect 58081 2397 58115 2431
rect 59369 2397 59403 2431
rect 60657 2397 60691 2431
rect 62129 2397 62163 2431
rect 63417 2397 63451 2431
rect 63877 2397 63911 2431
rect 65165 2397 65199 2431
rect 66453 2397 66487 2431
rect 67925 2397 67959 2431
rect 25789 2261 25823 2295
rect 31585 2261 31619 2295
rect 32873 2261 32907 2295
rect 33517 2261 33551 2295
rect 34805 2261 34839 2295
rect 36093 2261 36127 2295
rect 37381 2261 37415 2295
rect 38025 2261 38059 2295
rect 39957 2261 39991 2295
rect 40601 2261 40635 2295
rect 41889 2261 41923 2295
rect 43177 2261 43211 2295
rect 44465 2261 44499 2295
rect 45753 2261 45787 2295
rect 46397 2261 46431 2295
rect 47685 2261 47719 2295
rect 48973 2261 49007 2295
rect 50261 2261 50295 2295
rect 51549 2261 51583 2295
rect 52193 2261 52227 2295
rect 53481 2261 53515 2295
rect 54769 2261 54803 2295
rect 56057 2261 56091 2295
rect 57345 2261 57379 2295
rect 57989 2261 58023 2295
rect 59277 2261 59311 2295
rect 60565 2261 60599 2295
rect 61853 2261 61887 2295
rect 63141 2261 63175 2295
rect 63785 2261 63819 2295
rect 65073 2261 65107 2295
rect 66361 2261 66395 2295
rect 67649 2261 67683 2295
<< metal1 >>
rect 1104 97402 118864 97424
rect 1104 97350 4214 97402
rect 4266 97350 4278 97402
rect 4330 97350 4342 97402
rect 4394 97350 4406 97402
rect 4458 97350 4470 97402
rect 4522 97350 34934 97402
rect 34986 97350 34998 97402
rect 35050 97350 35062 97402
rect 35114 97350 35126 97402
rect 35178 97350 35190 97402
rect 35242 97350 65654 97402
rect 65706 97350 65718 97402
rect 65770 97350 65782 97402
rect 65834 97350 65846 97402
rect 65898 97350 65910 97402
rect 65962 97350 96374 97402
rect 96426 97350 96438 97402
rect 96490 97350 96502 97402
rect 96554 97350 96566 97402
rect 96618 97350 96630 97402
rect 96682 97350 118864 97402
rect 1104 97328 118864 97350
rect 55585 97291 55643 97297
rect 55585 97257 55597 97291
rect 55631 97288 55643 97291
rect 55766 97288 55772 97300
rect 55631 97260 55772 97288
rect 55631 97257 55643 97260
rect 55585 97251 55643 97257
rect 55766 97248 55772 97260
rect 55824 97248 55830 97300
rect 57698 97248 57704 97300
rect 57756 97288 57762 97300
rect 57977 97291 58035 97297
rect 57977 97288 57989 97291
rect 57756 97260 57989 97288
rect 57756 97248 57762 97260
rect 57977 97257 57989 97260
rect 58023 97257 58035 97291
rect 57977 97251 58035 97257
rect 58802 97248 58808 97300
rect 58860 97248 58866 97300
rect 60090 97248 60096 97300
rect 60148 97248 60154 97300
rect 60642 97248 60648 97300
rect 60700 97288 60706 97300
rect 60737 97291 60795 97297
rect 60737 97288 60749 97291
rect 60700 97260 60749 97288
rect 60700 97248 60706 97260
rect 60737 97257 60749 97260
rect 60783 97257 60795 97291
rect 60737 97251 60795 97257
rect 62666 97248 62672 97300
rect 62724 97248 62730 97300
rect 63310 97248 63316 97300
rect 63368 97248 63374 97300
rect 64598 97248 64604 97300
rect 64656 97248 64662 97300
rect 65242 97248 65248 97300
rect 65300 97248 65306 97300
rect 65334 97248 65340 97300
rect 65392 97288 65398 97300
rect 107838 97288 107844 97300
rect 65392 97260 107844 97288
rect 65392 97248 65398 97260
rect 107838 97248 107844 97260
rect 107896 97248 107902 97300
rect 67174 97180 67180 97232
rect 67232 97180 67238 97232
rect 67818 97180 67824 97232
rect 67876 97180 67882 97232
rect 70302 97180 70308 97232
rect 70360 97220 70366 97232
rect 70489 97223 70547 97229
rect 70489 97220 70501 97223
rect 70360 97192 70501 97220
rect 70360 97180 70366 97192
rect 70489 97189 70501 97192
rect 70535 97189 70547 97223
rect 70489 97183 70547 97189
rect 71682 97180 71688 97232
rect 71740 97180 71746 97232
rect 72326 97180 72332 97232
rect 72384 97180 72390 97232
rect 74350 97180 74356 97232
rect 74408 97180 74414 97232
rect 107470 97180 107476 97232
rect 107528 97180 107534 97232
rect 67634 97112 67640 97164
rect 67692 97152 67698 97164
rect 67692 97124 69980 97152
rect 67692 97112 67698 97124
rect 55769 97087 55827 97093
rect 55769 97053 55781 97087
rect 55815 97084 55827 97087
rect 57422 97084 57428 97096
rect 55815 97056 57428 97084
rect 55815 97053 55827 97056
rect 55769 97047 55827 97053
rect 57422 97044 57428 97056
rect 57480 97044 57486 97096
rect 58158 97044 58164 97096
rect 58216 97044 58222 97096
rect 58989 97087 59047 97093
rect 58989 97053 59001 97087
rect 59035 97084 59047 97087
rect 59262 97084 59268 97096
rect 59035 97056 59268 97084
rect 59035 97053 59047 97056
rect 58989 97047 59047 97053
rect 59262 97044 59268 97056
rect 59320 97044 59326 97096
rect 60277 97087 60335 97093
rect 60277 97053 60289 97087
rect 60323 97084 60335 97087
rect 60550 97084 60556 97096
rect 60323 97056 60556 97084
rect 60323 97053 60335 97056
rect 60277 97047 60335 97053
rect 60550 97044 60556 97056
rect 60608 97044 60614 97096
rect 60918 97044 60924 97096
rect 60976 97044 60982 97096
rect 62850 97044 62856 97096
rect 62908 97044 62914 97096
rect 63494 97044 63500 97096
rect 63552 97044 63558 97096
rect 64785 97087 64843 97093
rect 64785 97053 64797 97087
rect 64831 97084 64843 97087
rect 64966 97084 64972 97096
rect 64831 97056 64972 97084
rect 64831 97053 64843 97056
rect 64785 97047 64843 97053
rect 64966 97044 64972 97056
rect 65024 97044 65030 97096
rect 65429 97087 65487 97093
rect 65429 97053 65441 97087
rect 65475 97084 65487 97087
rect 66714 97084 66720 97096
rect 65475 97056 66720 97084
rect 65475 97053 65487 97056
rect 65429 97047 65487 97053
rect 66714 97044 66720 97056
rect 66772 97044 66778 97096
rect 67358 97044 67364 97096
rect 67416 97044 67422 97096
rect 68002 97044 68008 97096
rect 68060 97044 68066 97096
rect 69952 97093 69980 97124
rect 69937 97087 69995 97093
rect 69937 97053 69949 97087
rect 69983 97053 69995 97087
rect 69937 97047 69995 97053
rect 70026 97044 70032 97096
rect 70084 97084 70090 97096
rect 70305 97087 70363 97093
rect 70305 97084 70317 97087
rect 70084 97056 70317 97084
rect 70084 97044 70090 97056
rect 70305 97053 70317 97056
rect 70351 97053 70363 97087
rect 70305 97047 70363 97053
rect 71866 97044 71872 97096
rect 71924 97044 71930 97096
rect 72510 97044 72516 97096
rect 72568 97044 72574 97096
rect 74166 97044 74172 97096
rect 74224 97044 74230 97096
rect 107488 97084 107516 97180
rect 107657 97087 107715 97093
rect 107657 97084 107669 97087
rect 107488 97056 107669 97084
rect 107657 97053 107669 97056
rect 107703 97053 107715 97087
rect 107657 97047 107715 97053
rect 56594 96976 56600 97028
rect 56652 97016 56658 97028
rect 57609 97019 57667 97025
rect 57609 97016 57621 97019
rect 56652 96988 57621 97016
rect 56652 96976 56658 96988
rect 57609 96985 57621 96988
rect 57655 97016 57667 97019
rect 58253 97019 58311 97025
rect 58253 97016 58265 97019
rect 57655 96988 58265 97016
rect 57655 96985 57667 96988
rect 57609 96979 57667 96985
rect 58253 96985 58265 96988
rect 58299 96985 58311 97019
rect 58253 96979 58311 96985
rect 67450 96976 67456 97028
rect 67508 97016 67514 97028
rect 68189 97019 68247 97025
rect 68189 97016 68201 97019
rect 67508 96988 68201 97016
rect 67508 96976 67514 96988
rect 68189 96985 68201 96988
rect 68235 96985 68247 97019
rect 68189 96979 68247 96985
rect 56137 96951 56195 96957
rect 56137 96917 56149 96951
rect 56183 96948 56195 96951
rect 56226 96948 56232 96960
rect 56183 96920 56232 96948
rect 56183 96917 56195 96920
rect 56137 96911 56195 96917
rect 56226 96908 56232 96920
rect 56284 96908 56290 96960
rect 67634 96908 67640 96960
rect 67692 96908 67698 96960
rect 107838 96908 107844 96960
rect 107896 96948 107902 96960
rect 108025 96951 108083 96957
rect 108025 96948 108037 96951
rect 107896 96920 108037 96948
rect 107896 96908 107902 96920
rect 108025 96917 108037 96920
rect 108071 96917 108083 96951
rect 108025 96911 108083 96917
rect 1104 96858 118864 96880
rect 1104 96806 4874 96858
rect 4926 96806 4938 96858
rect 4990 96806 5002 96858
rect 5054 96806 5066 96858
rect 5118 96806 5130 96858
rect 5182 96806 35594 96858
rect 35646 96806 35658 96858
rect 35710 96806 35722 96858
rect 35774 96806 35786 96858
rect 35838 96806 35850 96858
rect 35902 96806 66314 96858
rect 66366 96806 66378 96858
rect 66430 96806 66442 96858
rect 66494 96806 66506 96858
rect 66558 96806 66570 96858
rect 66622 96806 97034 96858
rect 97086 96806 97098 96858
rect 97150 96806 97162 96858
rect 97214 96806 97226 96858
rect 97278 96806 97290 96858
rect 97342 96806 118864 96858
rect 1104 96784 118864 96806
rect 56226 96636 56232 96688
rect 56284 96676 56290 96688
rect 56778 96676 56784 96688
rect 56284 96648 56784 96676
rect 56284 96636 56290 96648
rect 56778 96636 56784 96648
rect 56836 96636 56842 96688
rect 69290 96568 69296 96620
rect 69348 96568 69354 96620
rect 68830 96432 68836 96484
rect 68888 96472 68894 96484
rect 69109 96475 69167 96481
rect 69109 96472 69121 96475
rect 68888 96444 69121 96472
rect 68888 96432 68894 96444
rect 69109 96441 69121 96444
rect 69155 96441 69167 96475
rect 69109 96435 69167 96441
rect 1104 96314 118864 96336
rect 1104 96262 4214 96314
rect 4266 96262 4278 96314
rect 4330 96262 4342 96314
rect 4394 96262 4406 96314
rect 4458 96262 4470 96314
rect 4522 96262 34934 96314
rect 34986 96262 34998 96314
rect 35050 96262 35062 96314
rect 35114 96262 35126 96314
rect 35178 96262 35190 96314
rect 35242 96262 65654 96314
rect 65706 96262 65718 96314
rect 65770 96262 65782 96314
rect 65834 96262 65846 96314
rect 65898 96262 65910 96314
rect 65962 96262 96374 96314
rect 96426 96262 96438 96314
rect 96490 96262 96502 96314
rect 96554 96262 96566 96314
rect 96618 96262 96630 96314
rect 96682 96262 118864 96314
rect 1104 96240 118864 96262
rect 58158 96160 58164 96212
rect 58216 96200 58222 96212
rect 58529 96203 58587 96209
rect 58529 96200 58541 96203
rect 58216 96172 58541 96200
rect 58216 96160 58222 96172
rect 58529 96169 58541 96172
rect 58575 96169 58587 96203
rect 58529 96163 58587 96169
rect 67821 96203 67879 96209
rect 67821 96169 67833 96203
rect 67867 96200 67879 96203
rect 68002 96200 68008 96212
rect 67867 96172 68008 96200
rect 67867 96169 67879 96172
rect 67821 96163 67879 96169
rect 68002 96160 68008 96172
rect 68060 96160 68066 96212
rect 73433 96203 73491 96209
rect 73433 96169 73445 96203
rect 73479 96200 73491 96203
rect 74166 96200 74172 96212
rect 73479 96172 74172 96200
rect 73479 96169 73491 96172
rect 73433 96163 73491 96169
rect 74166 96160 74172 96172
rect 74224 96160 74230 96212
rect 67450 96092 67456 96144
rect 67508 96092 67514 96144
rect 56778 96024 56784 96076
rect 56836 96024 56842 96076
rect 66073 96067 66131 96073
rect 66073 96033 66085 96067
rect 66119 96064 66131 96067
rect 67468 96064 67496 96092
rect 66119 96036 67496 96064
rect 66119 96033 66131 96036
rect 66073 96027 66131 96033
rect 70762 95956 70768 96008
rect 70820 95996 70826 96008
rect 71685 95999 71743 96005
rect 71685 95996 71697 95999
rect 70820 95968 71697 95996
rect 70820 95956 70826 95968
rect 71685 95965 71697 95968
rect 71731 95965 71743 95999
rect 71685 95959 71743 95965
rect 57054 95888 57060 95940
rect 57112 95888 57118 95940
rect 59170 95928 59176 95940
rect 58282 95900 59176 95928
rect 59170 95888 59176 95900
rect 59228 95888 59234 95940
rect 66349 95931 66407 95937
rect 66349 95897 66361 95931
rect 66395 95897 66407 95931
rect 69106 95928 69112 95940
rect 67574 95900 69112 95928
rect 66349 95891 66407 95897
rect 66364 95860 66392 95891
rect 69106 95888 69112 95900
rect 69164 95888 69170 95940
rect 71958 95888 71964 95940
rect 72016 95888 72022 95940
rect 74718 95928 74724 95940
rect 73186 95900 74724 95928
rect 74718 95888 74724 95900
rect 74776 95888 74782 95940
rect 66990 95860 66996 95872
rect 66364 95832 66996 95860
rect 66990 95820 66996 95832
rect 67048 95820 67054 95872
rect 1104 95770 118864 95792
rect 1104 95718 4874 95770
rect 4926 95718 4938 95770
rect 4990 95718 5002 95770
rect 5054 95718 5066 95770
rect 5118 95718 5130 95770
rect 5182 95718 35594 95770
rect 35646 95718 35658 95770
rect 35710 95718 35722 95770
rect 35774 95718 35786 95770
rect 35838 95718 35850 95770
rect 35902 95718 66314 95770
rect 66366 95718 66378 95770
rect 66430 95718 66442 95770
rect 66494 95718 66506 95770
rect 66558 95718 66570 95770
rect 66622 95718 97034 95770
rect 97086 95718 97098 95770
rect 97150 95718 97162 95770
rect 97214 95718 97226 95770
rect 97278 95718 97290 95770
rect 97342 95718 118864 95770
rect 1104 95696 118864 95718
rect 57422 95616 57428 95668
rect 57480 95616 57486 95668
rect 60918 95616 60924 95668
rect 60976 95656 60982 95668
rect 61013 95659 61071 95665
rect 61013 95656 61025 95659
rect 60976 95628 61025 95656
rect 60976 95616 60982 95628
rect 61013 95625 61025 95628
rect 61059 95625 61071 95659
rect 62758 95656 62764 95668
rect 61013 95619 61071 95625
rect 61764 95628 62764 95656
rect 54478 95548 54484 95600
rect 54536 95588 54542 95600
rect 55953 95591 56011 95597
rect 55953 95588 55965 95591
rect 54536 95560 55965 95588
rect 54536 95548 54542 95560
rect 55953 95557 55965 95560
rect 55999 95557 56011 95591
rect 57698 95588 57704 95600
rect 57178 95560 57704 95588
rect 55953 95551 56011 95557
rect 57698 95548 57704 95560
rect 57756 95548 57762 95600
rect 59541 95591 59599 95597
rect 59541 95588 59553 95591
rect 57808 95560 59553 95588
rect 57606 95480 57612 95532
rect 57664 95520 57670 95532
rect 57808 95520 57836 95560
rect 59541 95557 59553 95560
rect 59587 95557 59599 95591
rect 61764 95588 61792 95628
rect 62758 95616 62764 95628
rect 62816 95616 62822 95668
rect 62850 95616 62856 95668
rect 62908 95616 62914 95668
rect 64874 95656 64880 95668
rect 63880 95628 64880 95656
rect 63880 95588 63908 95628
rect 64874 95616 64880 95628
rect 64932 95616 64938 95668
rect 64966 95616 64972 95668
rect 65024 95616 65030 95668
rect 66622 95656 66628 95668
rect 65720 95628 66628 95656
rect 65720 95588 65748 95628
rect 66622 95616 66628 95628
rect 66680 95616 66686 95668
rect 66714 95616 66720 95668
rect 66772 95656 66778 95668
rect 66809 95659 66867 95665
rect 66809 95656 66821 95659
rect 66772 95628 66821 95656
rect 66772 95616 66778 95628
rect 66809 95625 66821 95628
rect 66855 95625 66867 95659
rect 71777 95659 71835 95665
rect 66809 95619 66867 95625
rect 68204 95628 70072 95656
rect 67082 95588 67088 95600
rect 60766 95560 61792 95588
rect 62606 95560 63908 95588
rect 64722 95560 65748 95588
rect 66562 95560 67088 95588
rect 59541 95551 59599 95557
rect 67082 95548 67088 95560
rect 67140 95548 67146 95600
rect 68204 95529 68232 95628
rect 69934 95588 69940 95600
rect 69690 95560 69940 95588
rect 69934 95548 69940 95560
rect 69992 95548 69998 95600
rect 70044 95588 70072 95628
rect 71777 95625 71789 95659
rect 71823 95656 71835 95659
rect 71866 95656 71872 95668
rect 71823 95628 71872 95656
rect 71823 95625 71835 95628
rect 71777 95619 71835 95625
rect 71866 95616 71872 95628
rect 71924 95616 71930 95668
rect 70578 95588 70584 95600
rect 70044 95560 70584 95588
rect 70044 95529 70072 95560
rect 70578 95548 70584 95560
rect 70636 95548 70642 95600
rect 71682 95588 71688 95600
rect 71530 95560 71688 95588
rect 71682 95548 71688 95560
rect 71740 95548 71746 95600
rect 57664 95492 57836 95520
rect 68189 95523 68247 95529
rect 57664 95480 57670 95492
rect 68189 95489 68201 95523
rect 68235 95489 68247 95523
rect 68189 95483 68247 95489
rect 70029 95523 70087 95529
rect 70029 95489 70041 95523
rect 70075 95489 70087 95523
rect 70029 95483 70087 95489
rect 55674 95412 55680 95464
rect 55732 95412 55738 95464
rect 57882 95412 57888 95464
rect 57940 95452 57946 95464
rect 59265 95455 59323 95461
rect 59265 95452 59277 95455
rect 57940 95424 59277 95452
rect 57940 95412 57946 95424
rect 59265 95421 59277 95424
rect 59311 95421 59323 95455
rect 61105 95455 61163 95461
rect 61105 95452 61117 95455
rect 59265 95415 59323 95421
rect 60568 95424 61117 95452
rect 59280 95316 59308 95415
rect 59538 95316 59544 95328
rect 59280 95288 59544 95316
rect 59538 95276 59544 95288
rect 59596 95316 59602 95328
rect 60568 95316 60596 95424
rect 61105 95421 61117 95424
rect 61151 95421 61163 95455
rect 61381 95455 61439 95461
rect 61381 95452 61393 95455
rect 61105 95415 61163 95421
rect 61212 95424 61393 95452
rect 60734 95344 60740 95396
rect 60792 95384 60798 95396
rect 61212 95384 61240 95424
rect 61381 95421 61393 95424
rect 61427 95421 61439 95455
rect 61381 95415 61439 95421
rect 63221 95455 63279 95461
rect 63221 95421 63233 95455
rect 63267 95421 63279 95455
rect 63221 95415 63279 95421
rect 63497 95455 63555 95461
rect 63497 95421 63509 95455
rect 63543 95452 63555 95455
rect 63586 95452 63592 95464
rect 63543 95424 63592 95452
rect 63543 95421 63555 95424
rect 63497 95415 63555 95421
rect 63236 95384 63264 95415
rect 63586 95412 63592 95424
rect 63644 95412 63650 95464
rect 65058 95452 65064 95464
rect 64524 95424 65064 95452
rect 60792 95356 61240 95384
rect 62408 95356 63264 95384
rect 60792 95344 60798 95356
rect 59596 95288 60596 95316
rect 59596 95276 59602 95288
rect 62022 95276 62028 95328
rect 62080 95316 62086 95328
rect 62408 95316 62436 95356
rect 62080 95288 62436 95316
rect 63236 95316 63264 95356
rect 64524 95316 64552 95424
rect 65058 95412 65064 95424
rect 65116 95412 65122 95464
rect 65337 95455 65395 95461
rect 65337 95452 65349 95455
rect 65168 95424 65349 95452
rect 64782 95344 64788 95396
rect 64840 95384 64846 95396
rect 65168 95384 65196 95424
rect 65337 95421 65349 95424
rect 65383 95421 65395 95455
rect 65337 95415 65395 95421
rect 67726 95412 67732 95464
rect 67784 95452 67790 95464
rect 68465 95455 68523 95461
rect 68465 95452 68477 95455
rect 67784 95424 68477 95452
rect 67784 95412 67790 95424
rect 68465 95421 68477 95424
rect 68511 95421 68523 95455
rect 68465 95415 68523 95421
rect 69014 95412 69020 95464
rect 69072 95452 69078 95464
rect 70305 95455 70363 95461
rect 70305 95452 70317 95455
rect 69072 95424 70317 95452
rect 69072 95412 69078 95424
rect 70305 95421 70317 95424
rect 70351 95421 70363 95455
rect 70305 95415 70363 95421
rect 64840 95356 65196 95384
rect 69937 95387 69995 95393
rect 64840 95344 64846 95356
rect 69937 95353 69949 95387
rect 69983 95384 69995 95387
rect 70026 95384 70032 95396
rect 69983 95356 70032 95384
rect 69983 95353 69995 95356
rect 69937 95347 69995 95353
rect 70026 95344 70032 95356
rect 70084 95344 70090 95396
rect 63236 95288 64552 95316
rect 62080 95276 62086 95288
rect 1104 95226 118864 95248
rect 1104 95174 4214 95226
rect 4266 95174 4278 95226
rect 4330 95174 4342 95226
rect 4394 95174 4406 95226
rect 4458 95174 4470 95226
rect 4522 95174 34934 95226
rect 34986 95174 34998 95226
rect 35050 95174 35062 95226
rect 35114 95174 35126 95226
rect 35178 95174 35190 95226
rect 35242 95174 65654 95226
rect 65706 95174 65718 95226
rect 65770 95174 65782 95226
rect 65834 95174 65846 95226
rect 65898 95174 65910 95226
rect 65962 95174 96374 95226
rect 96426 95174 96438 95226
rect 96490 95174 96502 95226
rect 96554 95174 96566 95226
rect 96618 95174 96630 95226
rect 96682 95174 118864 95226
rect 1104 95152 118864 95174
rect 59262 95072 59268 95124
rect 59320 95112 59326 95124
rect 59633 95115 59691 95121
rect 59633 95112 59645 95115
rect 59320 95084 59645 95112
rect 59320 95072 59326 95084
rect 59633 95081 59645 95084
rect 59679 95081 59691 95115
rect 59633 95075 59691 95081
rect 63494 95072 63500 95124
rect 63552 95112 63558 95124
rect 63773 95115 63831 95121
rect 63773 95112 63785 95115
rect 63552 95084 63785 95112
rect 63552 95072 63558 95084
rect 63773 95081 63785 95084
rect 63819 95081 63831 95115
rect 63773 95075 63831 95081
rect 67358 95072 67364 95124
rect 67416 95072 67422 95124
rect 69201 95115 69259 95121
rect 69201 95081 69213 95115
rect 69247 95112 69259 95115
rect 69290 95112 69296 95124
rect 69247 95084 69296 95112
rect 69247 95081 69259 95084
rect 69201 95075 69259 95081
rect 69290 95072 69296 95084
rect 69348 95072 69354 95124
rect 72510 95072 72516 95124
rect 72568 95072 72574 95124
rect 54662 94936 54668 94988
rect 54720 94976 54726 94988
rect 56045 94979 56103 94985
rect 56045 94976 56057 94979
rect 54720 94948 56057 94976
rect 54720 94936 54726 94948
rect 56045 94945 56057 94948
rect 56091 94945 56103 94979
rect 56045 94939 56103 94945
rect 56060 94908 56088 94939
rect 56778 94936 56784 94988
rect 56836 94976 56842 94988
rect 57882 94976 57888 94988
rect 56836 94948 57888 94976
rect 56836 94936 56842 94948
rect 57882 94936 57888 94948
rect 57940 94936 57946 94988
rect 62022 94936 62028 94988
rect 62080 94936 62086 94988
rect 65058 94936 65064 94988
rect 65116 94976 65122 94988
rect 65613 94979 65671 94985
rect 65613 94976 65625 94979
rect 65116 94948 65625 94976
rect 65116 94936 65122 94948
rect 65613 94945 65625 94948
rect 65659 94976 65671 94979
rect 66898 94976 66904 94988
rect 65659 94948 66904 94976
rect 65659 94945 65671 94948
rect 65613 94939 65671 94945
rect 66898 94936 66904 94948
rect 66956 94976 66962 94988
rect 67450 94976 67456 94988
rect 66956 94948 67456 94976
rect 66956 94936 66962 94948
rect 67450 94936 67456 94948
rect 67508 94936 67514 94988
rect 56870 94908 56876 94920
rect 56060 94880 56876 94908
rect 56870 94868 56876 94880
rect 56928 94868 56934 94920
rect 66990 94868 66996 94920
rect 67048 94868 67054 94920
rect 68830 94868 68836 94920
rect 68888 94868 68894 94920
rect 70762 94868 70768 94920
rect 70820 94868 70826 94920
rect 56229 94843 56287 94849
rect 56229 94809 56241 94843
rect 56275 94840 56287 94843
rect 57790 94840 57796 94852
rect 56275 94812 57796 94840
rect 56275 94809 56287 94812
rect 56229 94803 56287 94809
rect 57790 94800 57796 94812
rect 57848 94800 57854 94852
rect 58161 94843 58219 94849
rect 58161 94809 58173 94843
rect 58207 94809 58219 94843
rect 61746 94840 61752 94852
rect 59386 94812 61752 94840
rect 58161 94803 58219 94809
rect 55214 94732 55220 94784
rect 55272 94772 55278 94784
rect 56321 94775 56379 94781
rect 56321 94772 56333 94775
rect 55272 94744 56333 94772
rect 55272 94732 55278 94744
rect 56321 94741 56333 94744
rect 56367 94741 56379 94775
rect 56321 94735 56379 94741
rect 56689 94775 56747 94781
rect 56689 94741 56701 94775
rect 56735 94772 56747 94775
rect 58176 94772 58204 94803
rect 61746 94800 61752 94812
rect 61804 94800 61810 94852
rect 62298 94800 62304 94852
rect 62356 94800 62362 94852
rect 65242 94840 65248 94852
rect 63526 94812 65248 94840
rect 65242 94800 65248 94812
rect 65300 94800 65306 94852
rect 65889 94843 65947 94849
rect 65889 94809 65901 94843
rect 65935 94809 65947 94843
rect 65889 94803 65947 94809
rect 56735 94744 58204 94772
rect 56735 94741 56747 94744
rect 56689 94735 56747 94741
rect 64138 94732 64144 94784
rect 64196 94772 64202 94784
rect 65904 94772 65932 94803
rect 67174 94800 67180 94852
rect 67232 94840 67238 94852
rect 67729 94843 67787 94849
rect 67729 94840 67741 94843
rect 67232 94812 67741 94840
rect 67232 94800 67238 94812
rect 67729 94809 67741 94812
rect 67775 94809 67787 94843
rect 67729 94803 67787 94809
rect 69750 94800 69756 94852
rect 69808 94840 69814 94852
rect 71041 94843 71099 94849
rect 71041 94840 71053 94843
rect 69808 94812 71053 94840
rect 69808 94800 69814 94812
rect 71041 94809 71053 94812
rect 71087 94809 71099 94843
rect 72970 94840 72976 94852
rect 72266 94812 72976 94840
rect 71041 94803 71099 94809
rect 72970 94800 72976 94812
rect 73028 94800 73034 94852
rect 64196 94744 65932 94772
rect 64196 94732 64202 94744
rect 1104 94682 118864 94704
rect 1104 94630 4874 94682
rect 4926 94630 4938 94682
rect 4990 94630 5002 94682
rect 5054 94630 5066 94682
rect 5118 94630 5130 94682
rect 5182 94630 35594 94682
rect 35646 94630 35658 94682
rect 35710 94630 35722 94682
rect 35774 94630 35786 94682
rect 35838 94630 35850 94682
rect 35902 94630 66314 94682
rect 66366 94630 66378 94682
rect 66430 94630 66442 94682
rect 66494 94630 66506 94682
rect 66558 94630 66570 94682
rect 66622 94630 97034 94682
rect 97086 94630 97098 94682
rect 97150 94630 97162 94682
rect 97214 94630 97226 94682
rect 97278 94630 97290 94682
rect 97342 94630 118864 94682
rect 1104 94608 118864 94630
rect 55309 94571 55367 94577
rect 55309 94537 55321 94571
rect 55355 94568 55367 94571
rect 57054 94568 57060 94580
rect 55355 94540 57060 94568
rect 55355 94537 55367 94540
rect 55309 94531 55367 94537
rect 57054 94528 57060 94540
rect 57112 94528 57118 94580
rect 58345 94571 58403 94577
rect 58345 94537 58357 94571
rect 58391 94568 58403 94571
rect 59998 94568 60004 94580
rect 58391 94540 60004 94568
rect 58391 94537 58403 94540
rect 58345 94531 58403 94537
rect 59998 94528 60004 94540
rect 60056 94528 60062 94580
rect 60550 94528 60556 94580
rect 60608 94568 60614 94580
rect 61289 94571 61347 94577
rect 61289 94568 61301 94571
rect 60608 94540 61301 94568
rect 60608 94528 60614 94540
rect 61289 94537 61301 94540
rect 61335 94537 61347 94571
rect 61289 94531 61347 94537
rect 61746 94528 61752 94580
rect 61804 94528 61810 94580
rect 65242 94528 65248 94580
rect 65300 94568 65306 94580
rect 65337 94571 65395 94577
rect 65337 94568 65349 94571
rect 65300 94540 65349 94568
rect 65300 94528 65306 94540
rect 65337 94537 65349 94540
rect 65383 94537 65395 94571
rect 65337 94531 65395 94537
rect 57698 94460 57704 94512
rect 57756 94500 57762 94512
rect 59357 94503 59415 94509
rect 59357 94500 59369 94503
rect 57756 94472 59369 94500
rect 57756 94460 57762 94472
rect 59357 94469 59369 94472
rect 59403 94469 59415 94503
rect 60090 94500 60096 94512
rect 59357 94463 59415 94469
rect 59464 94472 60096 94500
rect 52454 94392 52460 94444
rect 52512 94432 52518 94444
rect 54941 94435 54999 94441
rect 54941 94432 54953 94435
rect 52512 94404 54953 94432
rect 52512 94392 52518 94404
rect 54941 94401 54953 94404
rect 54987 94401 54999 94435
rect 54941 94395 54999 94401
rect 55490 94392 55496 94444
rect 55548 94432 55554 94444
rect 55585 94435 55643 94441
rect 55585 94432 55597 94435
rect 55548 94404 55597 94432
rect 55548 94392 55554 94404
rect 55585 94401 55597 94404
rect 55631 94432 55643 94435
rect 55674 94432 55680 94444
rect 55631 94404 55680 94432
rect 55631 94401 55643 94404
rect 55585 94395 55643 94401
rect 55674 94392 55680 94404
rect 55732 94392 55738 94444
rect 55858 94441 55864 94444
rect 55852 94432 55864 94441
rect 55819 94404 55864 94432
rect 55852 94395 55864 94404
rect 55858 94392 55864 94395
rect 55916 94392 55922 94444
rect 58434 94392 58440 94444
rect 58492 94392 58498 94444
rect 59464 94441 59492 94472
rect 60090 94460 60096 94472
rect 60148 94460 60154 94512
rect 63218 94500 63224 94512
rect 61042 94472 63224 94500
rect 63218 94460 63224 94472
rect 63276 94460 63282 94512
rect 63328 94472 65472 94500
rect 59449 94435 59507 94441
rect 59449 94401 59461 94435
rect 59495 94401 59507 94435
rect 59449 94395 59507 94401
rect 59538 94392 59544 94444
rect 59596 94392 59602 94444
rect 61841 94435 61899 94441
rect 61841 94401 61853 94435
rect 61887 94401 61899 94435
rect 61841 94395 61899 94401
rect 53834 94324 53840 94376
rect 53892 94364 53898 94376
rect 54662 94364 54668 94376
rect 53892 94336 54668 94364
rect 53892 94324 53898 94336
rect 54662 94324 54668 94336
rect 54720 94324 54726 94376
rect 54849 94367 54907 94373
rect 54849 94333 54861 94367
rect 54895 94364 54907 94367
rect 55398 94364 55404 94376
rect 54895 94336 55404 94364
rect 54895 94333 54907 94336
rect 54849 94327 54907 94333
rect 55398 94324 55404 94336
rect 55456 94324 55462 94376
rect 56870 94324 56876 94376
rect 56928 94364 56934 94376
rect 57882 94364 57888 94376
rect 56928 94336 57888 94364
rect 56928 94324 56934 94336
rect 57882 94324 57888 94336
rect 57940 94364 57946 94376
rect 58161 94367 58219 94373
rect 58161 94364 58173 94367
rect 57940 94336 58173 94364
rect 57940 94324 57946 94336
rect 58161 94333 58173 94336
rect 58207 94333 58219 94367
rect 59817 94367 59875 94373
rect 59817 94364 59829 94367
rect 58161 94327 58219 94333
rect 58820 94336 59829 94364
rect 58820 94305 58848 94336
rect 59817 94333 59829 94336
rect 59863 94333 59875 94367
rect 59817 94327 59875 94333
rect 60182 94324 60188 94376
rect 60240 94364 60246 94376
rect 61856 94364 61884 94395
rect 63328 94376 63356 94472
rect 65444 94444 65472 94472
rect 64141 94435 64199 94441
rect 64141 94401 64153 94435
rect 64187 94432 64199 94435
rect 64187 94404 64460 94432
rect 64187 94401 64199 94404
rect 64141 94395 64199 94401
rect 63310 94364 63316 94376
rect 60240 94336 63316 94364
rect 60240 94324 60246 94336
rect 63310 94324 63316 94336
rect 63368 94324 63374 94376
rect 58805 94299 58863 94305
rect 58805 94265 58817 94299
rect 58851 94265 58863 94299
rect 63770 94296 63776 94308
rect 58805 94259 58863 94265
rect 63512 94268 63776 94296
rect 55493 94231 55551 94237
rect 55493 94197 55505 94231
rect 55539 94228 55551 94231
rect 55582 94228 55588 94240
rect 55539 94200 55588 94228
rect 55539 94197 55551 94200
rect 55493 94191 55551 94197
rect 55582 94188 55588 94200
rect 55640 94228 55646 94240
rect 55858 94228 55864 94240
rect 55640 94200 55864 94228
rect 55640 94188 55646 94200
rect 55858 94188 55864 94200
rect 55916 94188 55922 94240
rect 56965 94231 57023 94237
rect 56965 94197 56977 94231
rect 57011 94228 57023 94231
rect 63512 94228 63540 94268
rect 63770 94256 63776 94268
rect 63828 94256 63834 94308
rect 64432 94305 64460 94404
rect 65426 94392 65432 94444
rect 65484 94392 65490 94444
rect 64417 94299 64475 94305
rect 64417 94265 64429 94299
rect 64463 94296 64475 94299
rect 70486 94296 70492 94308
rect 64463 94268 70492 94296
rect 64463 94265 64475 94268
rect 64417 94259 64475 94265
rect 70486 94256 70492 94268
rect 70544 94256 70550 94308
rect 57011 94200 63540 94228
rect 57011 94197 57023 94200
rect 56965 94191 57023 94197
rect 63586 94188 63592 94240
rect 63644 94228 63650 94240
rect 63865 94231 63923 94237
rect 63865 94228 63877 94231
rect 63644 94200 63877 94228
rect 63644 94188 63650 94200
rect 63865 94197 63877 94200
rect 63911 94197 63923 94231
rect 63865 94191 63923 94197
rect 1104 94138 118864 94160
rect 1104 94086 4214 94138
rect 4266 94086 4278 94138
rect 4330 94086 4342 94138
rect 4394 94086 4406 94138
rect 4458 94086 4470 94138
rect 4522 94086 34934 94138
rect 34986 94086 34998 94138
rect 35050 94086 35062 94138
rect 35114 94086 35126 94138
rect 35178 94086 35190 94138
rect 35242 94086 65654 94138
rect 65706 94086 65718 94138
rect 65770 94086 65782 94138
rect 65834 94086 65846 94138
rect 65898 94086 65910 94138
rect 65962 94086 96374 94138
rect 96426 94086 96438 94138
rect 96490 94086 96502 94138
rect 96554 94086 96566 94138
rect 96618 94086 96630 94138
rect 96682 94086 118864 94138
rect 1104 94064 118864 94086
rect 57790 93984 57796 94036
rect 57848 93984 57854 94036
rect 57882 93984 57888 94036
rect 57940 94024 57946 94036
rect 60001 94027 60059 94033
rect 57940 93996 59492 94024
rect 57940 93984 57946 93996
rect 55582 93916 55588 93968
rect 55640 93916 55646 93968
rect 59464 93897 59492 93996
rect 60001 93993 60013 94027
rect 60047 94024 60059 94027
rect 60734 94024 60740 94036
rect 60047 93996 60740 94024
rect 60047 93993 60059 93996
rect 60001 93987 60059 93993
rect 60734 93984 60740 93996
rect 60792 93984 60798 94036
rect 64138 93984 64144 94036
rect 64196 93984 64202 94036
rect 66349 94027 66407 94033
rect 66349 93993 66361 94027
rect 66395 94024 66407 94027
rect 67174 94024 67180 94036
rect 66395 93996 67180 94024
rect 66395 93993 66407 93996
rect 66349 93987 66407 93993
rect 67174 93984 67180 93996
rect 67232 93984 67238 94036
rect 68830 93984 68836 94036
rect 68888 94024 68894 94036
rect 69937 94027 69995 94033
rect 69937 94024 69949 94027
rect 68888 93996 69949 94024
rect 68888 93984 68894 93996
rect 69937 93993 69949 93996
rect 69983 93993 69995 94027
rect 69937 93987 69995 93993
rect 65426 93916 65432 93968
rect 65484 93956 65490 93968
rect 65484 93928 66300 93956
rect 65484 93916 65490 93928
rect 59449 93891 59507 93897
rect 59449 93857 59461 93891
rect 59495 93888 59507 93891
rect 60553 93891 60611 93897
rect 60553 93888 60565 93891
rect 59495 93860 60565 93888
rect 59495 93857 59507 93860
rect 59449 93851 59507 93857
rect 60553 93857 60565 93860
rect 60599 93888 60611 93891
rect 61565 93891 61623 93897
rect 61565 93888 61577 93891
rect 60599 93860 61577 93888
rect 60599 93857 60611 93860
rect 60553 93851 60611 93857
rect 61565 93857 61577 93860
rect 61611 93888 61623 93891
rect 62393 93891 62451 93897
rect 62393 93888 62405 93891
rect 61611 93860 62405 93888
rect 61611 93857 61623 93860
rect 61565 93851 61623 93857
rect 62393 93857 62405 93860
rect 62439 93888 62451 93891
rect 63586 93888 63592 93900
rect 62439 93860 63592 93888
rect 62439 93857 62451 93860
rect 62393 93851 62451 93857
rect 63586 93848 63592 93860
rect 63644 93848 63650 93900
rect 64509 93891 64567 93897
rect 64509 93857 64521 93891
rect 64555 93888 64567 93891
rect 65705 93891 65763 93897
rect 65705 93888 65717 93891
rect 64555 93860 65717 93888
rect 64555 93857 64567 93860
rect 64509 93851 64567 93857
rect 65705 93857 65717 93860
rect 65751 93888 65763 93891
rect 66162 93888 66168 93900
rect 65751 93860 66168 93888
rect 65751 93857 65763 93860
rect 65705 93851 65763 93857
rect 66162 93848 66168 93860
rect 66220 93848 66226 93900
rect 55490 93780 55496 93832
rect 55548 93820 55554 93832
rect 56502 93820 56508 93832
rect 55548 93792 56508 93820
rect 55548 93780 55554 93792
rect 56502 93780 56508 93792
rect 56560 93820 56566 93832
rect 57149 93823 57207 93829
rect 57149 93820 57161 93823
rect 56560 93792 57161 93820
rect 56560 93780 56566 93792
rect 57149 93789 57161 93792
rect 57195 93789 57207 93823
rect 57149 93783 57207 93789
rect 59173 93823 59231 93829
rect 59173 93789 59185 93823
rect 59219 93820 59231 93823
rect 59538 93820 59544 93832
rect 59219 93792 59544 93820
rect 59219 93789 59231 93792
rect 59173 93783 59231 93789
rect 59538 93780 59544 93792
rect 59596 93780 59602 93832
rect 59630 93780 59636 93832
rect 59688 93780 59694 93832
rect 60090 93780 60096 93832
rect 60148 93820 60154 93832
rect 60277 93823 60335 93829
rect 60277 93820 60289 93823
rect 60148 93792 60289 93820
rect 60148 93780 60154 93792
rect 60277 93789 60289 93792
rect 60323 93789 60335 93823
rect 60277 93783 60335 93789
rect 60737 93823 60795 93829
rect 60737 93789 60749 93823
rect 60783 93820 60795 93823
rect 61470 93820 61476 93832
rect 60783 93792 61476 93820
rect 60783 93789 60795 93792
rect 60737 93783 60795 93789
rect 61470 93780 61476 93792
rect 61528 93780 61534 93832
rect 61654 93780 61660 93832
rect 61712 93820 61718 93832
rect 62577 93823 62635 93829
rect 62577 93820 62589 93823
rect 61712 93792 62589 93820
rect 61712 93780 61718 93792
rect 62577 93789 62589 93792
rect 62623 93789 62635 93823
rect 62577 93783 62635 93789
rect 62758 93780 62764 93832
rect 62816 93820 62822 93832
rect 63129 93823 63187 93829
rect 63129 93820 63141 93823
rect 62816 93792 63141 93820
rect 62816 93780 62822 93792
rect 63129 93789 63141 93792
rect 63175 93789 63187 93823
rect 63129 93783 63187 93789
rect 63221 93823 63279 93829
rect 63221 93789 63233 93823
rect 63267 93820 63279 93823
rect 63310 93820 63316 93832
rect 63267 93792 63316 93820
rect 63267 93789 63279 93792
rect 63221 93783 63279 93789
rect 63310 93780 63316 93792
rect 63368 93780 63374 93832
rect 63770 93780 63776 93832
rect 63828 93780 63834 93832
rect 64601 93823 64659 93829
rect 64601 93789 64613 93823
rect 64647 93820 64659 93823
rect 64690 93820 64696 93832
rect 64647 93792 64696 93820
rect 64647 93789 64659 93792
rect 64601 93783 64659 93789
rect 64690 93780 64696 93792
rect 64748 93780 64754 93832
rect 64874 93780 64880 93832
rect 64932 93820 64938 93832
rect 65245 93823 65303 93829
rect 65245 93820 65257 93823
rect 64932 93792 65257 93820
rect 64932 93780 64938 93792
rect 65245 93789 65257 93792
rect 65291 93789 65303 93823
rect 65245 93783 65303 93789
rect 65337 93823 65395 93829
rect 65337 93789 65349 93823
rect 65383 93820 65395 93823
rect 65426 93820 65432 93832
rect 65383 93792 65432 93820
rect 65383 93789 65395 93792
rect 65337 93783 65395 93789
rect 65426 93780 65432 93792
rect 65484 93780 65490 93832
rect 65886 93780 65892 93832
rect 65944 93780 65950 93832
rect 66272 93820 66300 93928
rect 66640 93860 67220 93888
rect 66640 93829 66668 93860
rect 66625 93823 66683 93829
rect 66625 93820 66637 93823
rect 66272 93792 66637 93820
rect 66625 93789 66637 93792
rect 66671 93789 66683 93823
rect 66625 93783 66683 93789
rect 67082 93780 67088 93832
rect 67140 93780 67146 93832
rect 67192 93829 67220 93860
rect 68572 93860 68784 93888
rect 67177 93823 67235 93829
rect 67177 93789 67189 93823
rect 67223 93820 67235 93823
rect 68373 93823 68431 93829
rect 68373 93820 68385 93823
rect 67223 93792 68385 93820
rect 67223 93789 67235 93792
rect 67177 93783 67235 93789
rect 68373 93789 68385 93792
rect 68419 93820 68431 93823
rect 68572 93820 68600 93860
rect 68756 93829 68784 93860
rect 70044 93860 70992 93888
rect 68419 93792 68600 93820
rect 68649 93823 68707 93829
rect 68419 93789 68431 93792
rect 68373 93783 68431 93789
rect 68649 93789 68661 93823
rect 68695 93789 68707 93823
rect 68649 93783 68707 93789
rect 68741 93823 68799 93829
rect 68741 93789 68753 93823
rect 68787 93789 68799 93823
rect 68741 93783 68799 93789
rect 53374 93644 53380 93696
rect 53432 93684 53438 93696
rect 54665 93687 54723 93693
rect 54665 93684 54677 93687
rect 53432 93656 54677 93684
rect 53432 93644 53438 93656
rect 54665 93653 54677 93656
rect 54711 93684 54723 93687
rect 55508 93684 55536 93780
rect 56904 93755 56962 93761
rect 56904 93721 56916 93755
rect 56950 93752 56962 93755
rect 58158 93752 58164 93764
rect 56950 93724 58164 93752
rect 56950 93721 56962 93724
rect 56904 93715 56962 93721
rect 58158 93712 58164 93724
rect 58216 93712 58222 93764
rect 58928 93755 58986 93761
rect 58928 93721 58940 93755
rect 58974 93752 58986 93755
rect 58974 93724 59216 93752
rect 58974 93721 58986 93724
rect 58928 93715 58986 93721
rect 54711 93656 55536 93684
rect 54711 93653 54723 93656
rect 54665 93647 54723 93653
rect 55766 93644 55772 93696
rect 55824 93644 55830 93696
rect 59188 93684 59216 93724
rect 59262 93712 59268 93764
rect 59320 93752 59326 93764
rect 60185 93755 60243 93761
rect 60185 93752 60197 93755
rect 59320 93724 60197 93752
rect 59320 93712 59326 93724
rect 60185 93721 60197 93724
rect 60231 93721 60243 93755
rect 60185 93715 60243 93721
rect 60366 93712 60372 93764
rect 60424 93752 60430 93764
rect 60829 93755 60887 93761
rect 60829 93752 60841 93755
rect 60424 93724 60841 93752
rect 60424 93712 60430 93724
rect 60829 93721 60841 93724
rect 60875 93721 60887 93755
rect 62298 93752 62304 93764
rect 60829 93715 60887 93721
rect 61212 93724 62304 93752
rect 59354 93684 59360 93696
rect 59188 93656 59360 93684
rect 59354 93644 59360 93656
rect 59412 93644 59418 93696
rect 59541 93687 59599 93693
rect 59541 93653 59553 93687
rect 59587 93684 59599 93687
rect 60642 93684 60648 93696
rect 59587 93656 60648 93684
rect 59587 93653 59599 93656
rect 59541 93647 59599 93653
rect 60642 93644 60648 93656
rect 60700 93644 60706 93696
rect 61212 93693 61240 93724
rect 62298 93712 62304 93724
rect 62356 93712 62362 93764
rect 63494 93752 63500 93764
rect 62408 93724 63500 93752
rect 61197 93687 61255 93693
rect 61197 93653 61209 93687
rect 61243 93653 61255 93687
rect 61197 93647 61255 93653
rect 61378 93644 61384 93696
rect 61436 93684 61442 93696
rect 61657 93687 61715 93693
rect 61657 93684 61669 93687
rect 61436 93656 61669 93684
rect 61436 93644 61442 93656
rect 61657 93653 61669 93656
rect 61703 93653 61715 93687
rect 61657 93647 61715 93653
rect 61746 93644 61752 93696
rect 61804 93644 61810 93696
rect 62117 93687 62175 93693
rect 62117 93653 62129 93687
rect 62163 93684 62175 93687
rect 62408 93684 62436 93724
rect 63494 93712 63500 93724
rect 63552 93712 63558 93764
rect 64782 93752 64788 93764
rect 63604 93724 64788 93752
rect 62163 93656 62436 93684
rect 62485 93687 62543 93693
rect 62163 93653 62175 93656
rect 62117 93647 62175 93653
rect 62485 93653 62497 93687
rect 62531 93684 62543 93687
rect 62850 93684 62856 93696
rect 62531 93656 62856 93684
rect 62531 93653 62543 93656
rect 62485 93647 62543 93653
rect 62850 93644 62856 93656
rect 62908 93644 62914 93696
rect 62945 93687 63003 93693
rect 62945 93653 62957 93687
rect 62991 93684 63003 93687
rect 63604 93684 63632 93724
rect 64782 93712 64788 93724
rect 64840 93712 64846 93764
rect 66806 93752 66812 93764
rect 65076 93724 66812 93752
rect 62991 93656 63632 93684
rect 63681 93687 63739 93693
rect 62991 93653 63003 93656
rect 62945 93647 63003 93653
rect 63681 93653 63693 93687
rect 63727 93684 63739 93687
rect 64506 93684 64512 93696
rect 63727 93656 64512 93684
rect 63727 93653 63739 93656
rect 63681 93647 63739 93653
rect 64506 93644 64512 93656
rect 64564 93644 64570 93696
rect 64598 93644 64604 93696
rect 64656 93684 64662 93696
rect 65076 93693 65104 93724
rect 66806 93712 66812 93724
rect 66864 93712 66870 93764
rect 67266 93712 67272 93764
rect 67324 93752 67330 93764
rect 68278 93752 68284 93764
rect 67324 93724 68284 93752
rect 67324 93712 67330 93724
rect 68278 93712 68284 93724
rect 68336 93712 68342 93764
rect 68664 93752 68692 93783
rect 69106 93780 69112 93832
rect 69164 93780 69170 93832
rect 70044 93829 70072 93860
rect 70964 93829 70992 93860
rect 69201 93823 69259 93829
rect 69201 93789 69213 93823
rect 69247 93820 69259 93823
rect 70029 93823 70087 93829
rect 70029 93820 70041 93823
rect 69247 93792 70041 93820
rect 69247 93789 69259 93792
rect 69201 93783 69259 93789
rect 70029 93789 70041 93792
rect 70075 93789 70087 93823
rect 70029 93783 70087 93789
rect 70949 93823 71007 93829
rect 70949 93789 70961 93823
rect 70995 93820 71007 93823
rect 72234 93820 72240 93832
rect 70995 93792 72240 93820
rect 70995 93789 71007 93792
rect 70949 93783 71007 93789
rect 69216 93752 69244 93783
rect 72234 93780 72240 93792
rect 72292 93780 72298 93832
rect 68664 93724 69244 93752
rect 70118 93712 70124 93764
rect 70176 93752 70182 93764
rect 70305 93755 70363 93761
rect 70305 93752 70317 93755
rect 70176 93724 70317 93752
rect 70176 93712 70182 93724
rect 70305 93721 70317 93724
rect 70351 93721 70363 93755
rect 70305 93715 70363 93721
rect 70486 93712 70492 93764
rect 70544 93752 70550 93764
rect 70544 93724 71176 93752
rect 70544 93712 70550 93724
rect 71148 93696 71176 93724
rect 64693 93687 64751 93693
rect 64693 93684 64705 93687
rect 64656 93656 64705 93684
rect 64656 93644 64662 93656
rect 64693 93653 64705 93656
rect 64739 93653 64751 93687
rect 64693 93647 64751 93653
rect 65061 93687 65119 93693
rect 65061 93653 65073 93687
rect 65107 93653 65119 93687
rect 65061 93647 65119 93653
rect 65978 93644 65984 93696
rect 66036 93644 66042 93696
rect 66533 93687 66591 93693
rect 66533 93653 66545 93687
rect 66579 93684 66591 93687
rect 66714 93684 66720 93696
rect 66579 93656 66720 93684
rect 66579 93653 66591 93656
rect 66533 93647 66591 93653
rect 66714 93644 66720 93656
rect 66772 93644 66778 93696
rect 66990 93644 66996 93696
rect 67048 93684 67054 93696
rect 68833 93687 68891 93693
rect 68833 93684 68845 93687
rect 67048 93656 68845 93684
rect 67048 93644 67054 93656
rect 68833 93653 68845 93656
rect 68879 93653 68891 93687
rect 68833 93647 68891 93653
rect 70854 93644 70860 93696
rect 70912 93644 70918 93696
rect 71130 93644 71136 93696
rect 71188 93644 71194 93696
rect 72142 93644 72148 93696
rect 72200 93684 72206 93696
rect 72237 93687 72295 93693
rect 72237 93684 72249 93687
rect 72200 93656 72249 93684
rect 72200 93644 72206 93656
rect 72237 93653 72249 93656
rect 72283 93653 72295 93687
rect 72237 93647 72295 93653
rect 1104 93594 118864 93616
rect 1104 93542 4874 93594
rect 4926 93542 4938 93594
rect 4990 93542 5002 93594
rect 5054 93542 5066 93594
rect 5118 93542 5130 93594
rect 5182 93542 35594 93594
rect 35646 93542 35658 93594
rect 35710 93542 35722 93594
rect 35774 93542 35786 93594
rect 35838 93542 35850 93594
rect 35902 93542 66314 93594
rect 66366 93542 66378 93594
rect 66430 93542 66442 93594
rect 66494 93542 66506 93594
rect 66558 93542 66570 93594
rect 66622 93542 97034 93594
rect 97086 93542 97098 93594
rect 97150 93542 97162 93594
rect 97214 93542 97226 93594
rect 97278 93542 97290 93594
rect 97342 93542 118864 93594
rect 1104 93520 118864 93542
rect 54478 93440 54484 93492
rect 54536 93440 54542 93492
rect 57606 93440 57612 93492
rect 57664 93480 57670 93492
rect 57701 93483 57759 93489
rect 57701 93480 57713 93483
rect 57664 93452 57713 93480
rect 57664 93440 57670 93452
rect 57701 93449 57713 93452
rect 57747 93449 57759 93483
rect 59630 93480 59636 93492
rect 57701 93443 57759 93449
rect 57808 93452 59636 93480
rect 54021 93415 54079 93421
rect 54021 93381 54033 93415
rect 54067 93412 54079 93415
rect 55766 93412 55772 93424
rect 54067 93384 55772 93412
rect 54067 93381 54079 93384
rect 54021 93375 54079 93381
rect 55766 93372 55772 93384
rect 55824 93372 55830 93424
rect 56226 93372 56232 93424
rect 56284 93412 56290 93424
rect 57808 93412 57836 93452
rect 59630 93440 59636 93452
rect 59688 93440 59694 93492
rect 59998 93440 60004 93492
rect 60056 93440 60062 93492
rect 60642 93440 60648 93492
rect 60700 93480 60706 93492
rect 61473 93483 61531 93489
rect 61473 93480 61485 93483
rect 60700 93452 61485 93480
rect 60700 93440 60706 93452
rect 61473 93449 61485 93452
rect 61519 93449 61531 93483
rect 61473 93443 61531 93449
rect 61562 93440 61568 93492
rect 61620 93480 61626 93492
rect 63405 93483 63463 93489
rect 63405 93480 63417 93483
rect 61620 93452 63417 93480
rect 61620 93440 61626 93452
rect 63405 93449 63417 93452
rect 63451 93449 63463 93483
rect 63405 93443 63463 93449
rect 63494 93440 63500 93492
rect 63552 93480 63558 93492
rect 65978 93480 65984 93492
rect 63552 93452 65984 93480
rect 63552 93440 63558 93452
rect 65978 93440 65984 93452
rect 66036 93440 66042 93492
rect 66625 93483 66683 93489
rect 66625 93449 66637 93483
rect 66671 93480 66683 93483
rect 69842 93480 69848 93492
rect 66671 93452 69848 93480
rect 66671 93449 66683 93452
rect 66625 93443 66683 93449
rect 69842 93440 69848 93452
rect 69900 93440 69906 93492
rect 69934 93440 69940 93492
rect 69992 93480 69998 93492
rect 70854 93480 70860 93492
rect 69992 93452 70860 93480
rect 69992 93440 69998 93452
rect 70854 93440 70860 93452
rect 70912 93440 70918 93492
rect 71682 93440 71688 93492
rect 71740 93480 71746 93492
rect 72697 93483 72755 93489
rect 72697 93480 72709 93483
rect 71740 93452 72709 93480
rect 71740 93440 71746 93452
rect 72697 93449 72709 93452
rect 72743 93449 72755 93483
rect 72697 93443 72755 93449
rect 72970 93440 72976 93492
rect 73028 93440 73034 93492
rect 74718 93440 74724 93492
rect 74776 93440 74782 93492
rect 56284 93384 57836 93412
rect 56284 93372 56290 93384
rect 58894 93372 58900 93424
rect 58952 93412 58958 93424
rect 59538 93412 59544 93424
rect 58952 93384 59544 93412
rect 58952 93372 58958 93384
rect 59538 93372 59544 93384
rect 59596 93412 59602 93424
rect 60734 93412 60740 93424
rect 59596 93384 60740 93412
rect 59596 93372 59602 93384
rect 46109 93347 46167 93353
rect 46109 93313 46121 93347
rect 46155 93344 46167 93347
rect 46155 93316 46336 93344
rect 46155 93313 46167 93316
rect 46109 93307 46167 93313
rect 46308 93285 46336 93316
rect 49326 93304 49332 93356
rect 49384 93344 49390 93356
rect 49769 93347 49827 93353
rect 49769 93344 49781 93347
rect 49384 93316 49781 93344
rect 49384 93304 49390 93316
rect 49769 93313 49781 93316
rect 49815 93313 49827 93347
rect 54113 93347 54171 93353
rect 54113 93344 54125 93347
rect 49769 93307 49827 93313
rect 50540 93316 54125 93344
rect 46293 93279 46351 93285
rect 46293 93245 46305 93279
rect 46339 93276 46351 93279
rect 46842 93276 46848 93288
rect 46339 93248 46848 93276
rect 46339 93245 46351 93248
rect 46293 93239 46351 93245
rect 46842 93236 46848 93248
rect 46900 93276 46906 93288
rect 46937 93279 46995 93285
rect 46937 93276 46949 93279
rect 46900 93248 46949 93276
rect 46900 93236 46906 93248
rect 46937 93245 46949 93248
rect 46983 93276 46995 93279
rect 47121 93279 47179 93285
rect 47121 93276 47133 93279
rect 46983 93248 47133 93276
rect 46983 93245 46995 93248
rect 46937 93239 46995 93245
rect 47121 93245 47133 93248
rect 47167 93276 47179 93279
rect 49237 93279 49295 93285
rect 49237 93276 49249 93279
rect 47167 93248 49249 93276
rect 47167 93245 47179 93248
rect 47121 93239 47179 93245
rect 49237 93245 49249 93248
rect 49283 93276 49295 93279
rect 49510 93276 49516 93288
rect 49283 93248 49516 93276
rect 49283 93245 49295 93248
rect 49237 93239 49295 93245
rect 49510 93236 49516 93248
rect 49568 93236 49574 93288
rect 49326 93168 49332 93220
rect 49384 93168 49390 93220
rect 46934 93100 46940 93152
rect 46992 93140 46998 93152
rect 50540 93140 50568 93316
rect 54113 93313 54125 93316
rect 54159 93313 54171 93347
rect 54113 93307 54171 93313
rect 54662 93304 54668 93356
rect 54720 93344 54726 93356
rect 56594 93344 56600 93356
rect 54720 93316 56600 93344
rect 54720 93304 54726 93316
rect 56594 93304 56600 93316
rect 56652 93304 56658 93356
rect 57333 93347 57391 93353
rect 57333 93344 57345 93347
rect 56704 93316 57345 93344
rect 53834 93236 53840 93288
rect 53892 93236 53898 93288
rect 53926 93236 53932 93288
rect 53984 93276 53990 93288
rect 56318 93276 56324 93288
rect 53984 93248 56324 93276
rect 53984 93236 53990 93248
rect 56318 93236 56324 93248
rect 56376 93236 56382 93288
rect 56413 93279 56471 93285
rect 56413 93245 56425 93279
rect 56459 93276 56471 93279
rect 56502 93276 56508 93288
rect 56459 93248 56508 93276
rect 56459 93245 56471 93248
rect 56413 93239 56471 93245
rect 56502 93236 56508 93248
rect 56560 93236 56566 93288
rect 50893 93211 50951 93217
rect 50893 93177 50905 93211
rect 50939 93208 50951 93211
rect 56704 93208 56732 93316
rect 57333 93313 57345 93316
rect 57379 93313 57391 93347
rect 57333 93307 57391 93313
rect 59653 93347 59711 93353
rect 59653 93313 59665 93347
rect 59699 93344 59711 93347
rect 59814 93344 59820 93356
rect 59699 93316 59820 93344
rect 59699 93313 59711 93316
rect 59653 93307 59711 93313
rect 59814 93304 59820 93316
rect 59872 93304 59878 93356
rect 59924 93353 59952 93384
rect 60734 93372 60740 93384
rect 60792 93412 60798 93424
rect 63586 93412 63592 93424
rect 60792 93384 61424 93412
rect 60792 93372 60798 93384
rect 61396 93353 61424 93384
rect 62868 93384 63592 93412
rect 62868 93353 62896 93384
rect 63586 93372 63592 93384
rect 63644 93412 63650 93424
rect 66898 93412 66904 93424
rect 63644 93384 66904 93412
rect 63644 93372 63650 93384
rect 59909 93347 59967 93353
rect 59909 93313 59921 93347
rect 59955 93313 59967 93347
rect 59909 93307 59967 93313
rect 61125 93347 61183 93353
rect 61125 93313 61137 93347
rect 61171 93344 61183 93347
rect 61381 93347 61439 93353
rect 61171 93316 61332 93344
rect 61171 93313 61183 93316
rect 61125 93307 61183 93313
rect 56870 93236 56876 93288
rect 56928 93276 56934 93288
rect 57057 93279 57115 93285
rect 57057 93276 57069 93279
rect 56928 93248 57069 93276
rect 56928 93236 56934 93248
rect 57057 93245 57069 93248
rect 57103 93245 57115 93279
rect 57057 93239 57115 93245
rect 57241 93279 57299 93285
rect 57241 93245 57253 93279
rect 57287 93245 57299 93279
rect 61304 93276 61332 93316
rect 61381 93313 61393 93347
rect 61427 93313 61439 93347
rect 61381 93307 61439 93313
rect 62597 93347 62655 93353
rect 62597 93313 62609 93347
rect 62643 93344 62655 93347
rect 62853 93347 62911 93353
rect 62643 93316 62804 93344
rect 62643 93313 62655 93316
rect 62597 93307 62655 93313
rect 62776 93276 62804 93316
rect 62853 93313 62865 93347
rect 62899 93313 62911 93347
rect 62853 93307 62911 93313
rect 63218 93304 63224 93356
rect 63276 93304 63282 93356
rect 63310 93304 63316 93356
rect 63368 93304 63374 93356
rect 64800 93353 64828 93384
rect 66272 93353 66300 93384
rect 66898 93372 66904 93384
rect 66956 93372 66962 93424
rect 68370 93372 68376 93424
rect 68428 93412 68434 93424
rect 70118 93412 70124 93424
rect 68428 93384 70124 93412
rect 68428 93372 68434 93384
rect 64529 93347 64587 93353
rect 64529 93313 64541 93347
rect 64575 93344 64587 93347
rect 64785 93347 64843 93353
rect 64575 93316 64736 93344
rect 64575 93313 64587 93316
rect 64529 93307 64587 93313
rect 63770 93276 63776 93288
rect 61304 93248 61884 93276
rect 62776 93248 63776 93276
rect 57241 93239 57299 93245
rect 50939 93180 56732 93208
rect 57256 93208 57284 93239
rect 58529 93211 58587 93217
rect 58529 93208 58541 93211
rect 57256 93180 58541 93208
rect 50939 93177 50951 93180
rect 50893 93171 50951 93177
rect 58529 93177 58541 93180
rect 58575 93177 58587 93211
rect 58529 93171 58587 93177
rect 46992 93112 50568 93140
rect 46992 93100 46998 93112
rect 52178 93100 52184 93152
rect 52236 93140 52242 93152
rect 56226 93140 56232 93152
rect 52236 93112 56232 93140
rect 52236 93100 52242 93112
rect 56226 93100 56232 93112
rect 56284 93100 56290 93152
rect 56318 93100 56324 93152
rect 56376 93140 56382 93152
rect 60366 93140 60372 93152
rect 56376 93112 60372 93140
rect 56376 93100 56382 93112
rect 60366 93100 60372 93112
rect 60424 93100 60430 93152
rect 60458 93100 60464 93152
rect 60516 93140 60522 93152
rect 61654 93140 61660 93152
rect 60516 93112 61660 93140
rect 60516 93100 60522 93112
rect 61654 93100 61660 93112
rect 61712 93100 61718 93152
rect 61856 93140 61884 93248
rect 63770 93236 63776 93248
rect 63828 93236 63834 93288
rect 64708 93276 64736 93316
rect 64785 93313 64797 93347
rect 64831 93313 64843 93347
rect 64785 93307 64843 93313
rect 66001 93347 66059 93353
rect 66001 93313 66013 93347
rect 66047 93344 66059 93347
rect 66257 93347 66315 93353
rect 66047 93316 66208 93344
rect 66047 93313 66059 93316
rect 66001 93307 66059 93313
rect 65242 93276 65248 93288
rect 64708 93248 65248 93276
rect 65242 93236 65248 93248
rect 65300 93236 65306 93288
rect 66180 93276 66208 93316
rect 66257 93313 66269 93347
rect 66303 93313 66315 93347
rect 66257 93307 66315 93313
rect 66346 93304 66352 93356
rect 66404 93344 66410 93356
rect 66404 93316 66484 93344
rect 66404 93304 66410 93316
rect 66456 93285 66484 93316
rect 66714 93304 66720 93356
rect 66772 93304 66778 93356
rect 67818 93304 67824 93356
rect 67876 93344 67882 93356
rect 68557 93347 68615 93353
rect 68557 93344 68569 93347
rect 67876 93316 68569 93344
rect 67876 93304 67882 93316
rect 68557 93313 68569 93316
rect 68603 93313 68615 93347
rect 68557 93307 68615 93313
rect 66441 93279 66499 93285
rect 66180 93248 66392 93276
rect 64782 93168 64788 93220
rect 64840 93208 64846 93220
rect 66364 93208 66392 93248
rect 66441 93245 66453 93279
rect 66487 93276 66499 93279
rect 68370 93276 68376 93288
rect 66487 93248 68376 93276
rect 66487 93245 66499 93248
rect 66441 93239 66499 93245
rect 68370 93236 68376 93248
rect 68428 93236 68434 93288
rect 69124 93285 69152 93384
rect 70118 93372 70124 93384
rect 70176 93372 70182 93424
rect 70213 93415 70271 93421
rect 70213 93381 70225 93415
rect 70259 93412 70271 93415
rect 72050 93412 72056 93424
rect 70259 93384 72056 93412
rect 70259 93381 70271 93384
rect 70213 93375 70271 93381
rect 72050 93372 72056 93384
rect 72108 93372 72114 93424
rect 72234 93372 72240 93424
rect 72292 93412 72298 93424
rect 72421 93415 72479 93421
rect 72292 93384 72372 93412
rect 72292 93372 72298 93384
rect 69198 93304 69204 93356
rect 69256 93344 69262 93356
rect 69385 93347 69443 93353
rect 69385 93344 69397 93347
rect 69256 93316 69397 93344
rect 69256 93304 69262 93316
rect 69385 93313 69397 93316
rect 69431 93313 69443 93347
rect 69385 93307 69443 93313
rect 70302 93304 70308 93356
rect 70360 93304 70366 93356
rect 71889 93347 71947 93353
rect 71889 93313 71901 93347
rect 71935 93344 71947 93347
rect 72344 93344 72372 93384
rect 72421 93381 72433 93415
rect 72467 93412 72479 93415
rect 72467 93384 73108 93412
rect 72467 93381 72479 93384
rect 72421 93375 72479 93381
rect 73080 93353 73108 93384
rect 73908 93384 75224 93412
rect 73908 93353 73936 93384
rect 72605 93347 72663 93353
rect 72605 93344 72617 93347
rect 71935 93316 72280 93344
rect 72344 93316 72617 93344
rect 71935 93313 71947 93316
rect 71889 93307 71947 93313
rect 68465 93279 68523 93285
rect 68465 93245 68477 93279
rect 68511 93276 68523 93279
rect 69109 93279 69167 93285
rect 68511 93248 69060 93276
rect 68511 93245 68523 93248
rect 68465 93239 68523 93245
rect 66806 93208 66812 93220
rect 64840 93180 65380 93208
rect 66364 93180 66812 93208
rect 64840 93168 64846 93180
rect 62850 93140 62856 93152
rect 61856 93112 62856 93140
rect 62850 93100 62856 93112
rect 62908 93100 62914 93152
rect 63402 93100 63408 93152
rect 63460 93140 63466 93152
rect 64877 93143 64935 93149
rect 64877 93140 64889 93143
rect 63460 93112 64889 93140
rect 63460 93100 63466 93112
rect 64877 93109 64889 93112
rect 64923 93109 64935 93143
rect 65352 93140 65380 93180
rect 66806 93168 66812 93180
rect 66864 93168 66870 93220
rect 67085 93211 67143 93217
rect 67085 93177 67097 93211
rect 67131 93208 67143 93211
rect 67726 93208 67732 93220
rect 67131 93180 67732 93208
rect 67131 93177 67143 93180
rect 67085 93171 67143 93177
rect 67726 93168 67732 93180
rect 67784 93168 67790 93220
rect 69032 93208 69060 93248
rect 69109 93245 69121 93279
rect 69155 93245 69167 93279
rect 69109 93239 69167 93245
rect 69293 93279 69351 93285
rect 69293 93245 69305 93279
rect 69339 93276 69351 93279
rect 69934 93276 69940 93288
rect 69339 93248 69940 93276
rect 69339 93245 69351 93248
rect 69293 93239 69351 93245
rect 69934 93236 69940 93248
rect 69992 93236 69998 93288
rect 70118 93236 70124 93288
rect 70176 93236 70182 93288
rect 72142 93236 72148 93288
rect 72200 93236 72206 93288
rect 72252 93276 72280 93316
rect 72605 93313 72617 93316
rect 72651 93313 72663 93347
rect 72605 93307 72663 93313
rect 73065 93347 73123 93353
rect 73065 93313 73077 93347
rect 73111 93344 73123 93347
rect 73433 93347 73491 93353
rect 73433 93344 73445 93347
rect 73111 93316 73445 93344
rect 73111 93313 73123 93316
rect 73065 93307 73123 93313
rect 73433 93313 73445 93316
rect 73479 93344 73491 93347
rect 73617 93347 73675 93353
rect 73617 93344 73629 93347
rect 73479 93316 73629 93344
rect 73479 93313 73491 93316
rect 73433 93307 73491 93313
rect 73617 93313 73629 93316
rect 73663 93344 73675 93347
rect 73893 93347 73951 93353
rect 73893 93344 73905 93347
rect 73663 93316 73905 93344
rect 73663 93313 73675 93316
rect 73617 93307 73675 93313
rect 73893 93313 73905 93316
rect 73939 93313 73951 93347
rect 73893 93307 73951 93313
rect 74445 93347 74503 93353
rect 74445 93313 74457 93347
rect 74491 93344 74503 93347
rect 74813 93347 74871 93353
rect 74813 93344 74825 93347
rect 74491 93316 74825 93344
rect 74491 93313 74503 93316
rect 74445 93307 74503 93313
rect 74813 93313 74825 93316
rect 74859 93344 74871 93347
rect 74859 93316 75040 93344
rect 74859 93313 74871 93316
rect 74813 93307 74871 93313
rect 74166 93276 74172 93288
rect 72252 93248 74172 93276
rect 74166 93236 74172 93248
rect 74224 93236 74230 93288
rect 75012 93217 75040 93316
rect 75196 93285 75224 93384
rect 75181 93279 75239 93285
rect 75181 93245 75193 93279
rect 75227 93276 75239 93279
rect 75227 93248 84194 93276
rect 75227 93245 75239 93248
rect 75181 93239 75239 93245
rect 70765 93211 70823 93217
rect 70765 93208 70777 93211
rect 69032 93180 70777 93208
rect 70765 93177 70777 93180
rect 70811 93177 70823 93211
rect 70765 93171 70823 93177
rect 74997 93211 75055 93217
rect 74997 93177 75009 93211
rect 75043 93208 75055 93211
rect 84166 93208 84194 93248
rect 107838 93208 107844 93220
rect 75043 93180 75408 93208
rect 84166 93180 107844 93208
rect 75043 93177 75055 93180
rect 74997 93171 75055 93177
rect 68554 93140 68560 93152
rect 65352 93112 68560 93140
rect 64877 93103 64935 93109
rect 68554 93100 68560 93112
rect 68612 93100 68618 93152
rect 68925 93143 68983 93149
rect 68925 93109 68937 93143
rect 68971 93140 68983 93143
rect 69014 93140 69020 93152
rect 68971 93112 69020 93140
rect 68971 93109 68983 93112
rect 68925 93103 68983 93109
rect 69014 93100 69020 93112
rect 69072 93100 69078 93152
rect 69750 93100 69756 93152
rect 69808 93100 69814 93152
rect 69842 93100 69848 93152
rect 69900 93140 69906 93152
rect 70578 93140 70584 93152
rect 69900 93112 70584 93140
rect 69900 93100 69906 93112
rect 70578 93100 70584 93112
rect 70636 93100 70642 93152
rect 70673 93143 70731 93149
rect 70673 93109 70685 93143
rect 70719 93140 70731 93143
rect 71958 93140 71964 93152
rect 70719 93112 71964 93140
rect 70719 93109 70731 93112
rect 70673 93103 70731 93109
rect 71958 93100 71964 93112
rect 72016 93100 72022 93152
rect 75380 93149 75408 93180
rect 107838 93168 107844 93180
rect 107896 93168 107902 93220
rect 75365 93143 75423 93149
rect 75365 93109 75377 93143
rect 75411 93140 75423 93143
rect 108574 93140 108580 93152
rect 75411 93112 108580 93140
rect 75411 93109 75423 93112
rect 75365 93103 75423 93109
rect 108574 93100 108580 93112
rect 108632 93100 108638 93152
rect 1104 93050 118864 93072
rect 1104 92998 4214 93050
rect 4266 92998 4278 93050
rect 4330 92998 4342 93050
rect 4394 92998 4406 93050
rect 4458 92998 4470 93050
rect 4522 92998 34934 93050
rect 34986 92998 34998 93050
rect 35050 92998 35062 93050
rect 35114 92998 35126 93050
rect 35178 92998 35190 93050
rect 35242 92998 65654 93050
rect 65706 92998 65718 93050
rect 65770 92998 65782 93050
rect 65834 92998 65846 93050
rect 65898 92998 65910 93050
rect 65962 92998 96374 93050
rect 96426 92998 96438 93050
rect 96490 92998 96502 93050
rect 96554 92998 96566 93050
rect 96618 92998 96630 93050
rect 96682 92998 118864 93050
rect 1104 92976 118864 92998
rect 46934 92896 46940 92948
rect 46992 92896 46998 92948
rect 48409 92939 48467 92945
rect 48409 92905 48421 92939
rect 48455 92936 48467 92939
rect 48455 92908 51764 92936
rect 48455 92905 48467 92908
rect 48409 92899 48467 92905
rect 51736 92868 51764 92908
rect 52178 92896 52184 92948
rect 52236 92896 52242 92948
rect 52454 92936 52460 92948
rect 52288 92908 52460 92936
rect 52288 92868 52316 92908
rect 52454 92896 52460 92908
rect 52512 92896 52518 92948
rect 53653 92939 53711 92945
rect 53653 92905 53665 92939
rect 53699 92936 53711 92939
rect 53926 92936 53932 92948
rect 53699 92908 53932 92936
rect 53699 92905 53711 92908
rect 53653 92899 53711 92905
rect 53926 92896 53932 92908
rect 53984 92896 53990 92948
rect 55125 92939 55183 92945
rect 55125 92905 55137 92939
rect 55171 92936 55183 92939
rect 55171 92908 55352 92936
rect 55171 92905 55183 92908
rect 55125 92899 55183 92905
rect 51736 92840 52316 92868
rect 55324 92868 55352 92908
rect 55398 92896 55404 92948
rect 55456 92936 55462 92948
rect 56505 92939 56563 92945
rect 56505 92936 56517 92939
rect 55456 92908 56517 92936
rect 55456 92896 55462 92908
rect 56505 92905 56517 92908
rect 56551 92905 56563 92939
rect 59541 92939 59599 92945
rect 56505 92899 56563 92905
rect 56612 92908 59124 92936
rect 56612 92868 56640 92908
rect 55324 92840 56640 92868
rect 59096 92868 59124 92908
rect 59541 92905 59553 92939
rect 59587 92936 59599 92939
rect 61286 92936 61292 92948
rect 59587 92908 61292 92936
rect 59587 92905 59599 92908
rect 59541 92899 59599 92905
rect 61286 92896 61292 92908
rect 61344 92896 61350 92948
rect 61378 92896 61384 92948
rect 61436 92936 61442 92948
rect 63402 92936 63408 92948
rect 61436 92908 63408 92936
rect 61436 92896 61442 92908
rect 63402 92896 63408 92908
rect 63460 92896 63466 92948
rect 63494 92896 63500 92948
rect 63552 92896 63558 92948
rect 65613 92939 65671 92945
rect 65613 92936 65625 92939
rect 63604 92908 65625 92936
rect 60458 92868 60464 92880
rect 59096 92840 60464 92868
rect 60458 92828 60464 92840
rect 60516 92828 60522 92880
rect 62942 92828 62948 92880
rect 63000 92868 63006 92880
rect 63604 92868 63632 92908
rect 65613 92905 65625 92908
rect 65659 92905 65671 92939
rect 67085 92939 67143 92945
rect 67085 92936 67097 92939
rect 65613 92899 65671 92905
rect 65720 92908 67097 92936
rect 63000 92840 63632 92868
rect 63000 92828 63006 92840
rect 64598 92828 64604 92880
rect 64656 92868 64662 92880
rect 65720 92868 65748 92908
rect 67085 92905 67097 92908
rect 67131 92905 67143 92939
rect 70302 92936 70308 92948
rect 67085 92899 67143 92905
rect 67560 92908 70308 92936
rect 67560 92868 67588 92908
rect 70302 92896 70308 92908
rect 70360 92896 70366 92948
rect 70578 92896 70584 92948
rect 70636 92936 70642 92948
rect 70765 92939 70823 92945
rect 70765 92936 70777 92939
rect 70636 92908 70777 92936
rect 70636 92896 70642 92908
rect 70765 92905 70777 92908
rect 70811 92905 70823 92939
rect 72237 92939 72295 92945
rect 72237 92936 72249 92939
rect 70765 92899 70823 92905
rect 71240 92908 72249 92936
rect 64656 92840 65748 92868
rect 67468 92840 67588 92868
rect 64656 92828 64662 92840
rect 46842 92760 46848 92812
rect 46900 92800 46906 92812
rect 47029 92803 47087 92809
rect 47029 92800 47041 92803
rect 46900 92772 47041 92800
rect 46900 92760 46906 92772
rect 47029 92769 47041 92772
rect 47075 92769 47087 92803
rect 47029 92763 47087 92769
rect 50614 92760 50620 92812
rect 50672 92760 50678 92812
rect 57974 92760 57980 92812
rect 58032 92760 58038 92812
rect 63586 92760 63592 92812
rect 63644 92760 63650 92812
rect 67468 92800 67496 92840
rect 68554 92828 68560 92880
rect 68612 92828 68618 92880
rect 69934 92828 69940 92880
rect 69992 92868 69998 92880
rect 71240 92868 71268 92908
rect 72237 92905 72249 92908
rect 72283 92905 72295 92939
rect 72237 92899 72295 92905
rect 69992 92840 71268 92868
rect 69992 92828 69998 92840
rect 66916 92772 67496 92800
rect 45557 92735 45615 92741
rect 45557 92701 45569 92735
rect 45603 92732 45615 92735
rect 45646 92732 45652 92744
rect 45603 92704 45652 92732
rect 45603 92701 45615 92704
rect 45557 92695 45615 92701
rect 45646 92692 45652 92704
rect 45704 92732 45710 92744
rect 46860 92732 46888 92760
rect 45704 92704 46888 92732
rect 45704 92692 45710 92704
rect 44174 92624 44180 92676
rect 44232 92664 44238 92676
rect 45373 92667 45431 92673
rect 45373 92664 45385 92667
rect 44232 92636 45385 92664
rect 44232 92624 44238 92636
rect 45373 92633 45385 92636
rect 45419 92664 45431 92667
rect 45802 92667 45860 92673
rect 45802 92664 45814 92667
rect 45419 92636 45814 92664
rect 45419 92633 45431 92636
rect 45373 92627 45431 92633
rect 45802 92633 45814 92636
rect 45848 92633 45860 92667
rect 45802 92627 45860 92633
rect 47118 92624 47124 92676
rect 47176 92664 47182 92676
rect 47274 92667 47332 92673
rect 47274 92664 47286 92667
rect 47176 92636 47286 92664
rect 47176 92624 47182 92636
rect 47274 92633 47286 92636
rect 47320 92664 47332 92667
rect 48501 92667 48559 92673
rect 48501 92664 48513 92667
rect 47320 92636 48513 92664
rect 47320 92633 47332 92636
rect 47274 92627 47332 92633
rect 48501 92633 48513 92636
rect 48547 92633 48559 92667
rect 50632 92664 50660 92760
rect 50801 92735 50859 92741
rect 50801 92701 50813 92735
rect 50847 92732 50859 92735
rect 52273 92735 52331 92741
rect 52273 92732 52285 92735
rect 50847 92704 52285 92732
rect 50847 92701 50859 92704
rect 50801 92695 50859 92701
rect 52273 92701 52285 92704
rect 52319 92732 52331 92735
rect 53374 92732 53380 92744
rect 52319 92704 53380 92732
rect 52319 92701 52331 92704
rect 52273 92695 52331 92701
rect 53374 92692 53380 92704
rect 53432 92732 53438 92744
rect 53745 92735 53803 92741
rect 53745 92732 53757 92735
rect 53432 92704 53757 92732
rect 53432 92692 53438 92704
rect 53745 92701 53757 92704
rect 53791 92701 53803 92735
rect 55493 92735 55551 92741
rect 55493 92732 55505 92735
rect 53745 92695 53803 92701
rect 55186 92704 55505 92732
rect 52546 92673 52552 92676
rect 51046 92667 51104 92673
rect 51046 92664 51058 92667
rect 50632 92636 51058 92664
rect 48501 92627 48559 92633
rect 51046 92633 51058 92636
rect 51092 92633 51104 92667
rect 52540 92664 52552 92673
rect 52507 92636 52552 92664
rect 51046 92627 51104 92633
rect 52540 92627 52552 92636
rect 52546 92624 52552 92627
rect 52604 92624 52610 92676
rect 54018 92673 54024 92676
rect 54012 92664 54024 92673
rect 53979 92636 54024 92664
rect 54012 92627 54024 92636
rect 54076 92664 54082 92676
rect 55186 92664 55214 92704
rect 55493 92701 55505 92704
rect 55539 92701 55551 92735
rect 55493 92695 55551 92701
rect 56502 92692 56508 92744
rect 56560 92732 56566 92744
rect 57885 92735 57943 92741
rect 57885 92732 57897 92735
rect 56560 92704 57897 92732
rect 56560 92692 56566 92704
rect 57885 92701 57897 92704
rect 57931 92701 57943 92735
rect 57885 92695 57943 92701
rect 58161 92735 58219 92741
rect 58161 92701 58173 92735
rect 58207 92732 58219 92735
rect 58894 92732 58900 92744
rect 58207 92704 58900 92732
rect 58207 92701 58219 92704
rect 58161 92695 58219 92701
rect 58894 92692 58900 92704
rect 58952 92692 58958 92744
rect 61933 92735 61991 92741
rect 61933 92701 61945 92735
rect 61979 92732 61991 92735
rect 63604 92732 63632 92760
rect 66916 92732 66944 92772
rect 61979 92704 63632 92732
rect 66640 92704 66944 92732
rect 66993 92735 67051 92741
rect 61979 92701 61991 92704
rect 61933 92695 61991 92701
rect 58434 92673 58440 92676
rect 54076 92636 55214 92664
rect 57640 92667 57698 92673
rect 54018 92624 54024 92627
rect 54076 92624 54082 92636
rect 57640 92633 57652 92667
rect 57686 92664 57698 92667
rect 57686 92636 58388 92664
rect 57686 92633 57698 92636
rect 57640 92627 57698 92633
rect 52564 92596 52592 92624
rect 55309 92599 55367 92605
rect 55309 92596 55321 92599
rect 52564 92568 55321 92596
rect 55309 92565 55321 92568
rect 55355 92565 55367 92599
rect 58360 92596 58388 92636
rect 58428 92627 58440 92673
rect 58492 92664 58498 92676
rect 58492 92636 58528 92664
rect 58434 92624 58440 92627
rect 58492 92624 58498 92636
rect 59262 92624 59268 92676
rect 59320 92664 59326 92676
rect 61749 92667 61807 92673
rect 61749 92664 61761 92667
rect 59320 92636 61761 92664
rect 59320 92624 59326 92636
rect 61749 92633 61761 92636
rect 61795 92664 61807 92667
rect 62178 92667 62236 92673
rect 62178 92664 62190 92667
rect 61795 92636 62190 92664
rect 61795 92633 61807 92636
rect 61749 92627 61807 92633
rect 62178 92633 62190 92636
rect 62224 92633 62236 92667
rect 62178 92627 62236 92633
rect 63218 92624 63224 92676
rect 63276 92624 63282 92676
rect 63494 92624 63500 92676
rect 63552 92664 63558 92676
rect 63834 92667 63892 92673
rect 63834 92664 63846 92667
rect 63552 92636 63846 92664
rect 63552 92624 63558 92636
rect 63834 92633 63846 92636
rect 63880 92633 63892 92667
rect 63834 92627 63892 92633
rect 59446 92596 59452 92608
rect 58360 92568 59452 92596
rect 55309 92559 55367 92565
rect 59446 92556 59452 92568
rect 59504 92556 59510 92608
rect 61286 92556 61292 92608
rect 61344 92596 61350 92608
rect 63236 92596 63264 92624
rect 61344 92568 63264 92596
rect 63313 92599 63371 92605
rect 61344 92556 61350 92568
rect 63313 92565 63325 92599
rect 63359 92596 63371 92599
rect 64874 92596 64880 92608
rect 63359 92568 64880 92596
rect 63359 92565 63371 92568
rect 63313 92559 63371 92565
rect 64874 92556 64880 92568
rect 64932 92556 64938 92608
rect 64969 92599 65027 92605
rect 64969 92565 64981 92599
rect 65015 92596 65027 92599
rect 66640 92596 66668 92704
rect 66993 92701 67005 92735
rect 67039 92732 67051 92735
rect 68465 92735 68523 92741
rect 68465 92732 68477 92735
rect 67039 92704 68477 92732
rect 67039 92701 67051 92704
rect 66993 92695 67051 92701
rect 68465 92701 68477 92704
rect 68511 92732 68523 92735
rect 69937 92735 69995 92741
rect 69937 92732 69949 92735
rect 68511 92704 69949 92732
rect 68511 92701 68523 92704
rect 68465 92695 68523 92701
rect 69584 92676 69612 92704
rect 69937 92701 69949 92704
rect 69983 92701 69995 92735
rect 69937 92695 69995 92701
rect 72142 92692 72148 92744
rect 72200 92732 72206 92744
rect 72970 92732 72976 92744
rect 72200 92704 72976 92732
rect 72200 92692 72206 92704
rect 72970 92692 72976 92704
rect 73028 92732 73034 92744
rect 73617 92735 73675 92741
rect 73617 92732 73629 92735
rect 73028 92704 73629 92732
rect 73028 92692 73034 92704
rect 73617 92701 73629 92704
rect 73663 92732 73675 92735
rect 73663 92704 73844 92732
rect 73663 92701 73675 92704
rect 73617 92695 73675 92701
rect 66748 92667 66806 92673
rect 66748 92633 66760 92667
rect 66794 92664 66806 92667
rect 67542 92664 67548 92676
rect 66794 92636 67548 92664
rect 66794 92633 66806 92636
rect 66748 92627 66806 92633
rect 67542 92624 67548 92636
rect 67600 92624 67606 92676
rect 68220 92667 68278 92673
rect 68220 92633 68232 92667
rect 68266 92664 68278 92667
rect 69198 92664 69204 92676
rect 68266 92636 69204 92664
rect 68266 92633 68278 92636
rect 68220 92627 68278 92633
rect 69198 92624 69204 92636
rect 69256 92624 69262 92676
rect 69566 92624 69572 92676
rect 69624 92624 69630 92676
rect 69692 92667 69750 92673
rect 69692 92633 69704 92667
rect 69738 92664 69750 92667
rect 70486 92664 70492 92676
rect 69738 92636 70492 92664
rect 69738 92633 69750 92636
rect 69692 92627 69750 92633
rect 70486 92624 70492 92636
rect 70544 92624 70550 92676
rect 71900 92667 71958 92673
rect 71900 92633 71912 92667
rect 71946 92664 71958 92667
rect 73246 92664 73252 92676
rect 71946 92636 73252 92664
rect 71946 92633 71958 92636
rect 71900 92627 71958 92633
rect 73246 92624 73252 92636
rect 73304 92624 73310 92676
rect 73372 92667 73430 92673
rect 73372 92633 73384 92667
rect 73418 92664 73430 92667
rect 73706 92664 73712 92676
rect 73418 92636 73712 92664
rect 73418 92633 73430 92636
rect 73372 92627 73430 92633
rect 73706 92624 73712 92636
rect 73764 92624 73770 92676
rect 73816 92605 73844 92704
rect 77389 92667 77447 92673
rect 77389 92633 77401 92667
rect 77435 92664 77447 92667
rect 77478 92664 77484 92676
rect 77435 92636 77484 92664
rect 77435 92633 77447 92636
rect 77389 92627 77447 92633
rect 77478 92624 77484 92636
rect 77536 92624 77542 92676
rect 79229 92667 79287 92673
rect 79229 92633 79241 92667
rect 79275 92633 79287 92667
rect 79229 92627 79287 92633
rect 65015 92568 66668 92596
rect 73801 92599 73859 92605
rect 65015 92565 65027 92568
rect 64969 92559 65027 92565
rect 73801 92565 73813 92599
rect 73847 92596 73859 92599
rect 74718 92596 74724 92608
rect 73847 92568 74724 92596
rect 73847 92565 73859 92568
rect 73801 92559 73859 92565
rect 74718 92556 74724 92568
rect 74776 92556 74782 92608
rect 79244 92596 79272 92627
rect 79410 92596 79416 92608
rect 79244 92568 79416 92596
rect 79410 92556 79416 92568
rect 79468 92556 79474 92608
rect 1104 92506 118864 92528
rect 1104 92454 4874 92506
rect 4926 92454 4938 92506
rect 4990 92454 5002 92506
rect 5054 92454 5066 92506
rect 5118 92454 5130 92506
rect 5182 92454 35594 92506
rect 35646 92454 35658 92506
rect 35710 92454 35722 92506
rect 35774 92454 35786 92506
rect 35838 92454 35850 92506
rect 35902 92454 66314 92506
rect 66366 92454 66378 92506
rect 66430 92454 66442 92506
rect 66494 92454 66506 92506
rect 66558 92454 66570 92506
rect 66622 92454 97034 92506
rect 97086 92454 97098 92506
rect 97150 92454 97162 92506
rect 97214 92454 97226 92506
rect 97278 92454 97290 92506
rect 97342 92454 113650 92506
rect 113702 92454 113714 92506
rect 113766 92454 113778 92506
rect 113830 92454 113842 92506
rect 113894 92454 113906 92506
rect 113958 92454 118864 92506
rect 1104 92432 118864 92454
rect 45646 92352 45652 92404
rect 45704 92352 45710 92404
rect 47121 92395 47179 92401
rect 47121 92392 47133 92395
rect 46952 92364 47133 92392
rect 46952 92265 46980 92364
rect 47121 92361 47133 92364
rect 47167 92392 47179 92395
rect 54662 92392 54668 92404
rect 47167 92364 54668 92392
rect 47167 92361 47179 92364
rect 47121 92355 47179 92361
rect 54662 92352 54668 92364
rect 54720 92352 54726 92404
rect 54757 92395 54815 92401
rect 54757 92361 54769 92395
rect 54803 92361 54815 92395
rect 54757 92355 54815 92361
rect 47305 92327 47363 92333
rect 47305 92293 47317 92327
rect 47351 92324 47363 92327
rect 47949 92327 48007 92333
rect 47949 92324 47961 92327
rect 47351 92296 47961 92324
rect 47351 92293 47363 92296
rect 47305 92287 47363 92293
rect 47949 92293 47961 92296
rect 47995 92324 48007 92327
rect 47995 92296 49556 92324
rect 47995 92293 48007 92296
rect 47949 92287 48007 92293
rect 48240 92265 48268 92296
rect 49528 92268 49556 92296
rect 52914 92284 52920 92336
rect 52972 92324 52978 92336
rect 54772 92324 54800 92355
rect 54846 92352 54852 92404
rect 54904 92392 54910 92404
rect 58342 92392 58348 92404
rect 54904 92364 58348 92392
rect 54904 92352 54910 92364
rect 58342 92352 58348 92364
rect 58400 92352 58406 92404
rect 60277 92395 60335 92401
rect 60277 92361 60289 92395
rect 60323 92361 60335 92395
rect 60277 92355 60335 92361
rect 56042 92324 56048 92336
rect 52972 92296 53788 92324
rect 54772 92296 56048 92324
rect 52972 92284 52978 92296
rect 46937 92259 46995 92265
rect 46937 92225 46949 92259
rect 46983 92225 46995 92259
rect 46937 92219 46995 92225
rect 48225 92259 48283 92265
rect 48225 92225 48237 92259
rect 48271 92225 48283 92259
rect 48481 92259 48539 92265
rect 48481 92256 48493 92259
rect 48225 92219 48283 92225
rect 48332 92228 48493 92256
rect 48332 92188 48360 92228
rect 48481 92225 48493 92228
rect 48527 92225 48539 92259
rect 48481 92219 48539 92225
rect 49510 92216 49516 92268
rect 49568 92256 49574 92268
rect 49973 92259 50031 92265
rect 49973 92256 49985 92259
rect 49568 92228 49985 92256
rect 49568 92216 49574 92228
rect 49973 92225 49985 92228
rect 50019 92256 50031 92259
rect 50433 92259 50491 92265
rect 50433 92256 50445 92259
rect 50019 92228 50445 92256
rect 50019 92225 50031 92228
rect 49973 92219 50031 92225
rect 50433 92225 50445 92228
rect 50479 92225 50491 92259
rect 50689 92259 50747 92265
rect 50689 92256 50701 92259
rect 50433 92219 50491 92225
rect 50540 92228 50701 92256
rect 50540 92188 50568 92228
rect 50689 92225 50701 92228
rect 50735 92225 50747 92259
rect 50689 92219 50747 92225
rect 53374 92216 53380 92268
rect 53432 92216 53438 92268
rect 53633 92259 53691 92265
rect 53633 92256 53645 92259
rect 53484 92228 53645 92256
rect 48056 92160 48360 92188
rect 50264 92160 50568 92188
rect 8202 92012 8208 92064
rect 8260 92052 8266 92064
rect 45646 92052 45652 92064
rect 8260 92024 45652 92052
rect 8260 92012 8266 92024
rect 45646 92012 45652 92024
rect 45704 92012 45710 92064
rect 46842 92012 46848 92064
rect 46900 92052 46906 92064
rect 48056 92061 48084 92160
rect 50264 92132 50292 92160
rect 53190 92148 53196 92200
rect 53248 92188 53254 92200
rect 53484 92188 53512 92228
rect 53633 92225 53645 92228
rect 53679 92225 53691 92259
rect 53760 92256 53788 92296
rect 56042 92284 56048 92296
rect 56100 92284 56106 92336
rect 56566 92327 56624 92333
rect 56566 92324 56578 92327
rect 56152 92296 56578 92324
rect 56152 92265 56180 92296
rect 56566 92293 56578 92296
rect 56612 92293 56624 92327
rect 60292 92324 60320 92355
rect 63494 92352 63500 92404
rect 63552 92392 63558 92404
rect 65061 92395 65119 92401
rect 65061 92392 65073 92395
rect 63552 92364 65073 92392
rect 63552 92352 63558 92364
rect 60292 92296 63724 92324
rect 56566 92287 56624 92293
rect 56137 92259 56195 92265
rect 56137 92256 56149 92259
rect 53760 92228 56149 92256
rect 53633 92219 53691 92225
rect 56137 92225 56149 92228
rect 56183 92225 56195 92259
rect 56137 92219 56195 92225
rect 56321 92259 56379 92265
rect 56321 92225 56333 92259
rect 56367 92256 56379 92259
rect 56410 92256 56416 92268
rect 56367 92228 56416 92256
rect 56367 92225 56379 92228
rect 56321 92219 56379 92225
rect 56410 92216 56416 92228
rect 56468 92216 56474 92268
rect 58894 92216 58900 92268
rect 58952 92216 58958 92268
rect 59153 92259 59211 92265
rect 59153 92256 59165 92259
rect 59004 92228 59165 92256
rect 59004 92188 59032 92228
rect 59153 92225 59165 92228
rect 59199 92225 59211 92259
rect 59153 92219 59211 92225
rect 60734 92216 60740 92268
rect 60792 92216 60798 92268
rect 60993 92259 61051 92265
rect 60993 92256 61005 92259
rect 60844 92228 61005 92256
rect 60844 92188 60872 92228
rect 60993 92225 61005 92228
rect 61039 92225 61051 92259
rect 60993 92219 61051 92225
rect 53248 92160 53512 92188
rect 58728 92160 59032 92188
rect 60568 92160 60872 92188
rect 63696 92188 63724 92296
rect 64892 92256 64920 92364
rect 65061 92361 65073 92364
rect 65107 92361 65119 92395
rect 65061 92355 65119 92361
rect 65334 92352 65340 92404
rect 65392 92352 65398 92404
rect 67634 92392 67640 92404
rect 66180 92364 67640 92392
rect 64969 92327 65027 92333
rect 64969 92293 64981 92327
rect 65015 92324 65027 92327
rect 65352 92324 65380 92352
rect 65015 92296 65380 92324
rect 65015 92293 65027 92296
rect 64969 92287 65027 92293
rect 66180 92256 66208 92364
rect 67634 92352 67640 92364
rect 67692 92392 67698 92404
rect 67692 92364 70992 92392
rect 67692 92352 67698 92364
rect 70964 92333 70992 92364
rect 72970 92352 72976 92404
rect 73028 92352 73034 92404
rect 77478 92352 77484 92404
rect 77536 92352 77542 92404
rect 69416 92327 69474 92333
rect 69416 92293 69428 92327
rect 69462 92324 69474 92327
rect 70949 92327 71007 92333
rect 69462 92296 70808 92324
rect 69462 92293 69474 92296
rect 69416 92287 69474 92293
rect 64892 92228 66208 92256
rect 69566 92216 69572 92268
rect 69624 92256 69630 92268
rect 69661 92259 69719 92265
rect 69661 92256 69673 92259
rect 69624 92228 69673 92256
rect 69624 92216 69630 92228
rect 69661 92225 69673 92228
rect 69707 92225 69719 92259
rect 69661 92219 69719 92225
rect 70305 92259 70363 92265
rect 70305 92225 70317 92259
rect 70351 92225 70363 92259
rect 70305 92219 70363 92225
rect 66714 92188 66720 92200
rect 63696 92160 66720 92188
rect 53248 92148 53254 92160
rect 58728 92132 58756 92160
rect 60568 92132 60596 92160
rect 66714 92148 66720 92160
rect 66772 92148 66778 92200
rect 50246 92080 50252 92132
rect 50304 92080 50310 92132
rect 51813 92123 51871 92129
rect 51813 92089 51825 92123
rect 51859 92120 51871 92123
rect 51859 92092 53420 92120
rect 51859 92089 51871 92092
rect 51813 92083 51871 92089
rect 48041 92055 48099 92061
rect 48041 92052 48053 92055
rect 46900 92024 48053 92052
rect 46900 92012 46906 92024
rect 48041 92021 48053 92024
rect 48087 92021 48099 92055
rect 48041 92015 48099 92021
rect 49602 92012 49608 92064
rect 49660 92012 49666 92064
rect 53190 92012 53196 92064
rect 53248 92012 53254 92064
rect 53392 92052 53420 92092
rect 58710 92080 58716 92132
rect 58768 92080 58774 92132
rect 60550 92080 60556 92132
rect 60608 92080 60614 92132
rect 62117 92123 62175 92129
rect 62117 92089 62129 92123
rect 62163 92120 62175 92123
rect 67818 92120 67824 92132
rect 62163 92092 67824 92120
rect 62163 92089 62175 92092
rect 62117 92083 62175 92089
rect 67818 92080 67824 92092
rect 67876 92080 67882 92132
rect 68278 92080 68284 92132
rect 68336 92080 68342 92132
rect 69676 92120 69704 92219
rect 70320 92120 70348 92219
rect 70780 92188 70808 92296
rect 70949 92293 70961 92327
rect 70995 92324 71007 92327
rect 72789 92327 72847 92333
rect 72789 92324 72801 92327
rect 70995 92296 72801 92324
rect 70995 92293 71007 92296
rect 70949 92287 71007 92293
rect 72789 92293 72801 92296
rect 72835 92324 72847 92327
rect 77496 92324 77524 92352
rect 72835 92296 77524 92324
rect 72835 92293 72847 92296
rect 72789 92287 72847 92293
rect 74465 92259 74523 92265
rect 74465 92225 74477 92259
rect 74511 92256 74523 92259
rect 74511 92228 74672 92256
rect 74511 92225 74523 92228
rect 74465 92219 74523 92225
rect 71866 92188 71872 92200
rect 70780 92160 71872 92188
rect 71866 92148 71872 92160
rect 71924 92148 71930 92200
rect 74644 92188 74672 92228
rect 74718 92216 74724 92268
rect 74776 92256 74782 92268
rect 74905 92259 74963 92265
rect 74905 92256 74917 92259
rect 74776 92228 74917 92256
rect 74776 92216 74782 92228
rect 74905 92225 74917 92228
rect 74951 92256 74963 92259
rect 77665 92259 77723 92265
rect 77665 92256 77677 92259
rect 74951 92228 77677 92256
rect 74951 92225 74963 92228
rect 74905 92219 74963 92225
rect 77665 92225 77677 92228
rect 77711 92256 77723 92259
rect 77711 92228 77984 92256
rect 77711 92225 77723 92228
rect 77665 92219 77723 92225
rect 75914 92188 75920 92200
rect 74644 92160 75920 92188
rect 75914 92148 75920 92160
rect 75972 92148 75978 92200
rect 70762 92120 70768 92132
rect 69676 92092 70768 92120
rect 70762 92080 70768 92092
rect 70820 92120 70826 92132
rect 71317 92123 71375 92129
rect 71317 92120 71329 92123
rect 70820 92092 71329 92120
rect 70820 92080 70826 92092
rect 71317 92089 71329 92092
rect 71363 92089 71375 92123
rect 71317 92083 71375 92089
rect 72050 92080 72056 92132
rect 72108 92120 72114 92132
rect 73341 92123 73399 92129
rect 73341 92120 73353 92123
rect 72108 92092 73353 92120
rect 72108 92080 72114 92092
rect 73341 92089 73353 92092
rect 73387 92089 73399 92123
rect 73341 92083 73399 92089
rect 54846 92052 54852 92064
rect 53392 92024 54852 92052
rect 54846 92012 54852 92024
rect 54904 92012 54910 92064
rect 57701 92055 57759 92061
rect 57701 92021 57713 92055
rect 57747 92052 57759 92055
rect 64690 92052 64696 92064
rect 57747 92024 64696 92052
rect 57747 92021 57759 92024
rect 57701 92015 57759 92021
rect 64690 92012 64696 92024
rect 64748 92012 64754 92064
rect 77956 92061 77984 92228
rect 100018 92120 100024 92132
rect 84166 92092 100024 92120
rect 77941 92055 77999 92061
rect 77941 92021 77953 92055
rect 77987 92052 77999 92055
rect 79410 92052 79416 92064
rect 77987 92024 79416 92052
rect 77987 92021 77999 92024
rect 77941 92015 77999 92021
rect 79410 92012 79416 92024
rect 79468 92052 79474 92064
rect 84166 92052 84194 92092
rect 100018 92080 100024 92092
rect 100076 92120 100082 92132
rect 100113 92123 100171 92129
rect 100113 92120 100125 92123
rect 100076 92092 100125 92120
rect 100076 92080 100082 92092
rect 100113 92089 100125 92092
rect 100159 92089 100171 92123
rect 100113 92083 100171 92089
rect 79468 92024 84194 92052
rect 79468 92012 79474 92024
rect 89438 92012 89444 92064
rect 89496 92012 89502 92064
rect 1104 91962 118864 91984
rect 1104 91910 4214 91962
rect 4266 91910 4278 91962
rect 4330 91910 4342 91962
rect 4394 91910 4406 91962
rect 4458 91910 4470 91962
rect 4522 91910 34934 91962
rect 34986 91910 34998 91962
rect 35050 91910 35062 91962
rect 35114 91910 35126 91962
rect 35178 91910 35190 91962
rect 35242 91910 65654 91962
rect 65706 91910 65718 91962
rect 65770 91910 65782 91962
rect 65834 91910 65846 91962
rect 65898 91910 65910 91962
rect 65962 91910 96374 91962
rect 96426 91910 96438 91962
rect 96490 91910 96502 91962
rect 96554 91910 96566 91962
rect 96618 91910 96630 91962
rect 96682 91910 112914 91962
rect 112966 91910 112978 91962
rect 113030 91910 113042 91962
rect 113094 91910 113106 91962
rect 113158 91910 113170 91962
rect 113222 91910 118864 91962
rect 1104 91888 118864 91910
rect 49602 91808 49608 91860
rect 49660 91848 49666 91860
rect 55214 91848 55220 91860
rect 49660 91820 55220 91848
rect 49660 91808 49666 91820
rect 55214 91808 55220 91820
rect 55272 91808 55278 91860
rect 56042 91808 56048 91860
rect 56100 91848 56106 91860
rect 61746 91848 61752 91860
rect 56100 91820 61752 91848
rect 56100 91808 56106 91820
rect 61746 91808 61752 91820
rect 61804 91808 61810 91860
rect 77478 91740 77484 91792
rect 77536 91780 77542 91792
rect 108298 91780 108304 91792
rect 77536 91752 108304 91780
rect 77536 91740 77542 91752
rect 108298 91740 108304 91752
rect 108356 91740 108362 91792
rect 1104 91418 7912 91440
rect 1104 91366 4874 91418
rect 4926 91366 4938 91418
rect 4990 91366 5002 91418
rect 5054 91366 5066 91418
rect 5118 91366 5130 91418
rect 5182 91366 7912 91418
rect 1104 91344 7912 91366
rect 108008 91418 118864 91440
rect 108008 91366 113650 91418
rect 113702 91366 113714 91418
rect 113766 91366 113778 91418
rect 113830 91366 113842 91418
rect 113894 91366 113906 91418
rect 113958 91366 118864 91418
rect 108008 91344 118864 91366
rect 1104 90874 7912 90896
rect 1104 90822 4214 90874
rect 4266 90822 4278 90874
rect 4330 90822 4342 90874
rect 4394 90822 4406 90874
rect 4458 90822 4470 90874
rect 4522 90822 7912 90874
rect 1104 90800 7912 90822
rect 108008 90874 118864 90896
rect 108008 90822 112914 90874
rect 112966 90822 112978 90874
rect 113030 90822 113042 90874
rect 113094 90822 113106 90874
rect 113158 90822 113170 90874
rect 113222 90822 118864 90874
rect 108008 90800 118864 90822
rect 71130 90380 71136 90432
rect 71188 90420 71194 90432
rect 108390 90420 108396 90432
rect 71188 90392 108396 90420
rect 71188 90380 71194 90392
rect 108390 90380 108396 90392
rect 108448 90380 108454 90432
rect 1104 90330 7912 90352
rect 1104 90278 4874 90330
rect 4926 90278 4938 90330
rect 4990 90278 5002 90330
rect 5054 90278 5066 90330
rect 5118 90278 5130 90330
rect 5182 90278 7912 90330
rect 1104 90256 7912 90278
rect 108008 90330 118864 90352
rect 108008 90278 113650 90330
rect 113702 90278 113714 90330
rect 113766 90278 113778 90330
rect 113830 90278 113842 90330
rect 113894 90278 113906 90330
rect 113958 90278 118864 90330
rect 108008 90256 118864 90278
rect 1104 89786 7912 89808
rect 1104 89734 4214 89786
rect 4266 89734 4278 89786
rect 4330 89734 4342 89786
rect 4394 89734 4406 89786
rect 4458 89734 4470 89786
rect 4522 89734 7912 89786
rect 1104 89712 7912 89734
rect 108008 89786 118864 89808
rect 108008 89734 112914 89786
rect 112966 89734 112978 89786
rect 113030 89734 113042 89786
rect 113094 89734 113106 89786
rect 113158 89734 113170 89786
rect 113222 89734 118864 89786
rect 108008 89712 118864 89734
rect 1104 89242 7912 89264
rect 1104 89190 4874 89242
rect 4926 89190 4938 89242
rect 4990 89190 5002 89242
rect 5054 89190 5066 89242
rect 5118 89190 5130 89242
rect 5182 89190 7912 89242
rect 1104 89168 7912 89190
rect 108008 89242 118864 89264
rect 108008 89190 113650 89242
rect 113702 89190 113714 89242
rect 113766 89190 113778 89242
rect 113830 89190 113842 89242
rect 113894 89190 113906 89242
rect 113958 89190 118864 89242
rect 108008 89168 118864 89190
rect 1104 88698 7912 88720
rect 1104 88646 4214 88698
rect 4266 88646 4278 88698
rect 4330 88646 4342 88698
rect 4394 88646 4406 88698
rect 4458 88646 4470 88698
rect 4522 88646 7912 88698
rect 1104 88624 7912 88646
rect 108008 88698 118864 88720
rect 108008 88646 112914 88698
rect 112966 88646 112978 88698
rect 113030 88646 113042 88698
rect 113094 88646 113106 88698
rect 113158 88646 113170 88698
rect 113222 88646 118864 88698
rect 108008 88624 118864 88646
rect 1104 88154 7912 88176
rect 1104 88102 4874 88154
rect 4926 88102 4938 88154
rect 4990 88102 5002 88154
rect 5054 88102 5066 88154
rect 5118 88102 5130 88154
rect 5182 88102 7912 88154
rect 1104 88080 7912 88102
rect 108008 88154 118864 88176
rect 108008 88102 113650 88154
rect 113702 88102 113714 88154
rect 113766 88102 113778 88154
rect 113830 88102 113842 88154
rect 113894 88102 113906 88154
rect 113958 88102 118864 88154
rect 108008 88080 118864 88102
rect 1104 87610 7912 87632
rect 1104 87558 4214 87610
rect 4266 87558 4278 87610
rect 4330 87558 4342 87610
rect 4394 87558 4406 87610
rect 4458 87558 4470 87610
rect 4522 87558 7912 87610
rect 1104 87536 7912 87558
rect 108008 87610 118864 87632
rect 108008 87558 112914 87610
rect 112966 87558 112978 87610
rect 113030 87558 113042 87610
rect 113094 87558 113106 87610
rect 113158 87558 113170 87610
rect 113222 87558 118864 87610
rect 108008 87536 118864 87558
rect 1104 87066 7912 87088
rect 1104 87014 4874 87066
rect 4926 87014 4938 87066
rect 4990 87014 5002 87066
rect 5054 87014 5066 87066
rect 5118 87014 5130 87066
rect 5182 87014 7912 87066
rect 1104 86992 7912 87014
rect 108008 87066 118864 87088
rect 108008 87014 113650 87066
rect 113702 87014 113714 87066
rect 113766 87014 113778 87066
rect 113830 87014 113842 87066
rect 113894 87014 113906 87066
rect 113958 87014 118864 87066
rect 108008 86992 118864 87014
rect 106182 86572 106188 86624
rect 106240 86612 106246 86624
rect 108301 86615 108359 86621
rect 108301 86612 108313 86615
rect 106240 86584 108313 86612
rect 106240 86572 106246 86584
rect 108301 86581 108313 86584
rect 108347 86581 108359 86615
rect 108301 86575 108359 86581
rect 1104 86522 7912 86544
rect 1104 86470 4214 86522
rect 4266 86470 4278 86522
rect 4330 86470 4342 86522
rect 4394 86470 4406 86522
rect 4458 86470 4470 86522
rect 4522 86470 7912 86522
rect 1104 86448 7912 86470
rect 108008 86522 118864 86544
rect 108008 86470 112914 86522
rect 112966 86470 112978 86522
rect 113030 86470 113042 86522
rect 113094 86470 113106 86522
rect 113158 86470 113170 86522
rect 113222 86470 118864 86522
rect 108008 86448 118864 86470
rect 1104 85978 7912 86000
rect 1104 85926 4874 85978
rect 4926 85926 4938 85978
rect 4990 85926 5002 85978
rect 5054 85926 5066 85978
rect 5118 85926 5130 85978
rect 5182 85926 7912 85978
rect 1104 85904 7912 85926
rect 108008 85978 118864 86000
rect 108008 85926 113650 85978
rect 113702 85926 113714 85978
rect 113766 85926 113778 85978
rect 113830 85926 113842 85978
rect 113894 85926 113906 85978
rect 113958 85926 118864 85978
rect 108008 85904 118864 85926
rect 1104 85434 7912 85456
rect 1104 85382 4214 85434
rect 4266 85382 4278 85434
rect 4330 85382 4342 85434
rect 4394 85382 4406 85434
rect 4458 85382 4470 85434
rect 4522 85382 7912 85434
rect 1104 85360 7912 85382
rect 108008 85434 118864 85456
rect 108008 85382 112914 85434
rect 112966 85382 112978 85434
rect 113030 85382 113042 85434
rect 113094 85382 113106 85434
rect 113158 85382 113170 85434
rect 113222 85382 118864 85434
rect 108008 85360 118864 85382
rect 1104 84890 7912 84912
rect 1104 84838 4874 84890
rect 4926 84838 4938 84890
rect 4990 84838 5002 84890
rect 5054 84838 5066 84890
rect 5118 84838 5130 84890
rect 5182 84838 7912 84890
rect 1104 84816 7912 84838
rect 108008 84890 118864 84912
rect 108008 84838 113650 84890
rect 113702 84838 113714 84890
rect 113766 84838 113778 84890
rect 113830 84838 113842 84890
rect 113894 84838 113906 84890
rect 113958 84838 118864 84890
rect 108008 84816 118864 84838
rect 1104 84346 7912 84368
rect 1104 84294 4214 84346
rect 4266 84294 4278 84346
rect 4330 84294 4342 84346
rect 4394 84294 4406 84346
rect 4458 84294 4470 84346
rect 4522 84294 7912 84346
rect 1104 84272 7912 84294
rect 108008 84346 118864 84368
rect 108008 84294 112914 84346
rect 112966 84294 112978 84346
rect 113030 84294 113042 84346
rect 113094 84294 113106 84346
rect 113158 84294 113170 84346
rect 113222 84294 118864 84346
rect 108008 84272 118864 84294
rect 1104 83802 7912 83824
rect 1104 83750 4874 83802
rect 4926 83750 4938 83802
rect 4990 83750 5002 83802
rect 5054 83750 5066 83802
rect 5118 83750 5130 83802
rect 5182 83750 7912 83802
rect 1104 83728 7912 83750
rect 108008 83802 118864 83824
rect 108008 83750 113650 83802
rect 113702 83750 113714 83802
rect 113766 83750 113778 83802
rect 113830 83750 113842 83802
rect 113894 83750 113906 83802
rect 113958 83750 118864 83802
rect 108008 83728 118864 83750
rect 1104 83258 7912 83280
rect 1104 83206 4214 83258
rect 4266 83206 4278 83258
rect 4330 83206 4342 83258
rect 4394 83206 4406 83258
rect 4458 83206 4470 83258
rect 4522 83206 7912 83258
rect 1104 83184 7912 83206
rect 108008 83258 118864 83280
rect 108008 83206 112914 83258
rect 112966 83206 112978 83258
rect 113030 83206 113042 83258
rect 113094 83206 113106 83258
rect 113158 83206 113170 83258
rect 113222 83206 118864 83258
rect 108008 83184 118864 83206
rect 1104 82714 7912 82736
rect 1104 82662 4874 82714
rect 4926 82662 4938 82714
rect 4990 82662 5002 82714
rect 5054 82662 5066 82714
rect 5118 82662 5130 82714
rect 5182 82662 7912 82714
rect 1104 82640 7912 82662
rect 108008 82714 118864 82736
rect 108008 82662 113650 82714
rect 113702 82662 113714 82714
rect 113766 82662 113778 82714
rect 113830 82662 113842 82714
rect 113894 82662 113906 82714
rect 113958 82662 118864 82714
rect 108008 82640 118864 82662
rect 1104 82170 7912 82192
rect 1104 82118 4214 82170
rect 4266 82118 4278 82170
rect 4330 82118 4342 82170
rect 4394 82118 4406 82170
rect 4458 82118 4470 82170
rect 4522 82118 7912 82170
rect 1104 82096 7912 82118
rect 108008 82170 118864 82192
rect 108008 82118 112914 82170
rect 112966 82118 112978 82170
rect 113030 82118 113042 82170
rect 113094 82118 113106 82170
rect 113158 82118 113170 82170
rect 113222 82118 118864 82170
rect 108008 82096 118864 82118
rect 1104 81626 7912 81648
rect 1104 81574 4874 81626
rect 4926 81574 4938 81626
rect 4990 81574 5002 81626
rect 5054 81574 5066 81626
rect 5118 81574 5130 81626
rect 5182 81574 7912 81626
rect 1104 81552 7912 81574
rect 108008 81626 118864 81648
rect 108008 81574 113650 81626
rect 113702 81574 113714 81626
rect 113766 81574 113778 81626
rect 113830 81574 113842 81626
rect 113894 81574 113906 81626
rect 113958 81574 118864 81626
rect 108008 81552 118864 81574
rect 1104 81082 7912 81104
rect 1104 81030 4214 81082
rect 4266 81030 4278 81082
rect 4330 81030 4342 81082
rect 4394 81030 4406 81082
rect 4458 81030 4470 81082
rect 4522 81030 7912 81082
rect 1104 81008 7912 81030
rect 108008 81082 118864 81104
rect 108008 81030 112914 81082
rect 112966 81030 112978 81082
rect 113030 81030 113042 81082
rect 113094 81030 113106 81082
rect 113158 81030 113170 81082
rect 113222 81030 118864 81082
rect 108008 81008 118864 81030
rect 1104 80538 7912 80560
rect 1104 80486 4874 80538
rect 4926 80486 4938 80538
rect 4990 80486 5002 80538
rect 5054 80486 5066 80538
rect 5118 80486 5130 80538
rect 5182 80486 7912 80538
rect 1104 80464 7912 80486
rect 108008 80538 118864 80560
rect 108008 80486 113650 80538
rect 113702 80486 113714 80538
rect 113766 80486 113778 80538
rect 113830 80486 113842 80538
rect 113894 80486 113906 80538
rect 113958 80486 118864 80538
rect 108008 80464 118864 80486
rect 1104 79994 7912 80016
rect 1104 79942 4214 79994
rect 4266 79942 4278 79994
rect 4330 79942 4342 79994
rect 4394 79942 4406 79994
rect 4458 79942 4470 79994
rect 4522 79942 7912 79994
rect 1104 79920 7912 79942
rect 108008 79994 118864 80016
rect 108008 79942 112914 79994
rect 112966 79942 112978 79994
rect 113030 79942 113042 79994
rect 113094 79942 113106 79994
rect 113158 79942 113170 79994
rect 113222 79942 118864 79994
rect 108008 79920 118864 79942
rect 1104 79450 7912 79472
rect 1104 79398 4874 79450
rect 4926 79398 4938 79450
rect 4990 79398 5002 79450
rect 5054 79398 5066 79450
rect 5118 79398 5130 79450
rect 5182 79398 7912 79450
rect 1104 79376 7912 79398
rect 108008 79450 118864 79472
rect 108008 79398 113650 79450
rect 113702 79398 113714 79450
rect 113766 79398 113778 79450
rect 113830 79398 113842 79450
rect 113894 79398 113906 79450
rect 113958 79398 118864 79450
rect 108008 79376 118864 79398
rect 1104 78906 7912 78928
rect 1104 78854 4214 78906
rect 4266 78854 4278 78906
rect 4330 78854 4342 78906
rect 4394 78854 4406 78906
rect 4458 78854 4470 78906
rect 4522 78854 7912 78906
rect 1104 78832 7912 78854
rect 108008 78906 118864 78928
rect 108008 78854 112914 78906
rect 112966 78854 112978 78906
rect 113030 78854 113042 78906
rect 113094 78854 113106 78906
rect 113158 78854 113170 78906
rect 113222 78854 118864 78906
rect 108008 78832 118864 78854
rect 1104 78362 7912 78384
rect 1104 78310 4874 78362
rect 4926 78310 4938 78362
rect 4990 78310 5002 78362
rect 5054 78310 5066 78362
rect 5118 78310 5130 78362
rect 5182 78310 7912 78362
rect 1104 78288 7912 78310
rect 108008 78362 118864 78384
rect 108008 78310 113650 78362
rect 113702 78310 113714 78362
rect 113766 78310 113778 78362
rect 113830 78310 113842 78362
rect 113894 78310 113906 78362
rect 113958 78310 118864 78362
rect 108008 78288 118864 78310
rect 1104 77818 7912 77840
rect 1104 77766 4214 77818
rect 4266 77766 4278 77818
rect 4330 77766 4342 77818
rect 4394 77766 4406 77818
rect 4458 77766 4470 77818
rect 4522 77766 7912 77818
rect 1104 77744 7912 77766
rect 108008 77818 118864 77840
rect 108008 77766 112914 77818
rect 112966 77766 112978 77818
rect 113030 77766 113042 77818
rect 113094 77766 113106 77818
rect 113158 77766 113170 77818
rect 113222 77766 118864 77818
rect 108008 77744 118864 77766
rect 1104 77274 7912 77296
rect 1104 77222 4874 77274
rect 4926 77222 4938 77274
rect 4990 77222 5002 77274
rect 5054 77222 5066 77274
rect 5118 77222 5130 77274
rect 5182 77222 7912 77274
rect 1104 77200 7912 77222
rect 108008 77274 118864 77296
rect 108008 77222 113650 77274
rect 113702 77222 113714 77274
rect 113766 77222 113778 77274
rect 113830 77222 113842 77274
rect 113894 77222 113906 77274
rect 113958 77222 118864 77274
rect 108008 77200 118864 77222
rect 1104 76730 7912 76752
rect 1104 76678 4214 76730
rect 4266 76678 4278 76730
rect 4330 76678 4342 76730
rect 4394 76678 4406 76730
rect 4458 76678 4470 76730
rect 4522 76678 7912 76730
rect 1104 76656 7912 76678
rect 108008 76730 118864 76752
rect 108008 76678 112914 76730
rect 112966 76678 112978 76730
rect 113030 76678 113042 76730
rect 113094 76678 113106 76730
rect 113158 76678 113170 76730
rect 113222 76678 118864 76730
rect 108008 76656 118864 76678
rect 1104 76186 7912 76208
rect 1104 76134 4874 76186
rect 4926 76134 4938 76186
rect 4990 76134 5002 76186
rect 5054 76134 5066 76186
rect 5118 76134 5130 76186
rect 5182 76134 7912 76186
rect 1104 76112 7912 76134
rect 108008 76186 118864 76208
rect 108008 76134 113650 76186
rect 113702 76134 113714 76186
rect 113766 76134 113778 76186
rect 113830 76134 113842 76186
rect 113894 76134 113906 76186
rect 113958 76134 118864 76186
rect 108008 76112 118864 76134
rect 1104 75642 7912 75664
rect 1104 75590 4214 75642
rect 4266 75590 4278 75642
rect 4330 75590 4342 75642
rect 4394 75590 4406 75642
rect 4458 75590 4470 75642
rect 4522 75590 7912 75642
rect 1104 75568 7912 75590
rect 108008 75642 118864 75664
rect 108008 75590 112914 75642
rect 112966 75590 112978 75642
rect 113030 75590 113042 75642
rect 113094 75590 113106 75642
rect 113158 75590 113170 75642
rect 113222 75590 118864 75642
rect 108008 75568 118864 75590
rect 1104 75098 7912 75120
rect 1104 75046 4874 75098
rect 4926 75046 4938 75098
rect 4990 75046 5002 75098
rect 5054 75046 5066 75098
rect 5118 75046 5130 75098
rect 5182 75046 7912 75098
rect 1104 75024 7912 75046
rect 108008 75098 118864 75120
rect 108008 75046 113650 75098
rect 113702 75046 113714 75098
rect 113766 75046 113778 75098
rect 113830 75046 113842 75098
rect 113894 75046 113906 75098
rect 113958 75046 118864 75098
rect 108008 75024 118864 75046
rect 1104 74554 7912 74576
rect 1104 74502 4214 74554
rect 4266 74502 4278 74554
rect 4330 74502 4342 74554
rect 4394 74502 4406 74554
rect 4458 74502 4470 74554
rect 4522 74502 7912 74554
rect 1104 74480 7912 74502
rect 108008 74554 118864 74576
rect 108008 74502 112914 74554
rect 112966 74502 112978 74554
rect 113030 74502 113042 74554
rect 113094 74502 113106 74554
rect 113158 74502 113170 74554
rect 113222 74502 118864 74554
rect 108008 74480 118864 74502
rect 1104 74010 7912 74032
rect 1104 73958 4874 74010
rect 4926 73958 4938 74010
rect 4990 73958 5002 74010
rect 5054 73958 5066 74010
rect 5118 73958 5130 74010
rect 5182 73958 7912 74010
rect 1104 73936 7912 73958
rect 108008 74010 118864 74032
rect 108008 73958 113650 74010
rect 113702 73958 113714 74010
rect 113766 73958 113778 74010
rect 113830 73958 113842 74010
rect 113894 73958 113906 74010
rect 113958 73958 118864 74010
rect 108008 73936 118864 73958
rect 1104 73466 7912 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 7912 73466
rect 1104 73392 7912 73414
rect 108008 73466 118864 73488
rect 108008 73414 112914 73466
rect 112966 73414 112978 73466
rect 113030 73414 113042 73466
rect 113094 73414 113106 73466
rect 113158 73414 113170 73466
rect 113222 73414 118864 73466
rect 108008 73392 118864 73414
rect 1104 72922 7912 72944
rect 1104 72870 4874 72922
rect 4926 72870 4938 72922
rect 4990 72870 5002 72922
rect 5054 72870 5066 72922
rect 5118 72870 5130 72922
rect 5182 72870 7912 72922
rect 1104 72848 7912 72870
rect 108008 72922 118864 72944
rect 108008 72870 113650 72922
rect 113702 72870 113714 72922
rect 113766 72870 113778 72922
rect 113830 72870 113842 72922
rect 113894 72870 113906 72922
rect 113958 72870 118864 72922
rect 108008 72848 118864 72870
rect 1104 72378 7912 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 7912 72378
rect 1104 72304 7912 72326
rect 108008 72378 118864 72400
rect 108008 72326 112914 72378
rect 112966 72326 112978 72378
rect 113030 72326 113042 72378
rect 113094 72326 113106 72378
rect 113158 72326 113170 72378
rect 113222 72326 118864 72378
rect 108008 72304 118864 72326
rect 1104 71834 7912 71856
rect 1104 71782 4874 71834
rect 4926 71782 4938 71834
rect 4990 71782 5002 71834
rect 5054 71782 5066 71834
rect 5118 71782 5130 71834
rect 5182 71782 7912 71834
rect 1104 71760 7912 71782
rect 108008 71834 118864 71856
rect 108008 71782 113650 71834
rect 113702 71782 113714 71834
rect 113766 71782 113778 71834
rect 113830 71782 113842 71834
rect 113894 71782 113906 71834
rect 113958 71782 118864 71834
rect 108008 71760 118864 71782
rect 1104 71290 7912 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 7912 71290
rect 1104 71216 7912 71238
rect 108008 71290 118864 71312
rect 108008 71238 112914 71290
rect 112966 71238 112978 71290
rect 113030 71238 113042 71290
rect 113094 71238 113106 71290
rect 113158 71238 113170 71290
rect 113222 71238 118864 71290
rect 108008 71216 118864 71238
rect 1104 70746 7912 70768
rect 1104 70694 4874 70746
rect 4926 70694 4938 70746
rect 4990 70694 5002 70746
rect 5054 70694 5066 70746
rect 5118 70694 5130 70746
rect 5182 70694 7912 70746
rect 1104 70672 7912 70694
rect 108008 70746 118864 70768
rect 108008 70694 113650 70746
rect 113702 70694 113714 70746
rect 113766 70694 113778 70746
rect 113830 70694 113842 70746
rect 113894 70694 113906 70746
rect 113958 70694 118864 70746
rect 108008 70672 118864 70694
rect 1104 70202 7912 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 7912 70202
rect 1104 70128 7912 70150
rect 108008 70202 118864 70224
rect 108008 70150 112914 70202
rect 112966 70150 112978 70202
rect 113030 70150 113042 70202
rect 113094 70150 113106 70202
rect 113158 70150 113170 70202
rect 113222 70150 118864 70202
rect 108008 70128 118864 70150
rect 1104 69658 7912 69680
rect 1104 69606 4874 69658
rect 4926 69606 4938 69658
rect 4990 69606 5002 69658
rect 5054 69606 5066 69658
rect 5118 69606 5130 69658
rect 5182 69606 7912 69658
rect 1104 69584 7912 69606
rect 108008 69658 118864 69680
rect 108008 69606 113650 69658
rect 113702 69606 113714 69658
rect 113766 69606 113778 69658
rect 113830 69606 113842 69658
rect 113894 69606 113906 69658
rect 113958 69606 118864 69658
rect 108008 69584 118864 69606
rect 1104 69114 7912 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 7912 69114
rect 1104 69040 7912 69062
rect 108008 69114 118864 69136
rect 108008 69062 112914 69114
rect 112966 69062 112978 69114
rect 113030 69062 113042 69114
rect 113094 69062 113106 69114
rect 113158 69062 113170 69114
rect 113222 69062 118864 69114
rect 108008 69040 118864 69062
rect 1104 68570 7912 68592
rect 1104 68518 4874 68570
rect 4926 68518 4938 68570
rect 4990 68518 5002 68570
rect 5054 68518 5066 68570
rect 5118 68518 5130 68570
rect 5182 68518 7912 68570
rect 1104 68496 7912 68518
rect 108008 68570 118864 68592
rect 108008 68518 113650 68570
rect 113702 68518 113714 68570
rect 113766 68518 113778 68570
rect 113830 68518 113842 68570
rect 113894 68518 113906 68570
rect 113958 68518 118864 68570
rect 108008 68496 118864 68518
rect 1104 68026 7912 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 7912 68026
rect 1104 67952 7912 67974
rect 108008 68026 118864 68048
rect 108008 67974 112914 68026
rect 112966 67974 112978 68026
rect 113030 67974 113042 68026
rect 113094 67974 113106 68026
rect 113158 67974 113170 68026
rect 113222 67974 118864 68026
rect 108008 67952 118864 67974
rect 1104 67482 7912 67504
rect 1104 67430 4874 67482
rect 4926 67430 4938 67482
rect 4990 67430 5002 67482
rect 5054 67430 5066 67482
rect 5118 67430 5130 67482
rect 5182 67430 7912 67482
rect 1104 67408 7912 67430
rect 108008 67482 118864 67504
rect 108008 67430 113650 67482
rect 113702 67430 113714 67482
rect 113766 67430 113778 67482
rect 113830 67430 113842 67482
rect 113894 67430 113906 67482
rect 113958 67430 118864 67482
rect 108008 67408 118864 67430
rect 108390 67328 108396 67380
rect 108448 67368 108454 67380
rect 109865 67371 109923 67377
rect 109865 67368 109877 67371
rect 108448 67340 109877 67368
rect 108448 67328 108454 67340
rect 109865 67337 109877 67340
rect 109911 67337 109923 67371
rect 109865 67331 109923 67337
rect 109517 67235 109575 67241
rect 109517 67201 109529 67235
rect 109563 67232 109575 67235
rect 109678 67232 109684 67244
rect 109563 67204 109684 67232
rect 109563 67201 109575 67204
rect 109517 67195 109575 67201
rect 109678 67192 109684 67204
rect 109736 67192 109742 67244
rect 109773 67167 109831 67173
rect 109773 67133 109785 67167
rect 109819 67164 109831 67167
rect 109819 67136 110000 67164
rect 109819 67133 109831 67136
rect 109773 67127 109831 67133
rect 109972 67040 110000 67136
rect 109954 66988 109960 67040
rect 110012 67028 110018 67040
rect 110049 67031 110107 67037
rect 110049 67028 110061 67031
rect 110012 67000 110061 67028
rect 110012 66988 110018 67000
rect 110049 66997 110061 67000
rect 110095 66997 110107 67031
rect 110049 66991 110107 66997
rect 1104 66938 7912 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 7912 66938
rect 1104 66864 7912 66886
rect 108008 66938 118864 66960
rect 108008 66886 112914 66938
rect 112966 66886 112978 66938
rect 113030 66886 113042 66938
rect 113094 66886 113106 66938
rect 113158 66886 113170 66938
rect 113222 66886 118864 66938
rect 108008 66864 118864 66886
rect 1104 66394 7912 66416
rect 1104 66342 4874 66394
rect 4926 66342 4938 66394
rect 4990 66342 5002 66394
rect 5054 66342 5066 66394
rect 5118 66342 5130 66394
rect 5182 66342 7912 66394
rect 1104 66320 7912 66342
rect 108008 66394 118864 66416
rect 108008 66342 113650 66394
rect 113702 66342 113714 66394
rect 113766 66342 113778 66394
rect 113830 66342 113842 66394
rect 113894 66342 113906 66394
rect 113958 66342 118864 66394
rect 108008 66320 118864 66342
rect 1104 65850 7912 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 7912 65850
rect 1104 65776 7912 65798
rect 108008 65850 118864 65872
rect 108008 65798 112914 65850
rect 112966 65798 112978 65850
rect 113030 65798 113042 65850
rect 113094 65798 113106 65850
rect 113158 65798 113170 65850
rect 113222 65798 118864 65850
rect 108008 65776 118864 65798
rect 1104 65306 7912 65328
rect 1104 65254 4874 65306
rect 4926 65254 4938 65306
rect 4990 65254 5002 65306
rect 5054 65254 5066 65306
rect 5118 65254 5130 65306
rect 5182 65254 7912 65306
rect 1104 65232 7912 65254
rect 108008 65306 118864 65328
rect 108008 65254 113650 65306
rect 113702 65254 113714 65306
rect 113766 65254 113778 65306
rect 113830 65254 113842 65306
rect 113894 65254 113906 65306
rect 113958 65254 118864 65306
rect 108008 65232 118864 65254
rect 1104 64762 7912 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 7912 64762
rect 1104 64688 7912 64710
rect 108008 64762 118864 64784
rect 108008 64710 112914 64762
rect 112966 64710 112978 64762
rect 113030 64710 113042 64762
rect 113094 64710 113106 64762
rect 113158 64710 113170 64762
rect 113222 64710 118864 64762
rect 108008 64688 118864 64710
rect 1104 64218 7912 64240
rect 1104 64166 4874 64218
rect 4926 64166 4938 64218
rect 4990 64166 5002 64218
rect 5054 64166 5066 64218
rect 5118 64166 5130 64218
rect 5182 64166 7912 64218
rect 1104 64144 7912 64166
rect 108008 64218 118864 64240
rect 108008 64166 113650 64218
rect 113702 64166 113714 64218
rect 113766 64166 113778 64218
rect 113830 64166 113842 64218
rect 113894 64166 113906 64218
rect 113958 64166 118864 64218
rect 108008 64144 118864 64166
rect 1104 63674 7912 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 7912 63674
rect 1104 63600 7912 63622
rect 108008 63674 118864 63696
rect 108008 63622 112914 63674
rect 112966 63622 112978 63674
rect 113030 63622 113042 63674
rect 113094 63622 113106 63674
rect 113158 63622 113170 63674
rect 113222 63622 118864 63674
rect 108008 63600 118864 63622
rect 1104 63130 7912 63152
rect 1104 63078 4874 63130
rect 4926 63078 4938 63130
rect 4990 63078 5002 63130
rect 5054 63078 5066 63130
rect 5118 63078 5130 63130
rect 5182 63078 7912 63130
rect 1104 63056 7912 63078
rect 108008 63130 118864 63152
rect 108008 63078 113650 63130
rect 113702 63078 113714 63130
rect 113766 63078 113778 63130
rect 113830 63078 113842 63130
rect 113894 63078 113906 63130
rect 113958 63078 118864 63130
rect 108008 63056 118864 63078
rect 1104 62586 7912 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 7912 62586
rect 1104 62512 7912 62534
rect 108008 62586 118864 62608
rect 108008 62534 112914 62586
rect 112966 62534 112978 62586
rect 113030 62534 113042 62586
rect 113094 62534 113106 62586
rect 113158 62534 113170 62586
rect 113222 62534 118864 62586
rect 108008 62512 118864 62534
rect 1104 62042 7912 62064
rect 1104 61990 4874 62042
rect 4926 61990 4938 62042
rect 4990 61990 5002 62042
rect 5054 61990 5066 62042
rect 5118 61990 5130 62042
rect 5182 61990 7912 62042
rect 1104 61968 7912 61990
rect 108008 62042 118864 62064
rect 108008 61990 113650 62042
rect 113702 61990 113714 62042
rect 113766 61990 113778 62042
rect 113830 61990 113842 62042
rect 113894 61990 113906 62042
rect 113958 61990 118864 62042
rect 108008 61968 118864 61990
rect 1104 61498 7912 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 7912 61498
rect 1104 61424 7912 61446
rect 108008 61498 118864 61520
rect 108008 61446 112914 61498
rect 112966 61446 112978 61498
rect 113030 61446 113042 61498
rect 113094 61446 113106 61498
rect 113158 61446 113170 61498
rect 113222 61446 118864 61498
rect 108008 61424 118864 61446
rect 1104 60954 7912 60976
rect 1104 60902 4874 60954
rect 4926 60902 4938 60954
rect 4990 60902 5002 60954
rect 5054 60902 5066 60954
rect 5118 60902 5130 60954
rect 5182 60902 7912 60954
rect 1104 60880 7912 60902
rect 108008 60954 118864 60976
rect 108008 60902 113650 60954
rect 113702 60902 113714 60954
rect 113766 60902 113778 60954
rect 113830 60902 113842 60954
rect 113894 60902 113906 60954
rect 113958 60902 118864 60954
rect 108008 60880 118864 60902
rect 1104 60410 7912 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 7912 60410
rect 1104 60336 7912 60358
rect 108008 60410 118864 60432
rect 108008 60358 112914 60410
rect 112966 60358 112978 60410
rect 113030 60358 113042 60410
rect 113094 60358 113106 60410
rect 113158 60358 113170 60410
rect 113222 60358 118864 60410
rect 108008 60336 118864 60358
rect 1104 59866 7912 59888
rect 1104 59814 4874 59866
rect 4926 59814 4938 59866
rect 4990 59814 5002 59866
rect 5054 59814 5066 59866
rect 5118 59814 5130 59866
rect 5182 59814 7912 59866
rect 1104 59792 7912 59814
rect 108008 59866 118864 59888
rect 108008 59814 113650 59866
rect 113702 59814 113714 59866
rect 113766 59814 113778 59866
rect 113830 59814 113842 59866
rect 113894 59814 113906 59866
rect 113958 59814 118864 59866
rect 108008 59792 118864 59814
rect 1104 59322 7912 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 7912 59322
rect 1104 59248 7912 59270
rect 108008 59322 118864 59344
rect 108008 59270 112914 59322
rect 112966 59270 112978 59322
rect 113030 59270 113042 59322
rect 113094 59270 113106 59322
rect 113158 59270 113170 59322
rect 113222 59270 118864 59322
rect 108008 59248 118864 59270
rect 1104 58778 7912 58800
rect 1104 58726 4874 58778
rect 4926 58726 4938 58778
rect 4990 58726 5002 58778
rect 5054 58726 5066 58778
rect 5118 58726 5130 58778
rect 5182 58726 7912 58778
rect 1104 58704 7912 58726
rect 108008 58778 118864 58800
rect 108008 58726 113650 58778
rect 113702 58726 113714 58778
rect 113766 58726 113778 58778
rect 113830 58726 113842 58778
rect 113894 58726 113906 58778
rect 113958 58726 118864 58778
rect 108008 58704 118864 58726
rect 1104 58234 7912 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 7912 58234
rect 1104 58160 7912 58182
rect 108008 58234 118864 58256
rect 108008 58182 112914 58234
rect 112966 58182 112978 58234
rect 113030 58182 113042 58234
rect 113094 58182 113106 58234
rect 113158 58182 113170 58234
rect 113222 58182 118864 58234
rect 108008 58160 118864 58182
rect 108301 57919 108359 57925
rect 108301 57885 108313 57919
rect 108347 57916 108359 57919
rect 109954 57916 109960 57928
rect 108347 57888 109960 57916
rect 108347 57885 108359 57888
rect 108301 57879 108359 57885
rect 109954 57876 109960 57888
rect 110012 57876 110018 57928
rect 108568 57851 108626 57857
rect 108568 57817 108580 57851
rect 108614 57848 108626 57851
rect 108666 57848 108672 57860
rect 108614 57820 108672 57848
rect 108614 57817 108626 57820
rect 108568 57811 108626 57817
rect 108666 57808 108672 57820
rect 108724 57848 108730 57860
rect 109773 57851 109831 57857
rect 109773 57848 109785 57851
rect 108724 57820 109785 57848
rect 108724 57808 108730 57820
rect 109773 57817 109785 57820
rect 109819 57817 109831 57851
rect 109773 57811 109831 57817
rect 109678 57740 109684 57792
rect 109736 57740 109742 57792
rect 1104 57690 7912 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 7912 57690
rect 1104 57616 7912 57638
rect 108008 57690 118864 57712
rect 108008 57638 113650 57690
rect 113702 57638 113714 57690
rect 113766 57638 113778 57690
rect 113830 57638 113842 57690
rect 113894 57638 113906 57690
rect 113958 57638 118864 57690
rect 108008 57616 118864 57638
rect 1104 57146 7912 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 7912 57146
rect 1104 57072 7912 57094
rect 108008 57146 118864 57168
rect 108008 57094 112914 57146
rect 112966 57094 112978 57146
rect 113030 57094 113042 57146
rect 113094 57094 113106 57146
rect 113158 57094 113170 57146
rect 113222 57094 118864 57146
rect 108008 57072 118864 57094
rect 1104 56602 7912 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 7912 56602
rect 1104 56528 7912 56550
rect 108008 56602 118864 56624
rect 108008 56550 113650 56602
rect 113702 56550 113714 56602
rect 113766 56550 113778 56602
rect 113830 56550 113842 56602
rect 113894 56550 113906 56602
rect 113958 56550 118864 56602
rect 108008 56528 118864 56550
rect 1104 56058 7912 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 7912 56058
rect 1104 55984 7912 56006
rect 108008 56058 118864 56080
rect 108008 56006 112914 56058
rect 112966 56006 112978 56058
rect 113030 56006 113042 56058
rect 113094 56006 113106 56058
rect 113158 56006 113170 56058
rect 113222 56006 118864 56058
rect 108008 55984 118864 56006
rect 1104 55514 7912 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 7912 55514
rect 1104 55440 7912 55462
rect 108008 55514 118864 55536
rect 108008 55462 113650 55514
rect 113702 55462 113714 55514
rect 113766 55462 113778 55514
rect 113830 55462 113842 55514
rect 113894 55462 113906 55514
rect 113958 55462 118864 55514
rect 108008 55440 118864 55462
rect 1104 54970 7912 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 7912 54970
rect 1104 54896 7912 54918
rect 108008 54970 118864 54992
rect 108008 54918 112914 54970
rect 112966 54918 112978 54970
rect 113030 54918 113042 54970
rect 113094 54918 113106 54970
rect 113158 54918 113170 54970
rect 113222 54918 118864 54970
rect 108008 54896 118864 54918
rect 108574 54816 108580 54868
rect 108632 54816 108638 54868
rect 108301 54655 108359 54661
rect 108301 54621 108313 54655
rect 108347 54652 108359 54655
rect 108574 54652 108580 54664
rect 108347 54624 108580 54652
rect 108347 54621 108359 54624
rect 108301 54615 108359 54621
rect 108574 54612 108580 54624
rect 108632 54612 108638 54664
rect 108393 54587 108451 54593
rect 108393 54553 108405 54587
rect 108439 54584 108451 54587
rect 109126 54584 109132 54596
rect 108439 54556 109132 54584
rect 108439 54553 108451 54556
rect 108393 54547 108451 54553
rect 109126 54544 109132 54556
rect 109184 54544 109190 54596
rect 1104 54426 7912 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 7912 54426
rect 1104 54352 7912 54374
rect 108008 54426 118864 54448
rect 108008 54374 113650 54426
rect 113702 54374 113714 54426
rect 113766 54374 113778 54426
rect 113830 54374 113842 54426
rect 113894 54374 113906 54426
rect 113958 54374 118864 54426
rect 108008 54352 118864 54374
rect 108298 54272 108304 54324
rect 108356 54272 108362 54324
rect 1104 53882 7912 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 7912 53882
rect 1104 53808 7912 53830
rect 108008 53882 118864 53904
rect 108008 53830 112914 53882
rect 112966 53830 112978 53882
rect 113030 53830 113042 53882
rect 113094 53830 113106 53882
rect 113158 53830 113170 53882
rect 113222 53830 118864 53882
rect 108008 53808 118864 53830
rect 108298 53524 108304 53576
rect 108356 53524 108362 53576
rect 110049 53499 110107 53505
rect 110049 53465 110061 53499
rect 110095 53465 110107 53499
rect 110049 53459 110107 53465
rect 109034 53388 109040 53440
rect 109092 53428 109098 53440
rect 109954 53428 109960 53440
rect 109092 53400 109960 53428
rect 109092 53388 109098 53400
rect 109954 53388 109960 53400
rect 110012 53428 110018 53440
rect 110064 53428 110092 53459
rect 110233 53431 110291 53437
rect 110233 53428 110245 53431
rect 110012 53400 110245 53428
rect 110012 53388 110018 53400
rect 110233 53397 110245 53400
rect 110279 53428 110291 53431
rect 110690 53428 110696 53440
rect 110279 53400 110696 53428
rect 110279 53397 110291 53400
rect 110233 53391 110291 53397
rect 110690 53388 110696 53400
rect 110748 53388 110754 53440
rect 1104 53338 7912 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 7912 53338
rect 1104 53264 7912 53286
rect 108008 53338 118864 53360
rect 108008 53286 113650 53338
rect 113702 53286 113714 53338
rect 113766 53286 113778 53338
rect 113830 53286 113842 53338
rect 113894 53286 113906 53338
rect 113958 53286 118864 53338
rect 108008 53264 118864 53286
rect 109034 53184 109040 53236
rect 109092 53184 109098 53236
rect 108761 53091 108819 53097
rect 108761 53057 108773 53091
rect 108807 53088 108819 53091
rect 109052 53088 109080 53184
rect 108807 53060 109080 53088
rect 108807 53057 108819 53060
rect 108761 53051 108819 53057
rect 1104 52794 7912 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 7912 52794
rect 1104 52720 7912 52742
rect 108008 52794 118864 52816
rect 108008 52742 112914 52794
rect 112966 52742 112978 52794
rect 113030 52742 113042 52794
rect 113094 52742 113106 52794
rect 113158 52742 113170 52794
rect 113222 52742 118864 52794
rect 108008 52720 118864 52742
rect 108301 52547 108359 52553
rect 108301 52513 108313 52547
rect 108347 52544 108359 52547
rect 109034 52544 109040 52556
rect 108347 52516 109040 52544
rect 108347 52513 108359 52516
rect 108301 52507 108359 52513
rect 109034 52504 109040 52516
rect 109092 52504 109098 52556
rect 110509 52479 110567 52485
rect 110509 52445 110521 52479
rect 110555 52476 110567 52479
rect 110690 52476 110696 52488
rect 110555 52448 110696 52476
rect 110555 52445 110567 52448
rect 110509 52439 110567 52445
rect 110690 52436 110696 52448
rect 110748 52436 110754 52488
rect 108574 52368 108580 52420
rect 108632 52368 108638 52420
rect 109126 52368 109132 52420
rect 109184 52368 109190 52420
rect 110325 52411 110383 52417
rect 110325 52377 110337 52411
rect 110371 52377 110383 52411
rect 110325 52371 110383 52377
rect 109402 52300 109408 52352
rect 109460 52340 109466 52352
rect 110340 52340 110368 52371
rect 109460 52312 110368 52340
rect 109460 52300 109466 52312
rect 1104 52250 7912 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 7912 52250
rect 1104 52176 7912 52198
rect 108008 52250 118864 52272
rect 108008 52198 113650 52250
rect 113702 52198 113714 52250
rect 113766 52198 113778 52250
rect 113830 52198 113842 52250
rect 113894 52198 113906 52250
rect 113958 52198 118864 52250
rect 108008 52176 118864 52198
rect 108298 52096 108304 52148
rect 108356 52096 108362 52148
rect 106918 52028 106924 52080
rect 106976 52068 106982 52080
rect 109313 52071 109371 52077
rect 109313 52068 109325 52071
rect 106976 52040 109325 52068
rect 106976 52028 106982 52040
rect 109313 52037 109325 52040
rect 109359 52068 109371 52071
rect 109589 52071 109647 52077
rect 109589 52068 109601 52071
rect 109359 52040 109601 52068
rect 109359 52037 109371 52040
rect 109313 52031 109371 52037
rect 109589 52037 109601 52040
rect 109635 52037 109647 52071
rect 109589 52031 109647 52037
rect 109037 52003 109095 52009
rect 109037 51969 109049 52003
rect 109083 52000 109095 52003
rect 109402 52000 109408 52012
rect 109083 51972 109408 52000
rect 109083 51969 109095 51972
rect 109037 51963 109095 51969
rect 109402 51960 109408 51972
rect 109460 51960 109466 52012
rect 1104 51706 7912 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 7912 51706
rect 1104 51632 7912 51654
rect 108008 51706 118864 51728
rect 108008 51654 112914 51706
rect 112966 51654 112978 51706
rect 113030 51654 113042 51706
rect 113094 51654 113106 51706
rect 113158 51654 113170 51706
rect 113222 51654 118864 51706
rect 108008 51632 118864 51654
rect 108298 51348 108304 51400
rect 108356 51348 108362 51400
rect 109586 51212 109592 51264
rect 109644 51212 109650 51264
rect 1104 51162 7912 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 7912 51162
rect 1104 51088 7912 51110
rect 108008 51162 118864 51184
rect 108008 51110 113650 51162
rect 113702 51110 113714 51162
rect 113766 51110 113778 51162
rect 113830 51110 113842 51162
rect 113894 51110 113906 51162
rect 113958 51110 118864 51162
rect 108008 51088 118864 51110
rect 108761 50983 108819 50989
rect 108761 50949 108773 50983
rect 108807 50980 108819 50983
rect 109586 50980 109592 50992
rect 108807 50952 109592 50980
rect 108807 50949 108819 50952
rect 108761 50943 108819 50949
rect 109586 50940 109592 50952
rect 109644 50940 109650 50992
rect 108666 50872 108672 50924
rect 108724 50912 108730 50924
rect 108853 50915 108911 50921
rect 108853 50912 108865 50915
rect 108724 50884 108865 50912
rect 108724 50872 108730 50884
rect 108853 50881 108865 50884
rect 108899 50912 108911 50915
rect 109129 50915 109187 50921
rect 109129 50912 109141 50915
rect 108899 50884 109141 50912
rect 108899 50881 108911 50884
rect 108853 50875 108911 50881
rect 109129 50881 109141 50884
rect 109175 50881 109187 50915
rect 109129 50875 109187 50881
rect 108942 50668 108948 50720
rect 109000 50668 109006 50720
rect 1104 50618 7912 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 7912 50618
rect 1104 50544 7912 50566
rect 108008 50618 118864 50640
rect 108008 50566 112914 50618
rect 112966 50566 112978 50618
rect 113030 50566 113042 50618
rect 113094 50566 113106 50618
rect 113158 50566 113170 50618
rect 113222 50566 118864 50618
rect 108008 50544 118864 50566
rect 108666 50464 108672 50516
rect 108724 50464 108730 50516
rect 108301 50303 108359 50309
rect 108301 50269 108313 50303
rect 108347 50300 108359 50303
rect 108666 50300 108672 50312
rect 108347 50272 108672 50300
rect 108347 50269 108359 50272
rect 108301 50263 108359 50269
rect 108666 50260 108672 50272
rect 108724 50260 108730 50312
rect 108393 50235 108451 50241
rect 108393 50201 108405 50235
rect 108439 50232 108451 50235
rect 109126 50232 109132 50244
rect 108439 50204 109132 50232
rect 108439 50201 108451 50204
rect 108393 50195 108451 50201
rect 109126 50192 109132 50204
rect 109184 50192 109190 50244
rect 1104 50074 7912 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 7912 50074
rect 1104 50000 7912 50022
rect 108008 50074 118864 50096
rect 108008 50022 113650 50074
rect 113702 50022 113714 50074
rect 113766 50022 113778 50074
rect 113830 50022 113842 50074
rect 113894 50022 113906 50074
rect 113958 50022 118864 50074
rect 108008 50000 118864 50022
rect 1104 49530 7912 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 7912 49530
rect 1104 49456 7912 49478
rect 108008 49530 118864 49552
rect 108008 49478 112914 49530
rect 112966 49478 112978 49530
rect 113030 49478 113042 49530
rect 113094 49478 113106 49530
rect 113158 49478 113170 49530
rect 113222 49478 118864 49530
rect 108008 49456 118864 49478
rect 108574 49376 108580 49428
rect 108632 49416 108638 49428
rect 108945 49419 109003 49425
rect 108945 49416 108957 49419
rect 108632 49388 108957 49416
rect 108632 49376 108638 49388
rect 108945 49385 108957 49388
rect 108991 49385 109003 49419
rect 108945 49379 109003 49385
rect 108666 49308 108672 49360
rect 108724 49308 108730 49360
rect 109129 49351 109187 49357
rect 109129 49317 109141 49351
rect 109175 49348 109187 49351
rect 109494 49348 109500 49360
rect 109175 49320 109500 49348
rect 109175 49317 109187 49320
rect 109129 49311 109187 49317
rect 109494 49308 109500 49320
rect 109552 49308 109558 49360
rect 108298 49172 108304 49224
rect 108356 49212 108362 49224
rect 108684 49212 108712 49308
rect 108356 49184 108712 49212
rect 108356 49172 108362 49184
rect 108393 49147 108451 49153
rect 108393 49113 108405 49147
rect 108439 49144 108451 49147
rect 109034 49144 109040 49156
rect 108439 49116 109040 49144
rect 108439 49113 108451 49116
rect 108393 49107 108451 49113
rect 109034 49104 109040 49116
rect 109092 49104 109098 49156
rect 109402 49104 109408 49156
rect 109460 49104 109466 49156
rect 1104 48986 7912 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 7912 48986
rect 1104 48912 7912 48934
rect 108008 48986 118864 49008
rect 108008 48934 113650 48986
rect 113702 48934 113714 48986
rect 113766 48934 113778 48986
rect 113830 48934 113842 48986
rect 113894 48934 113906 48986
rect 113958 48934 118864 48986
rect 108008 48912 118864 48934
rect 1104 48442 7912 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 7912 48442
rect 1104 48368 7912 48390
rect 108008 48442 118864 48464
rect 108008 48390 112914 48442
rect 112966 48390 112978 48442
rect 113030 48390 113042 48442
rect 113094 48390 113106 48442
rect 113158 48390 113170 48442
rect 113222 48390 118864 48442
rect 108008 48368 118864 48390
rect 109586 48152 109592 48204
rect 109644 48192 109650 48204
rect 110322 48192 110328 48204
rect 109644 48164 110328 48192
rect 109644 48152 109650 48164
rect 110322 48152 110328 48164
rect 110380 48152 110386 48204
rect 108942 48084 108948 48136
rect 109000 48084 109006 48136
rect 110046 48016 110052 48068
rect 110104 48016 110110 48068
rect 108574 47948 108580 48000
rect 108632 47948 108638 48000
rect 1104 47898 7912 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 7912 47898
rect 1104 47824 7912 47846
rect 108008 47898 118864 47920
rect 108008 47846 113650 47898
rect 113702 47846 113714 47898
rect 113766 47846 113778 47898
rect 113830 47846 113842 47898
rect 113894 47846 113906 47898
rect 113958 47846 118864 47898
rect 108008 47824 118864 47846
rect 1104 47354 7912 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 7912 47354
rect 1104 47280 7912 47302
rect 108008 47354 118864 47376
rect 108008 47302 112914 47354
rect 112966 47302 112978 47354
rect 113030 47302 113042 47354
rect 113094 47302 113106 47354
rect 113158 47302 113170 47354
rect 113222 47302 118864 47354
rect 108008 47280 118864 47302
rect 108669 47243 108727 47249
rect 108669 47209 108681 47243
rect 108715 47240 108727 47243
rect 108758 47240 108764 47252
rect 108715 47212 108764 47240
rect 108715 47209 108727 47212
rect 108669 47203 108727 47209
rect 108758 47200 108764 47212
rect 108816 47240 108822 47252
rect 110506 47240 110512 47252
rect 108816 47212 110512 47240
rect 108816 47200 108822 47212
rect 110506 47200 110512 47212
rect 110564 47240 110570 47252
rect 110693 47243 110751 47249
rect 110693 47240 110705 47243
rect 110564 47212 110705 47240
rect 110564 47200 110570 47212
rect 110693 47209 110705 47212
rect 110739 47209 110751 47243
rect 110693 47203 110751 47209
rect 110414 47064 110420 47116
rect 110472 47064 110478 47116
rect 109126 46928 109132 46980
rect 109184 46928 109190 46980
rect 110138 46928 110144 46980
rect 110196 46928 110202 46980
rect 1104 46810 7912 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 7912 46810
rect 1104 46736 7912 46758
rect 108008 46810 118864 46832
rect 108008 46758 113650 46810
rect 113702 46758 113714 46810
rect 113766 46758 113778 46810
rect 113830 46758 113842 46810
rect 113894 46758 113906 46810
rect 113958 46758 118864 46810
rect 108008 46736 118864 46758
rect 108574 46520 108580 46572
rect 108632 46560 108638 46572
rect 109221 46563 109279 46569
rect 109221 46560 109233 46563
rect 108632 46532 109233 46560
rect 108632 46520 108638 46532
rect 109221 46529 109233 46532
rect 109267 46529 109279 46563
rect 109221 46523 109279 46529
rect 109678 46316 109684 46368
rect 109736 46316 109742 46368
rect 1104 46266 7912 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 7912 46266
rect 1104 46192 7912 46214
rect 108008 46266 118864 46288
rect 108008 46214 112914 46266
rect 112966 46214 112978 46266
rect 113030 46214 113042 46266
rect 113094 46214 113106 46266
rect 113158 46214 113170 46266
rect 113222 46214 118864 46266
rect 108008 46192 118864 46214
rect 110322 46112 110328 46164
rect 110380 46112 110386 46164
rect 110340 46016 110368 46112
rect 110417 46019 110475 46025
rect 110417 46016 110429 46019
rect 110340 45988 110429 46016
rect 110417 45985 110429 45988
rect 110463 45985 110475 46019
rect 110417 45979 110475 45985
rect 108298 45908 108304 45960
rect 108356 45908 108362 45960
rect 109034 45908 109040 45960
rect 109092 45908 109098 45960
rect 110141 45883 110199 45889
rect 110141 45849 110153 45883
rect 110187 45880 110199 45883
rect 110414 45880 110420 45892
rect 110187 45852 110420 45880
rect 110187 45849 110199 45852
rect 110141 45843 110199 45849
rect 110414 45840 110420 45852
rect 110472 45840 110478 45892
rect 108393 45815 108451 45821
rect 108393 45781 108405 45815
rect 108439 45812 108451 45815
rect 108482 45812 108488 45824
rect 108439 45784 108488 45812
rect 108439 45781 108451 45784
rect 108393 45775 108451 45781
rect 108482 45772 108488 45784
rect 108540 45772 108546 45824
rect 108669 45815 108727 45821
rect 108669 45781 108681 45815
rect 108715 45812 108727 45815
rect 109218 45812 109224 45824
rect 108715 45784 109224 45812
rect 108715 45781 108727 45784
rect 108669 45775 108727 45781
rect 109218 45772 109224 45784
rect 109276 45772 109282 45824
rect 1104 45722 7912 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 7912 45722
rect 1104 45648 7912 45670
rect 108008 45722 118864 45744
rect 108008 45670 113650 45722
rect 113702 45670 113714 45722
rect 113766 45670 113778 45722
rect 113830 45670 113842 45722
rect 113894 45670 113906 45722
rect 113958 45670 118864 45722
rect 108008 45648 118864 45670
rect 108298 45568 108304 45620
rect 108356 45568 108362 45620
rect 109205 45543 109263 45549
rect 109205 45509 109217 45543
rect 109251 45540 109263 45543
rect 109310 45540 109316 45552
rect 109251 45512 109316 45540
rect 109251 45509 109263 45512
rect 109205 45503 109263 45509
rect 109310 45500 109316 45512
rect 109368 45500 109374 45552
rect 109402 45500 109408 45552
rect 109460 45500 109466 45552
rect 109494 45500 109500 45552
rect 109552 45540 109558 45552
rect 110601 45543 110659 45549
rect 110601 45540 110613 45543
rect 109552 45512 110613 45540
rect 109552 45500 109558 45512
rect 110601 45509 110613 45512
rect 110647 45509 110659 45543
rect 110601 45503 110659 45509
rect 108574 45432 108580 45484
rect 108632 45472 108638 45484
rect 108761 45475 108819 45481
rect 108761 45472 108773 45475
rect 108632 45444 108773 45472
rect 108632 45432 108638 45444
rect 108761 45441 108773 45444
rect 108807 45441 108819 45475
rect 109420 45472 109448 45500
rect 109586 45472 109592 45484
rect 109420 45444 109592 45472
rect 108761 45435 108819 45441
rect 109586 45432 109592 45444
rect 109644 45432 109650 45484
rect 109678 45432 109684 45484
rect 109736 45472 109742 45484
rect 110325 45475 110383 45481
rect 110325 45472 110337 45475
rect 109736 45444 110337 45472
rect 109736 45432 109742 45444
rect 110325 45441 110337 45444
rect 110371 45472 110383 45475
rect 110417 45475 110475 45481
rect 110417 45472 110429 45475
rect 110371 45444 110429 45472
rect 110371 45441 110383 45444
rect 110325 45435 110383 45441
rect 110417 45441 110429 45444
rect 110463 45441 110475 45475
rect 110417 45435 110475 45441
rect 110046 45404 110052 45416
rect 109052 45376 110052 45404
rect 109052 45345 109080 45376
rect 110046 45364 110052 45376
rect 110104 45364 110110 45416
rect 109037 45339 109095 45345
rect 109037 45305 109049 45339
rect 109083 45305 109095 45339
rect 110785 45339 110843 45345
rect 110785 45336 110797 45339
rect 109037 45299 109095 45305
rect 109236 45308 110797 45336
rect 108945 45271 109003 45277
rect 108945 45237 108957 45271
rect 108991 45268 109003 45271
rect 109126 45268 109132 45280
rect 108991 45240 109132 45268
rect 108991 45237 109003 45240
rect 108945 45231 109003 45237
rect 109126 45228 109132 45240
rect 109184 45228 109190 45280
rect 109236 45277 109264 45308
rect 110785 45305 110797 45308
rect 110831 45305 110843 45339
rect 110785 45299 110843 45305
rect 109221 45271 109279 45277
rect 109221 45237 109233 45271
rect 109267 45237 109279 45271
rect 109221 45231 109279 45237
rect 109586 45228 109592 45280
rect 109644 45268 109650 45280
rect 109773 45271 109831 45277
rect 109773 45268 109785 45271
rect 109644 45240 109785 45268
rect 109644 45228 109650 45240
rect 109773 45237 109785 45240
rect 109819 45237 109831 45271
rect 109773 45231 109831 45237
rect 1104 45178 7912 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 7912 45178
rect 1104 45104 7912 45126
rect 108008 45178 118864 45200
rect 108008 45126 112914 45178
rect 112966 45126 112978 45178
rect 113030 45126 113042 45178
rect 113094 45126 113106 45178
rect 113158 45126 113170 45178
rect 113222 45126 118864 45178
rect 108008 45104 118864 45126
rect 109310 45024 109316 45076
rect 109368 45064 109374 45076
rect 109497 45067 109555 45073
rect 109497 45064 109509 45067
rect 109368 45036 109509 45064
rect 109368 45024 109374 45036
rect 109497 45033 109509 45036
rect 109543 45033 109555 45067
rect 109497 45027 109555 45033
rect 109405 44863 109463 44869
rect 109405 44829 109417 44863
rect 109451 44860 109463 44863
rect 109494 44860 109500 44872
rect 109451 44832 109500 44860
rect 109451 44829 109463 44832
rect 109405 44823 109463 44829
rect 109494 44820 109500 44832
rect 109552 44820 109558 44872
rect 109586 44820 109592 44872
rect 109644 44820 109650 44872
rect 1104 44634 7912 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 7912 44634
rect 1104 44560 7912 44582
rect 108008 44634 118864 44656
rect 108008 44582 113650 44634
rect 113702 44582 113714 44634
rect 113766 44582 113778 44634
rect 113830 44582 113842 44634
rect 113894 44582 113906 44634
rect 113958 44582 118864 44634
rect 108008 44560 118864 44582
rect 1302 44344 1308 44396
rect 1360 44384 1366 44396
rect 1397 44387 1455 44393
rect 1397 44384 1409 44387
rect 1360 44356 1409 44384
rect 1360 44344 1366 44356
rect 1397 44353 1409 44356
rect 1443 44384 1455 44387
rect 1673 44387 1731 44393
rect 1673 44384 1685 44387
rect 1443 44356 1685 44384
rect 1443 44353 1455 44356
rect 1397 44347 1455 44353
rect 1673 44353 1685 44356
rect 1719 44353 1731 44387
rect 1673 44347 1731 44353
rect 108298 44344 108304 44396
rect 108356 44384 108362 44396
rect 108577 44387 108635 44393
rect 108577 44384 108589 44387
rect 108356 44356 108589 44384
rect 108356 44344 108362 44356
rect 108577 44353 108589 44356
rect 108623 44353 108635 44387
rect 108577 44347 108635 44353
rect 1581 44251 1639 44257
rect 1581 44217 1593 44251
rect 1627 44248 1639 44251
rect 108393 44251 108451 44257
rect 1627 44220 6914 44248
rect 1627 44217 1639 44220
rect 1581 44211 1639 44217
rect 6886 44180 6914 44220
rect 108393 44217 108405 44251
rect 108439 44248 108451 44251
rect 108850 44248 108856 44260
rect 108439 44220 108856 44248
rect 108439 44217 108451 44220
rect 108393 44211 108451 44217
rect 108850 44208 108856 44220
rect 108908 44208 108914 44260
rect 9674 44180 9680 44192
rect 6886 44152 9680 44180
rect 9674 44140 9680 44152
rect 9732 44140 9738 44192
rect 1104 44090 7912 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 7912 44090
rect 1104 44016 7912 44038
rect 108008 44090 118864 44112
rect 108008 44038 112914 44090
rect 112966 44038 112978 44090
rect 113030 44038 113042 44090
rect 113094 44038 113106 44090
rect 113158 44038 113170 44090
rect 113222 44038 118864 44090
rect 108008 44016 118864 44038
rect 108298 43936 108304 43988
rect 108356 43976 108362 43988
rect 108577 43979 108635 43985
rect 108577 43976 108589 43979
rect 108356 43948 108589 43976
rect 108356 43936 108362 43948
rect 108577 43945 108589 43948
rect 108623 43945 108635 43979
rect 108577 43939 108635 43945
rect 109589 43979 109647 43985
rect 109589 43945 109601 43979
rect 109635 43976 109647 43979
rect 110138 43976 110144 43988
rect 109635 43948 110144 43976
rect 109635 43945 109647 43948
rect 109589 43939 109647 43945
rect 110138 43936 110144 43948
rect 110196 43936 110202 43988
rect 110230 43936 110236 43988
rect 110288 43936 110294 43988
rect 110414 43936 110420 43988
rect 110472 43936 110478 43988
rect 109678 43800 109684 43852
rect 109736 43840 109742 43852
rect 109957 43843 110015 43849
rect 109957 43840 109969 43843
rect 109736 43812 109969 43840
rect 109736 43800 109742 43812
rect 109957 43809 109969 43812
rect 110003 43809 110015 43843
rect 109957 43803 110015 43809
rect 108298 43732 108304 43784
rect 108356 43732 108362 43784
rect 109770 43732 109776 43784
rect 109828 43732 109834 43784
rect 108393 43707 108451 43713
rect 108393 43673 108405 43707
rect 108439 43704 108451 43707
rect 108666 43704 108672 43716
rect 108439 43676 108672 43704
rect 108439 43673 108451 43676
rect 108393 43667 108451 43673
rect 108666 43664 108672 43676
rect 108724 43664 108730 43716
rect 109402 43664 109408 43716
rect 109460 43704 109466 43716
rect 110049 43707 110107 43713
rect 110049 43704 110061 43707
rect 109460 43676 110061 43704
rect 109460 43664 109466 43676
rect 110049 43673 110061 43676
rect 110095 43673 110107 43707
rect 110049 43667 110107 43673
rect 109862 43596 109868 43648
rect 109920 43636 109926 43648
rect 110249 43639 110307 43645
rect 110249 43636 110261 43639
rect 109920 43608 110261 43636
rect 109920 43596 109926 43608
rect 110249 43605 110261 43608
rect 110295 43605 110307 43639
rect 110249 43599 110307 43605
rect 1104 43546 7912 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 7912 43546
rect 1104 43472 7912 43494
rect 108008 43546 118864 43568
rect 108008 43494 113650 43546
rect 113702 43494 113714 43546
rect 113766 43494 113778 43546
rect 113830 43494 113842 43546
rect 113894 43494 113906 43546
rect 113958 43494 118864 43546
rect 108008 43472 118864 43494
rect 109589 43435 109647 43441
rect 109589 43401 109601 43435
rect 109635 43432 109647 43435
rect 110230 43432 110236 43444
rect 109635 43404 110236 43432
rect 109635 43401 109647 43404
rect 109589 43395 109647 43401
rect 110230 43392 110236 43404
rect 110288 43392 110294 43444
rect 109126 43324 109132 43376
rect 109184 43364 109190 43376
rect 109497 43367 109555 43373
rect 109497 43364 109509 43367
rect 109184 43336 109509 43364
rect 109184 43324 109190 43336
rect 109497 43333 109509 43336
rect 109543 43364 109555 43367
rect 109543 43336 109724 43364
rect 109543 43333 109555 43336
rect 109497 43327 109555 43333
rect 1302 43256 1308 43308
rect 1360 43296 1366 43308
rect 1397 43299 1455 43305
rect 1397 43296 1409 43299
rect 1360 43268 1409 43296
rect 1360 43256 1366 43268
rect 1397 43265 1409 43268
rect 1443 43296 1455 43299
rect 1673 43299 1731 43305
rect 1673 43296 1685 43299
rect 1443 43268 1685 43296
rect 1443 43265 1455 43268
rect 1397 43259 1455 43265
rect 1673 43265 1685 43268
rect 1719 43265 1731 43299
rect 1673 43259 1731 43265
rect 109218 43256 109224 43308
rect 109276 43296 109282 43308
rect 109313 43299 109371 43305
rect 109313 43296 109325 43299
rect 109276 43268 109325 43296
rect 109276 43256 109282 43268
rect 109313 43265 109325 43268
rect 109359 43265 109371 43299
rect 109313 43259 109371 43265
rect 109328 43228 109356 43259
rect 109586 43256 109592 43308
rect 109644 43256 109650 43308
rect 109696 43305 109724 43336
rect 109681 43299 109739 43305
rect 109681 43265 109693 43299
rect 109727 43265 109739 43299
rect 109681 43259 109739 43265
rect 109957 43299 110015 43305
rect 109957 43265 109969 43299
rect 110003 43265 110015 43299
rect 109957 43259 110015 43265
rect 109972 43228 110000 43259
rect 110138 43256 110144 43308
rect 110196 43296 110202 43308
rect 110417 43299 110475 43305
rect 110417 43296 110429 43299
rect 110196 43268 110429 43296
rect 110196 43256 110202 43268
rect 110417 43265 110429 43268
rect 110463 43265 110475 43299
rect 110417 43259 110475 43265
rect 109328 43200 110000 43228
rect 1581 43163 1639 43169
rect 1581 43129 1593 43163
rect 1627 43160 1639 43163
rect 9674 43160 9680 43172
rect 1627 43132 9680 43160
rect 1627 43129 1639 43132
rect 1581 43123 1639 43129
rect 9674 43120 9680 43132
rect 9732 43120 9738 43172
rect 109954 43120 109960 43172
rect 110012 43160 110018 43172
rect 110233 43163 110291 43169
rect 110233 43160 110245 43163
rect 110012 43132 110245 43160
rect 110012 43120 110018 43132
rect 110233 43129 110245 43132
rect 110279 43129 110291 43163
rect 110233 43123 110291 43129
rect 109586 43052 109592 43104
rect 109644 43092 109650 43104
rect 109865 43095 109923 43101
rect 109865 43092 109877 43095
rect 109644 43064 109877 43092
rect 109644 43052 109650 43064
rect 109865 43061 109877 43064
rect 109911 43061 109923 43095
rect 109865 43055 109923 43061
rect 110138 43052 110144 43104
rect 110196 43052 110202 43104
rect 1104 43002 7912 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 7912 43002
rect 1104 42928 7912 42950
rect 108008 43002 118864 43024
rect 108008 42950 112914 43002
rect 112966 42950 112978 43002
rect 113030 42950 113042 43002
rect 113094 42950 113106 43002
rect 113158 42950 113170 43002
rect 113222 42950 118864 43002
rect 108008 42928 118864 42950
rect 108298 42848 108304 42900
rect 108356 42888 108362 42900
rect 108669 42891 108727 42897
rect 108669 42888 108681 42891
rect 108356 42860 108681 42888
rect 108356 42848 108362 42860
rect 108408 42693 108436 42860
rect 108669 42857 108681 42860
rect 108715 42857 108727 42891
rect 108669 42851 108727 42857
rect 109862 42848 109868 42900
rect 109920 42848 109926 42900
rect 108393 42687 108451 42693
rect 108393 42653 108405 42687
rect 108439 42653 108451 42687
rect 108393 42647 108451 42653
rect 109405 42687 109463 42693
rect 109405 42653 109417 42687
rect 109451 42653 109463 42687
rect 109405 42647 109463 42653
rect 109420 42616 109448 42647
rect 109494 42644 109500 42696
rect 109552 42644 109558 42696
rect 109681 42687 109739 42693
rect 109681 42653 109693 42687
rect 109727 42684 109739 42687
rect 110138 42684 110144 42696
rect 109727 42656 110144 42684
rect 109727 42653 109739 42656
rect 109681 42647 109739 42653
rect 110138 42644 110144 42656
rect 110196 42644 110202 42696
rect 109586 42616 109592 42628
rect 109420 42588 109592 42616
rect 109586 42576 109592 42588
rect 109644 42616 109650 42628
rect 109862 42616 109868 42628
rect 109644 42588 109868 42616
rect 109644 42576 109650 42588
rect 109862 42576 109868 42588
rect 109920 42576 109926 42628
rect 108482 42508 108488 42560
rect 108540 42508 108546 42560
rect 1104 42458 7912 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 7912 42458
rect 1104 42384 7912 42406
rect 108008 42458 118864 42480
rect 108008 42406 113650 42458
rect 113702 42406 113714 42458
rect 113766 42406 113778 42458
rect 113830 42406 113842 42458
rect 113894 42406 113906 42458
rect 113958 42406 118864 42458
rect 108008 42384 118864 42406
rect 108574 42236 108580 42288
rect 108632 42276 108638 42288
rect 108632 42248 108882 42276
rect 108632 42236 108638 42248
rect 110322 42168 110328 42220
rect 110380 42168 110386 42220
rect 110046 42100 110052 42152
rect 110104 42100 110110 42152
rect 108577 42007 108635 42013
rect 108577 41973 108589 42007
rect 108623 42004 108635 42007
rect 109494 42004 109500 42016
rect 108623 41976 109500 42004
rect 108623 41973 108635 41976
rect 108577 41967 108635 41973
rect 109494 41964 109500 41976
rect 109552 41964 109558 42016
rect 1104 41914 7912 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 7912 41914
rect 1104 41840 7912 41862
rect 108008 41914 118864 41936
rect 108008 41862 112914 41914
rect 112966 41862 112978 41914
rect 113030 41862 113042 41914
rect 113094 41862 113106 41914
rect 113158 41862 113170 41914
rect 113222 41862 118864 41914
rect 108008 41840 118864 41862
rect 108298 41760 108304 41812
rect 108356 41800 108362 41812
rect 108577 41803 108635 41809
rect 108577 41800 108589 41803
rect 108356 41772 108589 41800
rect 108356 41760 108362 41772
rect 108577 41769 108589 41772
rect 108623 41769 108635 41803
rect 108577 41763 108635 41769
rect 109770 41760 109776 41812
rect 109828 41800 109834 41812
rect 109957 41803 110015 41809
rect 109957 41800 109969 41803
rect 109828 41772 109969 41800
rect 109828 41760 109834 41772
rect 109957 41769 109969 41772
rect 110003 41769 110015 41803
rect 109957 41763 110015 41769
rect 108942 41624 108948 41676
rect 109000 41664 109006 41676
rect 109589 41667 109647 41673
rect 109589 41664 109601 41667
rect 109000 41636 109601 41664
rect 109000 41624 109006 41636
rect 109589 41633 109601 41636
rect 109635 41633 109647 41667
rect 110506 41664 110512 41676
rect 109589 41627 109647 41633
rect 109696 41636 110512 41664
rect 108298 41556 108304 41608
rect 108356 41556 108362 41608
rect 109696 41605 109724 41636
rect 110506 41624 110512 41636
rect 110564 41624 110570 41676
rect 109405 41599 109463 41605
rect 109405 41565 109417 41599
rect 109451 41596 109463 41599
rect 109681 41599 109739 41605
rect 109681 41596 109693 41599
rect 109451 41568 109693 41596
rect 109451 41565 109463 41568
rect 109405 41559 109463 41565
rect 109681 41565 109693 41568
rect 109727 41565 109739 41599
rect 110230 41596 110236 41608
rect 109681 41559 109739 41565
rect 109880 41568 110236 41596
rect 109586 41488 109592 41540
rect 109644 41528 109650 41540
rect 109880 41528 109908 41568
rect 110230 41556 110236 41568
rect 110288 41596 110294 41608
rect 110693 41599 110751 41605
rect 110693 41596 110705 41599
rect 110288 41568 110705 41596
rect 110288 41556 110294 41568
rect 110693 41565 110705 41568
rect 110739 41565 110751 41599
rect 110693 41559 110751 41565
rect 110877 41599 110935 41605
rect 110877 41565 110889 41599
rect 110923 41565 110935 41599
rect 110877 41559 110935 41565
rect 109644 41500 109908 41528
rect 109644 41488 109650 41500
rect 110598 41488 110604 41540
rect 110656 41528 110662 41540
rect 110892 41528 110920 41559
rect 110656 41500 110920 41528
rect 110656 41488 110662 41500
rect 108390 41420 108396 41472
rect 108448 41420 108454 41472
rect 110782 41420 110788 41472
rect 110840 41420 110846 41472
rect 1104 41370 7912 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 7912 41370
rect 1104 41296 7912 41318
rect 108008 41370 118864 41392
rect 108008 41318 113650 41370
rect 113702 41318 113714 41370
rect 113766 41318 113778 41370
rect 113830 41318 113842 41370
rect 113894 41318 113906 41370
rect 113958 41318 118864 41370
rect 108008 41296 118864 41318
rect 1302 41080 1308 41132
rect 1360 41120 1366 41132
rect 1397 41123 1455 41129
rect 1397 41120 1409 41123
rect 1360 41092 1409 41120
rect 1360 41080 1366 41092
rect 1397 41089 1409 41092
rect 1443 41120 1455 41123
rect 1673 41123 1731 41129
rect 1673 41120 1685 41123
rect 1443 41092 1685 41120
rect 1443 41089 1455 41092
rect 1397 41083 1455 41089
rect 1673 41089 1685 41092
rect 1719 41089 1731 41123
rect 1673 41083 1731 41089
rect 108758 41080 108764 41132
rect 108816 41120 108822 41132
rect 108942 41120 108948 41132
rect 108816 41092 108948 41120
rect 108816 41080 108822 41092
rect 108942 41080 108948 41092
rect 109000 41080 109006 41132
rect 109678 41080 109684 41132
rect 109736 41120 109742 41132
rect 109862 41120 109868 41132
rect 109736 41092 109868 41120
rect 109736 41080 109742 41092
rect 109862 41080 109868 41092
rect 109920 41120 109926 41132
rect 109957 41123 110015 41129
rect 109957 41120 109969 41123
rect 109920 41092 109969 41120
rect 109920 41080 109926 41092
rect 109957 41089 109969 41092
rect 110003 41089 110015 41123
rect 109957 41083 110015 41089
rect 110230 41080 110236 41132
rect 110288 41120 110294 41132
rect 110417 41123 110475 41129
rect 110417 41120 110429 41123
rect 110288 41092 110429 41120
rect 110288 41080 110294 41092
rect 110417 41089 110429 41092
rect 110463 41089 110475 41123
rect 110417 41083 110475 41089
rect 110598 41080 110604 41132
rect 110656 41080 110662 41132
rect 110874 41080 110880 41132
rect 110932 41080 110938 41132
rect 1581 40987 1639 40993
rect 1581 40953 1593 40987
rect 1627 40984 1639 40987
rect 9674 40984 9680 40996
rect 1627 40956 9680 40984
rect 1627 40953 1639 40956
rect 1581 40947 1639 40953
rect 9674 40944 9680 40956
rect 9732 40944 9738 40996
rect 108942 40944 108948 40996
rect 109000 40984 109006 40996
rect 110322 40984 110328 40996
rect 109000 40956 110328 40984
rect 109000 40944 109006 40956
rect 110322 40944 110328 40956
rect 110380 40944 110386 40996
rect 110141 40919 110199 40925
rect 110141 40885 110153 40919
rect 110187 40916 110199 40919
rect 110230 40916 110236 40928
rect 110187 40888 110236 40916
rect 110187 40885 110199 40888
rect 110141 40879 110199 40885
rect 110230 40876 110236 40888
rect 110288 40876 110294 40928
rect 110506 40876 110512 40928
rect 110564 40916 110570 40928
rect 111061 40919 111119 40925
rect 111061 40916 111073 40919
rect 110564 40888 111073 40916
rect 110564 40876 110570 40888
rect 111061 40885 111073 40888
rect 111107 40885 111119 40919
rect 111061 40879 111119 40885
rect 1104 40826 7912 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 7912 40826
rect 1104 40752 7912 40774
rect 108008 40826 118864 40848
rect 108008 40774 112914 40826
rect 112966 40774 112978 40826
rect 113030 40774 113042 40826
rect 113094 40774 113106 40826
rect 113158 40774 113170 40826
rect 113222 40774 118864 40826
rect 108008 40752 118864 40774
rect 110046 40672 110052 40724
rect 110104 40712 110110 40724
rect 110141 40715 110199 40721
rect 110141 40712 110153 40715
rect 110104 40684 110153 40712
rect 110104 40672 110110 40684
rect 110141 40681 110153 40684
rect 110187 40681 110199 40715
rect 110141 40675 110199 40681
rect 110322 40672 110328 40724
rect 110380 40672 110386 40724
rect 109678 40604 109684 40656
rect 109736 40604 109742 40656
rect 110598 40604 110604 40656
rect 110656 40644 110662 40656
rect 110693 40647 110751 40653
rect 110693 40644 110705 40647
rect 110656 40616 110705 40644
rect 110656 40604 110662 40616
rect 110693 40613 110705 40616
rect 110739 40613 110751 40647
rect 110693 40607 110751 40613
rect 108301 40579 108359 40585
rect 108301 40545 108313 40579
rect 108347 40576 108359 40579
rect 108942 40576 108948 40588
rect 108347 40548 108948 40576
rect 108347 40545 108359 40548
rect 108301 40539 108359 40545
rect 108942 40536 108948 40548
rect 109000 40536 109006 40588
rect 109696 40576 109724 40604
rect 110969 40579 111027 40585
rect 110969 40576 110981 40579
rect 109696 40548 110981 40576
rect 110969 40545 110981 40548
rect 111015 40545 111027 40579
rect 110969 40539 111027 40545
rect 1302 40468 1308 40520
rect 1360 40508 1366 40520
rect 1397 40511 1455 40517
rect 1397 40508 1409 40511
rect 1360 40480 1409 40508
rect 1360 40468 1366 40480
rect 1397 40477 1409 40480
rect 1443 40508 1455 40511
rect 1673 40511 1731 40517
rect 1673 40508 1685 40511
rect 1443 40480 1685 40508
rect 1443 40477 1455 40480
rect 1397 40471 1455 40477
rect 1673 40477 1685 40480
rect 1719 40477 1731 40511
rect 1673 40471 1731 40477
rect 109862 40468 109868 40520
rect 109920 40508 109926 40520
rect 111061 40511 111119 40517
rect 109920 40480 110552 40508
rect 109920 40468 109926 40480
rect 9674 40440 9680 40452
rect 1596 40412 9680 40440
rect 1596 40381 1624 40412
rect 9674 40400 9680 40412
rect 9732 40400 9738 40452
rect 108574 40400 108580 40452
rect 108632 40400 108638 40452
rect 108850 40400 108856 40452
rect 108908 40440 108914 40452
rect 110524 40449 110552 40480
rect 111061 40477 111073 40511
rect 111107 40508 111119 40511
rect 113450 40508 113456 40520
rect 111107 40480 113456 40508
rect 111107 40477 111119 40480
rect 111061 40471 111119 40477
rect 113450 40468 113456 40480
rect 113508 40468 113514 40520
rect 110509 40443 110567 40449
rect 108908 40412 109066 40440
rect 110064 40412 110460 40440
rect 108908 40400 108914 40412
rect 110064 40381 110092 40412
rect 1581 40375 1639 40381
rect 1581 40341 1593 40375
rect 1627 40341 1639 40375
rect 1581 40335 1639 40341
rect 110049 40375 110107 40381
rect 110049 40341 110061 40375
rect 110095 40341 110107 40375
rect 110049 40335 110107 40341
rect 110138 40332 110144 40384
rect 110196 40372 110202 40384
rect 110299 40375 110357 40381
rect 110299 40372 110311 40375
rect 110196 40344 110311 40372
rect 110196 40332 110202 40344
rect 110299 40341 110311 40344
rect 110345 40341 110357 40375
rect 110432 40372 110460 40412
rect 110509 40409 110521 40443
rect 110555 40409 110567 40443
rect 110509 40403 110567 40409
rect 110598 40372 110604 40384
rect 110432 40344 110604 40372
rect 110299 40335 110357 40341
rect 110598 40332 110604 40344
rect 110656 40332 110662 40384
rect 1104 40282 7912 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 7912 40282
rect 1104 40208 7912 40230
rect 108008 40282 118864 40304
rect 108008 40230 113650 40282
rect 113702 40230 113714 40282
rect 113766 40230 113778 40282
rect 113830 40230 113842 40282
rect 113894 40230 113906 40282
rect 113958 40230 118864 40282
rect 108008 40208 118864 40230
rect 109957 40171 110015 40177
rect 109957 40137 109969 40171
rect 110003 40168 110015 40171
rect 110138 40168 110144 40180
rect 110003 40140 110144 40168
rect 110003 40137 110015 40140
rect 109957 40131 110015 40137
rect 110138 40128 110144 40140
rect 110196 40128 110202 40180
rect 110414 40128 110420 40180
rect 110472 40128 110478 40180
rect 110782 40128 110788 40180
rect 110840 40128 110846 40180
rect 109512 40072 110092 40100
rect 109512 40044 109540 40072
rect 109494 39992 109500 40044
rect 109552 39992 109558 40044
rect 109586 39992 109592 40044
rect 109644 39992 109650 40044
rect 109678 39992 109684 40044
rect 109736 39992 109742 40044
rect 109773 40035 109831 40041
rect 109773 40001 109785 40035
rect 109819 40032 109831 40035
rect 109954 40032 109960 40044
rect 109819 40004 109960 40032
rect 109819 40001 109831 40004
rect 109773 39995 109831 40001
rect 109954 39992 109960 40004
rect 110012 39992 110018 40044
rect 110064 40041 110092 40072
rect 110506 40060 110512 40112
rect 110564 40100 110570 40112
rect 110564 40072 110644 40100
rect 110564 40060 110570 40072
rect 110616 40041 110644 40072
rect 110800 40041 110828 40128
rect 110874 40060 110880 40112
rect 110932 40060 110938 40112
rect 110049 40035 110107 40041
rect 110049 40001 110061 40035
rect 110095 40001 110107 40035
rect 110049 39995 110107 40001
rect 110601 40035 110659 40041
rect 110601 40001 110613 40035
rect 110647 40001 110659 40035
rect 110601 39995 110659 40001
rect 110749 40035 110828 40041
rect 110749 40001 110761 40035
rect 110795 40004 110828 40035
rect 110969 40035 111027 40041
rect 110795 40001 110807 40004
rect 110749 39995 110807 40001
rect 110969 40001 110981 40035
rect 111015 40001 111027 40035
rect 110969 39995 111027 40001
rect 111107 40035 111165 40041
rect 111107 40001 111119 40035
rect 111153 40032 111165 40035
rect 111334 40032 111340 40044
rect 111153 40004 111340 40032
rect 111153 40001 111165 40004
rect 111107 39995 111165 40001
rect 110414 39924 110420 39976
rect 110472 39964 110478 39976
rect 110984 39964 111012 39995
rect 111334 39992 111340 40004
rect 111392 39992 111398 40044
rect 110472 39936 111012 39964
rect 110472 39924 110478 39936
rect 110138 39788 110144 39840
rect 110196 39828 110202 39840
rect 110233 39831 110291 39837
rect 110233 39828 110245 39831
rect 110196 39800 110245 39828
rect 110196 39788 110202 39800
rect 110233 39797 110245 39800
rect 110279 39797 110291 39831
rect 110233 39791 110291 39797
rect 111150 39788 111156 39840
rect 111208 39828 111214 39840
rect 111245 39831 111303 39837
rect 111245 39828 111257 39831
rect 111208 39800 111257 39828
rect 111208 39788 111214 39800
rect 111245 39797 111257 39800
rect 111291 39797 111303 39831
rect 111245 39791 111303 39797
rect 1104 39738 7912 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 7912 39738
rect 1104 39664 7912 39686
rect 108008 39738 118864 39760
rect 108008 39686 112914 39738
rect 112966 39686 112978 39738
rect 113030 39686 113042 39738
rect 113094 39686 113106 39738
rect 113158 39686 113170 39738
rect 113222 39686 118864 39738
rect 108008 39664 118864 39686
rect 109770 39584 109776 39636
rect 109828 39624 109834 39636
rect 110230 39624 110236 39636
rect 109828 39596 110236 39624
rect 109828 39584 109834 39596
rect 110230 39584 110236 39596
rect 110288 39584 110294 39636
rect 110690 39584 110696 39636
rect 110748 39584 110754 39636
rect 110233 39491 110291 39497
rect 110233 39457 110245 39491
rect 110279 39488 110291 39491
rect 110414 39488 110420 39500
rect 110279 39460 110420 39488
rect 110279 39457 110291 39460
rect 110233 39451 110291 39457
rect 110414 39448 110420 39460
rect 110472 39488 110478 39500
rect 110708 39488 110736 39584
rect 110472 39460 110736 39488
rect 110472 39448 110478 39460
rect 110509 39423 110567 39429
rect 110509 39389 110521 39423
rect 110555 39389 110567 39423
rect 110509 39383 110567 39389
rect 106918 39312 106924 39364
rect 106976 39352 106982 39364
rect 106976 39324 108620 39352
rect 106976 39312 106982 39324
rect 108206 39244 108212 39296
rect 108264 39284 108270 39296
rect 108485 39287 108543 39293
rect 108485 39284 108497 39287
rect 108264 39256 108497 39284
rect 108264 39244 108270 39256
rect 108485 39253 108497 39256
rect 108531 39253 108543 39287
rect 108592 39284 108620 39324
rect 108666 39312 108672 39364
rect 108724 39352 108730 39364
rect 108724 39324 108790 39352
rect 108724 39312 108730 39324
rect 109678 39312 109684 39364
rect 109736 39352 109742 39364
rect 109957 39355 110015 39361
rect 109957 39352 109969 39355
rect 109736 39324 109969 39352
rect 109736 39312 109742 39324
rect 109957 39321 109969 39324
rect 110003 39321 110015 39355
rect 109957 39315 110015 39321
rect 110230 39312 110236 39364
rect 110288 39352 110294 39364
rect 110524 39352 110552 39383
rect 110288 39324 110552 39352
rect 110288 39312 110294 39324
rect 110325 39287 110383 39293
rect 110325 39284 110337 39287
rect 108592 39256 110337 39284
rect 108485 39247 108543 39253
rect 110325 39253 110337 39256
rect 110371 39253 110383 39287
rect 110325 39247 110383 39253
rect 1104 39194 7912 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 7912 39194
rect 1104 39120 7912 39142
rect 108008 39194 118864 39216
rect 108008 39142 113650 39194
rect 113702 39142 113714 39194
rect 113766 39142 113778 39194
rect 113830 39142 113842 39194
rect 113894 39142 113906 39194
rect 113958 39142 118864 39194
rect 108008 39120 118864 39142
rect 109494 39040 109500 39092
rect 109552 39040 109558 39092
rect 109586 39040 109592 39092
rect 109644 39080 109650 39092
rect 109644 39052 109908 39080
rect 109644 39040 109650 39052
rect 109681 39015 109739 39021
rect 109681 38981 109693 39015
rect 109727 39012 109739 39015
rect 109770 39012 109776 39024
rect 109727 38984 109776 39012
rect 109727 38981 109739 38984
rect 109681 38975 109739 38981
rect 109770 38972 109776 38984
rect 109828 38972 109834 39024
rect 109880 39021 109908 39052
rect 110322 39040 110328 39092
rect 110380 39040 110386 39092
rect 110506 39040 110512 39092
rect 110564 39080 110570 39092
rect 110601 39083 110659 39089
rect 110601 39080 110613 39083
rect 110564 39052 110613 39080
rect 110564 39040 110570 39052
rect 110601 39049 110613 39052
rect 110647 39049 110659 39083
rect 110601 39043 110659 39049
rect 109865 39015 109923 39021
rect 109865 38981 109877 39015
rect 109911 38981 109923 39015
rect 110616 39012 110644 39043
rect 110969 39015 111027 39021
rect 110969 39012 110981 39015
rect 110616 38984 110981 39012
rect 109865 38975 109923 38981
rect 110969 38981 110981 38984
rect 111015 38981 111027 39015
rect 110969 38975 111027 38981
rect 109589 38947 109647 38953
rect 109589 38913 109601 38947
rect 109635 38913 109647 38947
rect 109589 38907 109647 38913
rect 109604 38876 109632 38907
rect 109954 38904 109960 38956
rect 110012 38904 110018 38956
rect 110233 38947 110291 38953
rect 110233 38913 110245 38947
rect 110279 38913 110291 38947
rect 110233 38907 110291 38913
rect 111153 38947 111211 38953
rect 111153 38913 111165 38947
rect 111199 38944 111211 38947
rect 111334 38944 111340 38956
rect 111199 38916 111340 38944
rect 111199 38913 111211 38916
rect 111153 38907 111211 38913
rect 109972 38876 110000 38904
rect 109604 38848 110000 38876
rect 109313 38811 109371 38817
rect 109313 38777 109325 38811
rect 109359 38808 109371 38811
rect 109586 38808 109592 38820
rect 109359 38780 109592 38808
rect 109359 38777 109371 38780
rect 109313 38771 109371 38777
rect 109586 38768 109592 38780
rect 109644 38808 109650 38820
rect 110248 38808 110276 38907
rect 111334 38904 111340 38916
rect 111392 38904 111398 38956
rect 109644 38780 110276 38808
rect 109644 38768 109650 38780
rect 110138 38700 110144 38752
rect 110196 38700 110202 38752
rect 110785 38743 110843 38749
rect 110785 38709 110797 38743
rect 110831 38740 110843 38743
rect 110966 38740 110972 38752
rect 110831 38712 110972 38740
rect 110831 38709 110843 38712
rect 110785 38703 110843 38709
rect 110966 38700 110972 38712
rect 111024 38700 111030 38752
rect 1104 38650 7912 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 7912 38650
rect 1104 38576 7912 38598
rect 108008 38650 118864 38672
rect 108008 38598 112914 38650
rect 112966 38598 112978 38650
rect 113030 38598 113042 38650
rect 113094 38598 113106 38650
rect 113158 38598 113170 38650
rect 113222 38598 118864 38650
rect 108008 38576 118864 38598
rect 110874 38496 110880 38548
rect 110932 38536 110938 38548
rect 111705 38539 111763 38545
rect 111705 38536 111717 38539
rect 110932 38508 111717 38536
rect 110932 38496 110938 38508
rect 111705 38505 111717 38508
rect 111751 38505 111763 38539
rect 111705 38499 111763 38505
rect 108942 38428 108948 38480
rect 109000 38468 109006 38480
rect 109000 38428 109034 38468
rect 109006 38400 109034 38428
rect 110325 38403 110383 38409
rect 110325 38400 110337 38403
rect 109006 38372 110337 38400
rect 110325 38369 110337 38372
rect 110371 38369 110383 38403
rect 110325 38363 110383 38369
rect 1210 38292 1216 38344
rect 1268 38332 1274 38344
rect 1397 38335 1455 38341
rect 1397 38332 1409 38335
rect 1268 38304 1409 38332
rect 1268 38292 1274 38304
rect 1397 38301 1409 38304
rect 1443 38332 1455 38335
rect 1673 38335 1731 38341
rect 1673 38332 1685 38335
rect 1443 38304 1685 38332
rect 1443 38301 1455 38304
rect 1397 38295 1455 38301
rect 1673 38301 1685 38304
rect 1719 38301 1731 38335
rect 1673 38295 1731 38301
rect 111886 38292 111892 38344
rect 111944 38292 111950 38344
rect 112073 38335 112131 38341
rect 112073 38301 112085 38335
rect 112119 38332 112131 38335
rect 112346 38332 112352 38344
rect 112119 38304 112352 38332
rect 112119 38301 112131 38304
rect 112073 38295 112131 38301
rect 112346 38292 112352 38304
rect 112404 38292 112410 38344
rect 9674 38264 9680 38276
rect 1596 38236 9680 38264
rect 1596 38205 1624 38236
rect 9674 38224 9680 38236
rect 9732 38224 9738 38276
rect 108482 38224 108488 38276
rect 108540 38264 108546 38276
rect 108540 38236 108882 38264
rect 108540 38224 108546 38236
rect 110046 38224 110052 38276
rect 110104 38224 110110 38276
rect 1581 38199 1639 38205
rect 1581 38165 1593 38199
rect 1627 38165 1639 38199
rect 1581 38159 1639 38165
rect 108577 38199 108635 38205
rect 108577 38165 108589 38199
rect 108623 38196 108635 38199
rect 108666 38196 108672 38208
rect 108623 38168 108672 38196
rect 108623 38165 108635 38168
rect 108577 38159 108635 38165
rect 108666 38156 108672 38168
rect 108724 38156 108730 38208
rect 1104 38106 7912 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 7912 38106
rect 1104 38032 7912 38054
rect 108008 38106 118864 38128
rect 108008 38054 113650 38106
rect 113702 38054 113714 38106
rect 113766 38054 113778 38106
rect 113830 38054 113842 38106
rect 113894 38054 113906 38106
rect 113958 38054 118864 38106
rect 108008 38032 118864 38054
rect 108574 37952 108580 38004
rect 108632 37992 108638 38004
rect 109129 37995 109187 38001
rect 109129 37992 109141 37995
rect 108632 37964 109141 37992
rect 108632 37952 108638 37964
rect 109129 37961 109141 37964
rect 109175 37961 109187 37995
rect 109129 37955 109187 37961
rect 109773 37995 109831 38001
rect 109773 37961 109785 37995
rect 109819 37992 109831 37995
rect 109862 37992 109868 38004
rect 109819 37964 109868 37992
rect 109819 37961 109831 37964
rect 109773 37955 109831 37961
rect 109862 37952 109868 37964
rect 109920 37952 109926 38004
rect 109310 37933 109316 37936
rect 109297 37927 109316 37933
rect 109297 37893 109309 37927
rect 109297 37887 109316 37893
rect 109310 37884 109316 37887
rect 109368 37884 109374 37936
rect 109402 37884 109408 37936
rect 109460 37924 109466 37936
rect 109497 37927 109555 37933
rect 109497 37924 109509 37927
rect 109460 37896 109509 37924
rect 109460 37884 109466 37896
rect 109497 37893 109509 37896
rect 109543 37893 109555 37927
rect 109497 37887 109555 37893
rect 110138 37884 110144 37936
rect 110196 37924 110202 37936
rect 110196 37896 110736 37924
rect 110196 37884 110202 37896
rect 1302 37816 1308 37868
rect 1360 37856 1366 37868
rect 1397 37859 1455 37865
rect 1397 37856 1409 37859
rect 1360 37828 1409 37856
rect 1360 37816 1366 37828
rect 1397 37825 1409 37828
rect 1443 37856 1455 37859
rect 1673 37859 1731 37865
rect 1673 37856 1685 37859
rect 1443 37828 1685 37856
rect 1443 37825 1455 37828
rect 1397 37819 1455 37825
rect 1673 37825 1685 37828
rect 1719 37825 1731 37859
rect 1673 37819 1731 37825
rect 110417 37859 110475 37865
rect 110417 37825 110429 37859
rect 110463 37856 110475 37859
rect 110598 37856 110604 37868
rect 110463 37828 110604 37856
rect 110463 37825 110475 37828
rect 110417 37819 110475 37825
rect 110598 37816 110604 37828
rect 110656 37816 110662 37868
rect 110708 37865 110736 37896
rect 110693 37859 110751 37865
rect 110693 37825 110705 37859
rect 110739 37825 110751 37859
rect 110693 37819 110751 37825
rect 112533 37859 112591 37865
rect 112533 37825 112545 37859
rect 112579 37856 112591 37859
rect 112806 37856 112812 37868
rect 112579 37828 112812 37856
rect 112579 37825 112591 37828
rect 112533 37819 112591 37825
rect 112806 37816 112812 37828
rect 112864 37816 112870 37868
rect 113450 37816 113456 37868
rect 113508 37816 113514 37868
rect 113913 37859 113971 37865
rect 113913 37825 113925 37859
rect 113959 37856 113971 37859
rect 114554 37856 114560 37868
rect 113959 37828 114560 37856
rect 113959 37825 113971 37828
rect 113913 37819 113971 37825
rect 114554 37816 114560 37828
rect 114612 37816 114618 37868
rect 110049 37791 110107 37797
rect 110049 37757 110061 37791
rect 110095 37788 110107 37791
rect 110322 37788 110328 37800
rect 110095 37760 110328 37788
rect 110095 37757 110107 37760
rect 110049 37751 110107 37757
rect 110322 37748 110328 37760
rect 110380 37748 110386 37800
rect 110782 37748 110788 37800
rect 110840 37748 110846 37800
rect 111886 37748 111892 37800
rect 111944 37788 111950 37800
rect 112257 37791 112315 37797
rect 112257 37788 112269 37791
rect 111944 37760 112269 37788
rect 111944 37748 111950 37760
rect 112257 37757 112269 37760
rect 112303 37757 112315 37791
rect 112257 37751 112315 37757
rect 1581 37723 1639 37729
rect 1581 37689 1593 37723
rect 1627 37720 1639 37723
rect 9490 37720 9496 37732
rect 1627 37692 9496 37720
rect 1627 37689 1639 37692
rect 1581 37683 1639 37689
rect 9490 37680 9496 37692
rect 9548 37680 9554 37732
rect 108758 37680 108764 37732
rect 108816 37720 108822 37732
rect 108816 37692 109356 37720
rect 108816 37680 108822 37692
rect 109328 37661 109356 37692
rect 111058 37680 111064 37732
rect 111116 37680 111122 37732
rect 112272 37720 112300 37751
rect 112346 37748 112352 37800
rect 112404 37748 112410 37800
rect 112441 37791 112499 37797
rect 112441 37757 112453 37791
rect 112487 37788 112499 37791
rect 113468 37788 113496 37816
rect 112487 37760 113496 37788
rect 112487 37757 112499 37760
rect 112441 37751 112499 37757
rect 113818 37748 113824 37800
rect 113876 37748 113882 37800
rect 112272 37692 112484 37720
rect 112456 37664 112484 37692
rect 109313 37655 109371 37661
rect 109313 37621 109325 37655
rect 109359 37621 109371 37655
rect 109313 37615 109371 37621
rect 109954 37612 109960 37664
rect 110012 37652 110018 37664
rect 110141 37655 110199 37661
rect 110141 37652 110153 37655
rect 110012 37624 110153 37652
rect 110012 37612 110018 37624
rect 110141 37621 110153 37624
rect 110187 37621 110199 37655
rect 110141 37615 110199 37621
rect 110279 37655 110337 37661
rect 110279 37621 110291 37655
rect 110325 37652 110337 37655
rect 110506 37652 110512 37664
rect 110325 37624 110512 37652
rect 110325 37621 110337 37624
rect 110279 37615 110337 37621
rect 110506 37612 110512 37624
rect 110564 37612 110570 37664
rect 111242 37612 111248 37664
rect 111300 37652 111306 37664
rect 112073 37655 112131 37661
rect 112073 37652 112085 37655
rect 111300 37624 112085 37652
rect 111300 37612 111306 37624
rect 112073 37621 112085 37624
rect 112119 37621 112131 37655
rect 112073 37615 112131 37621
rect 112438 37612 112444 37664
rect 112496 37612 112502 37664
rect 114094 37612 114100 37664
rect 114152 37612 114158 37664
rect 114462 37612 114468 37664
rect 114520 37612 114526 37664
rect 1104 37562 7912 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 7912 37562
rect 1104 37488 7912 37510
rect 108008 37562 118864 37584
rect 108008 37510 112914 37562
rect 112966 37510 112978 37562
rect 113030 37510 113042 37562
rect 113094 37510 113106 37562
rect 113158 37510 113170 37562
rect 113222 37510 118864 37562
rect 108008 37488 118864 37510
rect 108482 37408 108488 37460
rect 108540 37448 108546 37460
rect 108850 37448 108856 37460
rect 108540 37420 108856 37448
rect 108540 37408 108546 37420
rect 108850 37408 108856 37420
rect 108908 37448 108914 37460
rect 109313 37451 109371 37457
rect 109313 37448 109325 37451
rect 108908 37420 109325 37448
rect 108908 37408 108914 37420
rect 109313 37417 109325 37420
rect 109359 37417 109371 37451
rect 109313 37411 109371 37417
rect 109497 37451 109555 37457
rect 109497 37417 109509 37451
rect 109543 37448 109555 37451
rect 110046 37448 110052 37460
rect 109543 37420 110052 37448
rect 109543 37417 109555 37420
rect 109497 37411 109555 37417
rect 110046 37408 110052 37420
rect 110104 37408 110110 37460
rect 110782 37408 110788 37460
rect 110840 37448 110846 37460
rect 111061 37451 111119 37457
rect 111061 37448 111073 37451
rect 110840 37420 111073 37448
rect 110840 37408 110846 37420
rect 111061 37417 111073 37420
rect 111107 37417 111119 37451
rect 113542 37448 113548 37460
rect 111061 37411 111119 37417
rect 112824 37420 113548 37448
rect 112824 37392 112852 37420
rect 113542 37408 113548 37420
rect 113600 37408 113606 37460
rect 111242 37340 111248 37392
rect 111300 37340 111306 37392
rect 112806 37340 112812 37392
rect 112864 37340 112870 37392
rect 113269 37383 113327 37389
rect 113269 37349 113281 37383
rect 113315 37380 113327 37383
rect 113450 37380 113456 37392
rect 113315 37352 113456 37380
rect 113315 37349 113327 37352
rect 113269 37343 113327 37349
rect 107010 37272 107016 37324
rect 107068 37312 107074 37324
rect 109681 37315 109739 37321
rect 109681 37312 109693 37315
rect 107068 37284 109693 37312
rect 107068 37272 107074 37284
rect 109681 37281 109693 37284
rect 109727 37281 109739 37315
rect 109681 37275 109739 37281
rect 109402 37244 109408 37256
rect 109144 37216 109408 37244
rect 109144 37185 109172 37216
rect 109402 37204 109408 37216
rect 109460 37204 109466 37256
rect 109865 37247 109923 37253
rect 109865 37213 109877 37247
rect 109911 37244 109923 37247
rect 110138 37244 110144 37256
rect 109911 37216 110144 37244
rect 109911 37213 109923 37216
rect 109865 37207 109923 37213
rect 110138 37204 110144 37216
rect 110196 37204 110202 37256
rect 112625 37247 112683 37253
rect 112625 37213 112637 37247
rect 112671 37244 112683 37247
rect 113174 37244 113180 37256
rect 112671 37216 113180 37244
rect 112671 37213 112683 37216
rect 112625 37207 112683 37213
rect 113174 37204 113180 37216
rect 113232 37244 113238 37256
rect 113284 37244 113312 37343
rect 113450 37340 113456 37352
rect 113508 37340 113514 37392
rect 113818 37272 113824 37324
rect 113876 37312 113882 37324
rect 113876 37284 115060 37312
rect 113876 37272 113882 37284
rect 115032 37256 115060 37284
rect 116394 37272 116400 37324
rect 116452 37272 116458 37324
rect 113232 37216 113312 37244
rect 113545 37247 113603 37253
rect 113232 37204 113238 37216
rect 113545 37213 113557 37247
rect 113591 37213 113603 37247
rect 113545 37207 113603 37213
rect 113913 37247 113971 37253
rect 113913 37213 113925 37247
rect 113959 37244 113971 37247
rect 114002 37244 114008 37256
rect 113959 37216 114008 37244
rect 113959 37213 113971 37216
rect 113913 37207 113971 37213
rect 109129 37179 109187 37185
rect 109129 37145 109141 37179
rect 109175 37145 109187 37179
rect 109420 37176 109448 37204
rect 109954 37176 109960 37188
rect 109420 37148 109960 37176
rect 109129 37139 109187 37145
rect 109954 37136 109960 37148
rect 110012 37136 110018 37188
rect 111521 37179 111579 37185
rect 111521 37145 111533 37179
rect 111567 37176 111579 37179
rect 111702 37176 111708 37188
rect 111567 37148 111708 37176
rect 111567 37145 111579 37148
rect 111521 37139 111579 37145
rect 111702 37136 111708 37148
rect 111760 37176 111766 37188
rect 112257 37179 112315 37185
rect 112257 37176 112269 37179
rect 111760 37148 112269 37176
rect 111760 37136 111766 37148
rect 112257 37145 112269 37148
rect 112303 37145 112315 37179
rect 113560 37176 113588 37207
rect 114002 37204 114008 37216
rect 114060 37204 114066 37256
rect 114278 37204 114284 37256
rect 114336 37204 114342 37256
rect 114370 37204 114376 37256
rect 114428 37204 114434 37256
rect 114480 37216 114876 37244
rect 114186 37176 114192 37188
rect 113560 37148 114192 37176
rect 112257 37139 112315 37145
rect 114186 37136 114192 37148
rect 114244 37176 114250 37188
rect 114480 37176 114508 37216
rect 114848 37188 114876 37216
rect 115014 37204 115020 37256
rect 115072 37244 115078 37256
rect 115109 37247 115167 37253
rect 115109 37244 115121 37247
rect 115072 37216 115121 37244
rect 115072 37204 115078 37216
rect 115109 37213 115121 37216
rect 115155 37213 115167 37247
rect 115109 37207 115167 37213
rect 115293 37247 115351 37253
rect 115293 37213 115305 37247
rect 115339 37244 115351 37247
rect 116302 37244 116308 37256
rect 115339 37216 116308 37244
rect 115339 37213 115351 37216
rect 115293 37207 115351 37213
rect 116302 37204 116308 37216
rect 116360 37204 116366 37256
rect 114244 37148 114508 37176
rect 114244 37136 114250 37148
rect 114554 37136 114560 37188
rect 114612 37176 114618 37188
rect 114741 37179 114799 37185
rect 114741 37176 114753 37179
rect 114612 37148 114753 37176
rect 114612 37136 114618 37148
rect 114741 37145 114753 37148
rect 114787 37145 114799 37179
rect 114741 37139 114799 37145
rect 108850 37068 108856 37120
rect 108908 37108 108914 37120
rect 109329 37111 109387 37117
rect 109329 37108 109341 37111
rect 108908 37080 109341 37108
rect 108908 37068 108914 37080
rect 109329 37077 109341 37080
rect 109375 37077 109387 37111
rect 109329 37071 109387 37077
rect 112438 37068 112444 37120
rect 112496 37068 112502 37120
rect 112530 37068 112536 37120
rect 112588 37068 112594 37120
rect 114756 37108 114784 37139
rect 114830 37136 114836 37188
rect 114888 37136 114894 37188
rect 115845 37111 115903 37117
rect 115845 37108 115857 37111
rect 114756 37080 115857 37108
rect 115845 37077 115857 37080
rect 115891 37077 115903 37111
rect 115845 37071 115903 37077
rect 116210 37068 116216 37120
rect 116268 37068 116274 37120
rect 116305 37111 116363 37117
rect 116305 37077 116317 37111
rect 116351 37108 116363 37111
rect 116486 37108 116492 37120
rect 116351 37080 116492 37108
rect 116351 37077 116363 37080
rect 116305 37071 116363 37077
rect 116486 37068 116492 37080
rect 116544 37068 116550 37120
rect 1104 37018 7912 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 7912 37018
rect 1104 36944 7912 36966
rect 108008 37018 118864 37040
rect 108008 36966 113650 37018
rect 113702 36966 113714 37018
rect 113766 36966 113778 37018
rect 113830 36966 113842 37018
rect 113894 36966 113906 37018
rect 113958 36966 118864 37018
rect 108008 36944 118864 36966
rect 110233 36907 110291 36913
rect 110233 36873 110245 36907
rect 110279 36904 110291 36907
rect 110414 36904 110420 36916
rect 110279 36876 110420 36904
rect 110279 36873 110291 36876
rect 110233 36867 110291 36873
rect 108390 36796 108396 36848
rect 108448 36836 108454 36848
rect 108448 36808 108606 36836
rect 108448 36796 108454 36808
rect 110049 36771 110107 36777
rect 110049 36737 110061 36771
rect 110095 36768 110107 36771
rect 110248 36768 110276 36867
rect 110414 36864 110420 36876
rect 110472 36864 110478 36916
rect 112438 36864 112444 36916
rect 112496 36904 112502 36916
rect 113269 36907 113327 36913
rect 113269 36904 113281 36907
rect 112496 36876 113281 36904
rect 112496 36864 112502 36876
rect 113269 36873 113281 36876
rect 113315 36873 113327 36907
rect 113269 36867 113327 36873
rect 114557 36907 114615 36913
rect 114557 36873 114569 36907
rect 114603 36904 114615 36907
rect 114646 36904 114652 36916
rect 114603 36876 114652 36904
rect 114603 36873 114615 36876
rect 114557 36867 114615 36873
rect 114646 36864 114652 36876
rect 114704 36864 114710 36916
rect 114741 36907 114799 36913
rect 114741 36873 114753 36907
rect 114787 36904 114799 36907
rect 114830 36904 114836 36916
rect 114787 36876 114836 36904
rect 114787 36873 114799 36876
rect 114741 36867 114799 36873
rect 114830 36864 114836 36876
rect 114888 36864 114894 36916
rect 116118 36904 116124 36916
rect 115216 36876 116124 36904
rect 111058 36796 111064 36848
rect 111116 36836 111122 36848
rect 111153 36839 111211 36845
rect 111153 36836 111165 36839
rect 111116 36808 111165 36836
rect 111116 36796 111122 36808
rect 111153 36805 111165 36808
rect 111199 36805 111211 36839
rect 111153 36799 111211 36805
rect 112349 36839 112407 36845
rect 112349 36805 112361 36839
rect 112395 36836 112407 36839
rect 112806 36836 112812 36848
rect 112395 36808 112812 36836
rect 112395 36805 112407 36808
rect 112349 36799 112407 36805
rect 112806 36796 112812 36808
rect 112864 36796 112870 36848
rect 114094 36836 114100 36848
rect 113744 36808 114100 36836
rect 110095 36740 110276 36768
rect 110095 36737 110107 36740
rect 110049 36731 110107 36737
rect 111886 36728 111892 36780
rect 111944 36768 111950 36780
rect 112441 36771 112499 36777
rect 112441 36768 112453 36771
rect 111944 36740 112453 36768
rect 111944 36728 111950 36740
rect 112441 36737 112453 36740
rect 112487 36737 112499 36771
rect 113174 36768 113180 36780
rect 112441 36731 112499 36737
rect 112640 36740 113180 36768
rect 109770 36660 109776 36712
rect 109828 36660 109834 36712
rect 110782 36660 110788 36712
rect 110840 36660 110846 36712
rect 111006 36703 111064 36709
rect 111006 36669 111018 36703
rect 111052 36700 111064 36703
rect 111150 36700 111156 36712
rect 111052 36672 111156 36700
rect 111052 36669 111064 36672
rect 111006 36663 111064 36669
rect 111150 36660 111156 36672
rect 111208 36660 111214 36712
rect 112257 36703 112315 36709
rect 112257 36669 112269 36703
rect 112303 36700 112315 36703
rect 112640 36700 112668 36740
rect 113174 36728 113180 36740
rect 113232 36728 113238 36780
rect 113358 36728 113364 36780
rect 113416 36768 113422 36780
rect 113744 36777 113772 36808
rect 114094 36796 114100 36808
rect 114152 36796 114158 36848
rect 114189 36839 114247 36845
rect 114189 36805 114201 36839
rect 114235 36836 114247 36839
rect 114462 36836 114468 36848
rect 114235 36808 114468 36836
rect 114235 36805 114247 36808
rect 114189 36799 114247 36805
rect 114462 36796 114468 36808
rect 114520 36796 114526 36848
rect 115106 36796 115112 36848
rect 115164 36796 115170 36848
rect 113545 36771 113603 36777
rect 113545 36768 113557 36771
rect 113416 36740 113557 36768
rect 113416 36728 113422 36740
rect 113545 36737 113557 36740
rect 113591 36737 113603 36771
rect 113545 36731 113603 36737
rect 113637 36771 113695 36777
rect 113637 36737 113649 36771
rect 113683 36737 113695 36771
rect 113637 36731 113695 36737
rect 113729 36771 113787 36777
rect 113729 36737 113741 36771
rect 113775 36737 113787 36771
rect 113729 36731 113787 36737
rect 113652 36700 113680 36731
rect 113910 36728 113916 36780
rect 113968 36728 113974 36780
rect 114002 36728 114008 36780
rect 114060 36728 114066 36780
rect 114278 36728 114284 36780
rect 114336 36728 114342 36780
rect 114370 36728 114376 36780
rect 114428 36728 114434 36780
rect 114646 36728 114652 36780
rect 114704 36728 114710 36780
rect 114922 36728 114928 36780
rect 114980 36728 114986 36780
rect 115014 36728 115020 36780
rect 115072 36728 115078 36780
rect 115216 36777 115244 36876
rect 116118 36864 116124 36876
rect 116176 36864 116182 36916
rect 116210 36864 116216 36916
rect 116268 36864 116274 36916
rect 115477 36839 115535 36845
rect 115477 36805 115489 36839
rect 115523 36836 115535 36839
rect 115566 36836 115572 36848
rect 115523 36808 115572 36836
rect 115523 36805 115535 36808
rect 115477 36799 115535 36805
rect 115566 36796 115572 36808
rect 115624 36836 115630 36848
rect 116394 36836 116400 36848
rect 115624 36808 116400 36836
rect 115624 36796 115630 36808
rect 116394 36796 116400 36808
rect 116452 36796 116458 36848
rect 115201 36771 115259 36777
rect 115201 36737 115213 36771
rect 115247 36737 115259 36771
rect 115201 36731 115259 36737
rect 115216 36700 115244 36731
rect 115842 36728 115848 36780
rect 115900 36777 115906 36780
rect 115900 36771 115928 36777
rect 115916 36737 115928 36771
rect 115900 36731 115928 36737
rect 115900 36728 115906 36731
rect 116118 36728 116124 36780
rect 116176 36768 116182 36780
rect 116305 36771 116363 36777
rect 116305 36768 116317 36771
rect 116176 36740 116317 36768
rect 116176 36728 116182 36740
rect 116305 36737 116317 36740
rect 116351 36737 116363 36771
rect 116305 36731 116363 36737
rect 112303 36672 112668 36700
rect 112824 36672 113680 36700
rect 114480 36672 115244 36700
rect 115753 36703 115811 36709
rect 112303 36669 112315 36672
rect 112257 36663 112315 36669
rect 108298 36524 108304 36576
rect 108356 36524 108362 36576
rect 110690 36524 110696 36576
rect 110748 36524 110754 36576
rect 110874 36524 110880 36576
rect 110932 36524 110938 36576
rect 112162 36524 112168 36576
rect 112220 36564 112226 36576
rect 112824 36573 112852 36672
rect 113358 36592 113364 36644
rect 113416 36632 113422 36644
rect 114480 36632 114508 36672
rect 115753 36669 115765 36703
rect 115799 36669 115811 36703
rect 116320 36700 116348 36731
rect 116486 36728 116492 36780
rect 116544 36728 116550 36780
rect 116673 36771 116731 36777
rect 116673 36737 116685 36771
rect 116719 36768 116731 36771
rect 116765 36771 116823 36777
rect 116765 36768 116777 36771
rect 116719 36740 116777 36768
rect 116719 36737 116731 36740
rect 116673 36731 116731 36737
rect 116765 36737 116777 36740
rect 116811 36737 116823 36771
rect 116765 36731 116823 36737
rect 116946 36728 116952 36780
rect 117004 36728 117010 36780
rect 117130 36700 117136 36712
rect 116320 36672 117136 36700
rect 115753 36663 115811 36669
rect 113416 36604 114508 36632
rect 115768 36632 115796 36663
rect 117130 36660 117136 36672
rect 117188 36660 117194 36712
rect 116949 36635 117007 36641
rect 116949 36632 116961 36635
rect 115768 36604 116961 36632
rect 113416 36592 113422 36604
rect 116949 36601 116961 36604
rect 116995 36601 117007 36635
rect 116949 36595 117007 36601
rect 112809 36567 112867 36573
rect 112809 36564 112821 36567
rect 112220 36536 112821 36564
rect 112220 36524 112226 36536
rect 112809 36533 112821 36536
rect 112855 36533 112867 36567
rect 112809 36527 112867 36533
rect 113910 36524 113916 36576
rect 113968 36564 113974 36576
rect 114925 36567 114983 36573
rect 114925 36564 114937 36567
rect 113968 36536 114937 36564
rect 113968 36524 113974 36536
rect 114925 36533 114937 36536
rect 114971 36533 114983 36567
rect 114925 36527 114983 36533
rect 115198 36524 115204 36576
rect 115256 36564 115262 36576
rect 115385 36567 115443 36573
rect 115385 36564 115397 36567
rect 115256 36536 115397 36564
rect 115256 36524 115262 36536
rect 115385 36533 115397 36536
rect 115431 36533 115443 36567
rect 115385 36527 115443 36533
rect 1104 36474 7912 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 7912 36474
rect 1104 36400 7912 36422
rect 108008 36474 118864 36496
rect 108008 36422 112914 36474
rect 112966 36422 112978 36474
rect 113030 36422 113042 36474
rect 113094 36422 113106 36474
rect 113158 36422 113170 36474
rect 113222 36422 118864 36474
rect 108008 36400 118864 36422
rect 109313 36363 109371 36369
rect 109313 36329 109325 36363
rect 109359 36360 109371 36363
rect 109402 36360 109408 36372
rect 109359 36332 109408 36360
rect 109359 36329 109371 36332
rect 109313 36323 109371 36329
rect 109402 36320 109408 36332
rect 109460 36320 109466 36372
rect 109497 36363 109555 36369
rect 109497 36329 109509 36363
rect 109543 36360 109555 36363
rect 109678 36360 109684 36372
rect 109543 36332 109684 36360
rect 109543 36329 109555 36332
rect 109497 36323 109555 36329
rect 109678 36320 109684 36332
rect 109736 36320 109742 36372
rect 110782 36320 110788 36372
rect 110840 36320 110846 36372
rect 111797 36363 111855 36369
rect 111797 36329 111809 36363
rect 111843 36360 111855 36363
rect 112530 36360 112536 36372
rect 111843 36332 112536 36360
rect 111843 36329 111855 36332
rect 111797 36323 111855 36329
rect 112530 36320 112536 36332
rect 112588 36320 112594 36372
rect 113358 36360 113364 36372
rect 112916 36332 113364 36360
rect 112346 36252 112352 36304
rect 112404 36292 112410 36304
rect 112916 36292 112944 36332
rect 113358 36320 113364 36332
rect 113416 36320 113422 36372
rect 114465 36363 114523 36369
rect 114465 36329 114477 36363
rect 114511 36360 114523 36363
rect 115014 36360 115020 36372
rect 114511 36332 115020 36360
rect 114511 36329 114523 36332
rect 114465 36323 114523 36329
rect 115014 36320 115020 36332
rect 115072 36320 115078 36372
rect 115566 36320 115572 36372
rect 115624 36320 115630 36372
rect 116581 36363 116639 36369
rect 116581 36329 116593 36363
rect 116627 36360 116639 36363
rect 116946 36360 116952 36372
rect 116627 36332 116952 36360
rect 116627 36329 116639 36332
rect 116581 36323 116639 36329
rect 116946 36320 116952 36332
rect 117004 36320 117010 36372
rect 112404 36264 112944 36292
rect 112993 36295 113051 36301
rect 112404 36252 112410 36264
rect 112993 36261 113005 36295
rect 113039 36292 113051 36295
rect 113542 36292 113548 36304
rect 113039 36264 113548 36292
rect 113039 36261 113051 36264
rect 112993 36255 113051 36261
rect 113542 36252 113548 36264
rect 113600 36292 113606 36304
rect 114370 36292 114376 36304
rect 113600 36264 114376 36292
rect 113600 36252 113606 36264
rect 114370 36252 114376 36264
rect 114428 36252 114434 36304
rect 114922 36252 114928 36304
rect 114980 36292 114986 36304
rect 115382 36292 115388 36304
rect 114980 36264 115388 36292
rect 114980 36252 114986 36264
rect 115382 36252 115388 36264
rect 115440 36292 115446 36304
rect 116397 36295 116455 36301
rect 116397 36292 116409 36295
rect 115440 36264 116409 36292
rect 115440 36252 115446 36264
rect 116397 36261 116409 36264
rect 116443 36261 116455 36295
rect 116397 36255 116455 36261
rect 110966 36184 110972 36236
rect 111024 36184 111030 36236
rect 113361 36227 113419 36233
rect 113361 36224 113373 36227
rect 112272 36196 113373 36224
rect 107102 36116 107108 36168
rect 107160 36156 107166 36168
rect 110141 36159 110199 36165
rect 110141 36156 110153 36159
rect 107160 36128 110153 36156
rect 107160 36116 107166 36128
rect 110141 36125 110153 36128
rect 110187 36125 110199 36159
rect 110141 36119 110199 36125
rect 110230 36116 110236 36168
rect 110288 36156 110294 36168
rect 110325 36159 110383 36165
rect 110325 36156 110337 36159
rect 110288 36128 110337 36156
rect 110288 36116 110294 36128
rect 110325 36125 110337 36128
rect 110371 36156 110383 36159
rect 111061 36159 111119 36165
rect 111061 36156 111073 36159
rect 110371 36128 111073 36156
rect 110371 36125 110383 36128
rect 110325 36119 110383 36125
rect 111061 36125 111073 36128
rect 111107 36125 111119 36159
rect 111061 36119 111119 36125
rect 111976 36159 112034 36165
rect 111976 36125 111988 36159
rect 112022 36156 112034 36159
rect 112272 36156 112300 36196
rect 113361 36193 113373 36196
rect 113407 36193 113419 36227
rect 113637 36227 113695 36233
rect 113637 36224 113649 36227
rect 113361 36187 113419 36193
rect 113468 36196 113649 36224
rect 112022 36128 112300 36156
rect 112022 36125 112034 36128
rect 111976 36119 112034 36125
rect 112346 36116 112352 36168
rect 112404 36116 112410 36168
rect 112438 36116 112444 36168
rect 112496 36116 112502 36168
rect 112530 36116 112536 36168
rect 112588 36156 112594 36168
rect 112588 36128 112760 36156
rect 112588 36116 112594 36128
rect 109034 36048 109040 36100
rect 109092 36088 109098 36100
rect 109129 36091 109187 36097
rect 109129 36088 109141 36091
rect 109092 36060 109141 36088
rect 109092 36048 109098 36060
rect 109129 36057 109141 36060
rect 109175 36088 109187 36091
rect 109862 36088 109868 36100
rect 109175 36060 109868 36088
rect 109175 36057 109187 36060
rect 109129 36051 109187 36057
rect 109862 36048 109868 36060
rect 109920 36048 109926 36100
rect 112070 36048 112076 36100
rect 112128 36048 112134 36100
rect 112162 36048 112168 36100
rect 112220 36048 112226 36100
rect 112732 36088 112760 36128
rect 112806 36116 112812 36168
rect 112864 36156 112870 36168
rect 112901 36159 112959 36165
rect 112901 36156 112913 36159
rect 112864 36128 112913 36156
rect 112864 36116 112870 36128
rect 112901 36125 112913 36128
rect 112947 36125 112959 36159
rect 112901 36119 112959 36125
rect 113082 36116 113088 36168
rect 113140 36156 113146 36168
rect 113177 36159 113235 36165
rect 113177 36156 113189 36159
rect 113140 36128 113189 36156
rect 113140 36116 113146 36128
rect 113177 36125 113189 36128
rect 113223 36125 113235 36159
rect 113177 36119 113235 36125
rect 113266 36116 113272 36168
rect 113324 36156 113330 36168
rect 113468 36156 113496 36196
rect 113637 36193 113649 36196
rect 113683 36193 113695 36227
rect 113637 36187 113695 36193
rect 113729 36227 113787 36233
rect 113729 36193 113741 36227
rect 113775 36224 113787 36227
rect 114094 36224 114100 36236
rect 113775 36196 114100 36224
rect 113775 36193 113787 36196
rect 113729 36187 113787 36193
rect 114094 36184 114100 36196
rect 114152 36184 114158 36236
rect 115017 36227 115075 36233
rect 115017 36224 115029 36227
rect 114572 36196 115029 36224
rect 113324 36128 113496 36156
rect 113545 36159 113603 36165
rect 113324 36116 113330 36128
rect 113545 36125 113557 36159
rect 113591 36125 113603 36159
rect 113545 36119 113603 36125
rect 113560 36088 113588 36119
rect 113818 36116 113824 36168
rect 113876 36116 113882 36168
rect 114002 36116 114008 36168
rect 114060 36116 114066 36168
rect 114462 36088 114468 36100
rect 112732 36060 114468 36088
rect 114462 36048 114468 36060
rect 114520 36048 114526 36100
rect 109218 35980 109224 36032
rect 109276 36020 109282 36032
rect 109329 36023 109387 36029
rect 109329 36020 109341 36023
rect 109276 35992 109341 36020
rect 109276 35980 109282 35992
rect 109329 35989 109341 35992
rect 109375 35989 109387 36023
rect 109329 35983 109387 35989
rect 113266 35980 113272 36032
rect 113324 36020 113330 36032
rect 113818 36020 113824 36032
rect 113324 35992 113824 36020
rect 113324 35980 113330 35992
rect 113818 35980 113824 35992
rect 113876 36020 113882 36032
rect 114572 36020 114600 36196
rect 115017 36193 115029 36196
rect 115063 36224 115075 36227
rect 115198 36224 115204 36236
rect 115063 36196 115204 36224
rect 115063 36193 115075 36196
rect 115017 36187 115075 36193
rect 115198 36184 115204 36196
rect 115256 36184 115262 36236
rect 116118 36224 116124 36236
rect 115860 36196 116124 36224
rect 115293 36159 115351 36165
rect 115293 36125 115305 36159
rect 115339 36156 115351 36159
rect 115750 36156 115756 36168
rect 115339 36128 115756 36156
rect 115339 36125 115351 36128
rect 115293 36119 115351 36125
rect 115198 36048 115204 36100
rect 115256 36088 115262 36100
rect 115308 36088 115336 36119
rect 115750 36116 115756 36128
rect 115808 36116 115814 36168
rect 115860 36165 115888 36196
rect 116118 36184 116124 36196
rect 116176 36184 116182 36236
rect 116489 36227 116547 36233
rect 116489 36193 116501 36227
rect 116535 36224 116547 36227
rect 117406 36224 117412 36236
rect 116535 36196 117412 36224
rect 116535 36193 116547 36196
rect 116489 36187 116547 36193
rect 117406 36184 117412 36196
rect 117464 36184 117470 36236
rect 115845 36159 115903 36165
rect 115845 36125 115857 36159
rect 115891 36125 115903 36159
rect 115845 36119 115903 36125
rect 116029 36159 116087 36165
rect 116029 36125 116041 36159
rect 116075 36156 116087 36159
rect 116075 36128 116348 36156
rect 116075 36125 116087 36128
rect 116029 36119 116087 36125
rect 115256 36060 115336 36088
rect 115256 36048 115262 36060
rect 115474 36048 115480 36100
rect 115532 36088 115538 36100
rect 115569 36091 115627 36097
rect 115569 36088 115581 36091
rect 115532 36060 115581 36088
rect 115532 36048 115538 36060
rect 115569 36057 115581 36060
rect 115615 36088 115627 36091
rect 116121 36091 116179 36097
rect 116121 36088 116133 36091
rect 115615 36060 116133 36088
rect 115615 36057 115627 36060
rect 115569 36051 115627 36057
rect 116121 36057 116133 36060
rect 116167 36057 116179 36091
rect 116320 36088 116348 36128
rect 116854 36116 116860 36168
rect 116912 36116 116918 36168
rect 116946 36116 116952 36168
rect 117004 36116 117010 36168
rect 117130 36116 117136 36168
rect 117188 36116 117194 36168
rect 116486 36088 116492 36100
rect 116320 36060 116492 36088
rect 116121 36051 116179 36057
rect 116486 36048 116492 36060
rect 116544 36088 116550 36100
rect 116964 36088 116992 36116
rect 116544 36060 116992 36088
rect 116544 36048 116550 36060
rect 113876 35992 114600 36020
rect 113876 35980 113882 35992
rect 114830 35980 114836 36032
rect 114888 35980 114894 36032
rect 114922 35980 114928 36032
rect 114980 35980 114986 36032
rect 115290 35980 115296 36032
rect 115348 36020 115354 36032
rect 115385 36023 115443 36029
rect 115385 36020 115397 36023
rect 115348 35992 115397 36020
rect 115348 35980 115354 35992
rect 115385 35989 115397 35992
rect 115431 36020 115443 36023
rect 115845 36023 115903 36029
rect 115845 36020 115857 36023
rect 115431 35992 115857 36020
rect 115431 35989 115443 35992
rect 115385 35983 115443 35989
rect 115845 35989 115857 35992
rect 115891 35989 115903 36023
rect 115845 35983 115903 35989
rect 116765 36023 116823 36029
rect 116765 35989 116777 36023
rect 116811 36020 116823 36023
rect 117314 36020 117320 36032
rect 116811 35992 117320 36020
rect 116811 35989 116823 35992
rect 116765 35983 116823 35989
rect 117314 35980 117320 35992
rect 117372 35980 117378 36032
rect 1104 35930 7912 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 7912 35930
rect 1104 35856 7912 35878
rect 108008 35930 118864 35952
rect 108008 35878 113650 35930
rect 113702 35878 113714 35930
rect 113766 35878 113778 35930
rect 113830 35878 113842 35930
rect 113894 35878 113906 35930
rect 113958 35878 118864 35930
rect 108008 35856 118864 35878
rect 1581 35819 1639 35825
rect 1581 35785 1593 35819
rect 1627 35816 1639 35819
rect 1627 35788 6914 35816
rect 1627 35785 1639 35788
rect 1581 35779 1639 35785
rect 6886 35748 6914 35788
rect 108758 35776 108764 35828
rect 108816 35776 108822 35828
rect 108942 35816 108948 35828
rect 108868 35788 108948 35816
rect 9490 35748 9496 35760
rect 6886 35720 9496 35748
rect 9490 35708 9496 35720
rect 9548 35708 9554 35760
rect 108868 35757 108896 35788
rect 108942 35776 108948 35788
rect 109000 35776 109006 35828
rect 109221 35819 109279 35825
rect 109221 35785 109233 35819
rect 109267 35785 109279 35819
rect 109221 35779 109279 35785
rect 108853 35751 108911 35757
rect 108853 35717 108865 35751
rect 108899 35717 108911 35751
rect 108853 35711 108911 35717
rect 109034 35708 109040 35760
rect 109092 35757 109098 35760
rect 109092 35751 109111 35757
rect 109099 35717 109111 35751
rect 109236 35748 109264 35779
rect 109310 35776 109316 35828
rect 109368 35776 109374 35828
rect 111886 35776 111892 35828
rect 111944 35776 111950 35828
rect 113358 35776 113364 35828
rect 113416 35816 113422 35828
rect 114002 35816 114008 35828
rect 113416 35788 114008 35816
rect 113416 35776 113422 35788
rect 114002 35776 114008 35788
rect 114060 35776 114066 35828
rect 114741 35819 114799 35825
rect 114741 35785 114753 35819
rect 114787 35816 114799 35819
rect 114830 35816 114836 35828
rect 114787 35788 114836 35816
rect 114787 35785 114799 35788
rect 114741 35779 114799 35785
rect 114830 35776 114836 35788
rect 114888 35776 114894 35828
rect 116946 35776 116952 35828
rect 117004 35776 117010 35828
rect 117133 35819 117191 35825
rect 117133 35785 117145 35819
rect 117179 35785 117191 35819
rect 117133 35779 117191 35785
rect 109770 35748 109776 35760
rect 109236 35720 109776 35748
rect 109092 35711 109111 35717
rect 109092 35708 109098 35711
rect 109770 35708 109776 35720
rect 109828 35708 109834 35760
rect 111702 35748 111708 35760
rect 110524 35720 111708 35748
rect 1302 35640 1308 35692
rect 1360 35680 1366 35692
rect 1397 35683 1455 35689
rect 1397 35680 1409 35683
rect 1360 35652 1409 35680
rect 1360 35640 1366 35652
rect 1397 35649 1409 35652
rect 1443 35680 1455 35683
rect 1673 35683 1731 35689
rect 1673 35680 1685 35683
rect 1443 35652 1685 35680
rect 1443 35649 1455 35652
rect 1397 35643 1455 35649
rect 1673 35649 1685 35652
rect 1719 35649 1731 35683
rect 1673 35643 1731 35649
rect 108577 35683 108635 35689
rect 108577 35649 108589 35683
rect 108623 35649 108635 35683
rect 108577 35643 108635 35649
rect 108761 35683 108819 35689
rect 108761 35649 108773 35683
rect 108807 35680 108819 35683
rect 109497 35683 109555 35689
rect 108807 35652 109034 35680
rect 108807 35649 108819 35652
rect 108761 35643 108819 35649
rect 108390 35504 108396 35556
rect 108448 35544 108454 35556
rect 108592 35544 108620 35643
rect 109006 35612 109034 35652
rect 109497 35649 109509 35683
rect 109543 35649 109555 35683
rect 109497 35643 109555 35649
rect 109512 35612 109540 35643
rect 109586 35640 109592 35692
rect 109644 35680 109650 35692
rect 109681 35683 109739 35689
rect 109681 35680 109693 35683
rect 109644 35652 109693 35680
rect 109644 35640 109650 35652
rect 109681 35649 109693 35652
rect 109727 35649 109739 35683
rect 109681 35643 109739 35649
rect 109957 35683 110015 35689
rect 109957 35649 109969 35683
rect 110003 35649 110015 35683
rect 109957 35643 110015 35649
rect 109972 35612 110000 35643
rect 110414 35640 110420 35692
rect 110472 35640 110478 35692
rect 110524 35621 110552 35720
rect 111702 35708 111708 35720
rect 111760 35708 111766 35760
rect 112993 35751 113051 35757
rect 112993 35717 113005 35751
rect 113039 35748 113051 35751
rect 113637 35751 113695 35757
rect 113637 35748 113649 35751
rect 113039 35720 113649 35748
rect 113039 35717 113051 35720
rect 112993 35711 113051 35717
rect 113637 35717 113649 35720
rect 113683 35748 113695 35751
rect 114278 35748 114284 35760
rect 113683 35720 114284 35748
rect 113683 35717 113695 35720
rect 113637 35711 113695 35717
rect 114278 35708 114284 35720
rect 114336 35708 114342 35760
rect 117148 35748 117176 35779
rect 117406 35776 117412 35828
rect 117464 35776 117470 35828
rect 117961 35751 118019 35757
rect 117961 35748 117973 35751
rect 116412 35720 117176 35748
rect 117332 35720 117973 35748
rect 110598 35640 110604 35692
rect 110656 35680 110662 35692
rect 111061 35683 111119 35689
rect 111061 35680 111073 35683
rect 110656 35652 111073 35680
rect 110656 35640 110662 35652
rect 111061 35649 111073 35652
rect 111107 35649 111119 35683
rect 111061 35643 111119 35649
rect 111521 35683 111579 35689
rect 111521 35649 111533 35683
rect 111567 35680 111579 35683
rect 112530 35680 112536 35692
rect 111567 35652 112536 35680
rect 111567 35649 111579 35652
rect 111521 35643 111579 35649
rect 112530 35640 112536 35652
rect 112588 35640 112594 35692
rect 112806 35640 112812 35692
rect 112864 35680 112870 35692
rect 112901 35683 112959 35689
rect 112901 35680 112913 35683
rect 112864 35652 112913 35680
rect 112864 35640 112870 35652
rect 112901 35649 112913 35652
rect 112947 35649 112959 35683
rect 112901 35643 112959 35649
rect 113082 35640 113088 35692
rect 113140 35640 113146 35692
rect 113542 35640 113548 35692
rect 113600 35640 113606 35692
rect 113729 35683 113787 35689
rect 113729 35649 113741 35683
rect 113775 35649 113787 35683
rect 113729 35643 113787 35649
rect 113913 35683 113971 35689
rect 113913 35649 113925 35683
rect 113959 35649 113971 35683
rect 113913 35643 113971 35649
rect 114005 35683 114063 35689
rect 114005 35649 114017 35683
rect 114051 35680 114063 35683
rect 114051 35652 114324 35680
rect 114051 35649 114063 35652
rect 114005 35643 114063 35649
rect 109006 35584 110000 35612
rect 109586 35544 109592 35556
rect 108448 35516 109592 35544
rect 108448 35504 108454 35516
rect 109586 35504 109592 35516
rect 109644 35504 109650 35556
rect 109972 35544 110000 35584
rect 110509 35615 110567 35621
rect 110509 35581 110521 35615
rect 110555 35581 110567 35615
rect 110509 35575 110567 35581
rect 110785 35615 110843 35621
rect 110785 35581 110797 35615
rect 110831 35612 110843 35615
rect 110966 35612 110972 35624
rect 110831 35584 110972 35612
rect 110831 35581 110843 35584
rect 110785 35575 110843 35581
rect 110966 35572 110972 35584
rect 111024 35572 111030 35624
rect 111610 35572 111616 35624
rect 111668 35572 111674 35624
rect 113100 35612 113128 35640
rect 112548 35584 113128 35612
rect 112548 35556 112576 35584
rect 113450 35572 113456 35624
rect 113508 35612 113514 35624
rect 113744 35612 113772 35643
rect 113508 35584 113772 35612
rect 113928 35612 113956 35643
rect 114186 35612 114192 35624
rect 113928 35584 114192 35612
rect 113508 35572 113514 35584
rect 114186 35572 114192 35584
rect 114244 35572 114250 35624
rect 110877 35547 110935 35553
rect 110877 35544 110889 35547
rect 109972 35516 110889 35544
rect 110877 35513 110889 35516
rect 110923 35513 110935 35547
rect 110877 35507 110935 35513
rect 112530 35504 112536 35556
rect 112588 35504 112594 35556
rect 114296 35544 114324 35652
rect 114370 35640 114376 35692
rect 114428 35640 114434 35692
rect 115198 35640 115204 35692
rect 115256 35640 115262 35692
rect 115290 35640 115296 35692
rect 115348 35640 115354 35692
rect 115474 35640 115480 35692
rect 115532 35640 115538 35692
rect 115569 35683 115627 35689
rect 115569 35649 115581 35683
rect 115615 35649 115627 35683
rect 115569 35643 115627 35649
rect 114462 35572 114468 35624
rect 114520 35572 114526 35624
rect 115584 35612 115612 35643
rect 115934 35612 115940 35624
rect 115492 35584 115940 35612
rect 115492 35544 115520 35584
rect 115934 35572 115940 35584
rect 115992 35572 115998 35624
rect 116026 35572 116032 35624
rect 116084 35612 116090 35624
rect 116412 35621 116440 35720
rect 116578 35640 116584 35692
rect 116636 35640 116642 35692
rect 117038 35640 117044 35692
rect 117096 35680 117102 35692
rect 117332 35689 117360 35720
rect 117961 35717 117973 35720
rect 118007 35717 118019 35751
rect 117961 35711 118019 35717
rect 117317 35683 117375 35689
rect 117317 35680 117329 35683
rect 117096 35652 117329 35680
rect 117096 35640 117102 35652
rect 117317 35649 117329 35652
rect 117363 35649 117375 35683
rect 117317 35643 117375 35649
rect 117593 35683 117651 35689
rect 117593 35649 117605 35683
rect 117639 35680 117651 35683
rect 118145 35683 118203 35689
rect 117639 35652 117820 35680
rect 117639 35649 117651 35652
rect 117593 35643 117651 35649
rect 116397 35615 116455 35621
rect 116397 35612 116409 35615
rect 116084 35584 116409 35612
rect 116084 35572 116090 35584
rect 116397 35581 116409 35584
rect 116443 35581 116455 35615
rect 116397 35575 116455 35581
rect 116489 35615 116547 35621
rect 116489 35581 116501 35615
rect 116535 35581 116547 35615
rect 116489 35575 116547 35581
rect 114296 35516 115520 35544
rect 115566 35504 115572 35556
rect 115624 35544 115630 35556
rect 116504 35544 116532 35575
rect 115624 35516 116532 35544
rect 117792 35544 117820 35652
rect 118145 35649 118157 35683
rect 118191 35649 118203 35683
rect 118145 35643 118203 35649
rect 117866 35572 117872 35624
rect 117924 35612 117930 35624
rect 118160 35612 118188 35643
rect 118234 35640 118240 35692
rect 118292 35640 118298 35692
rect 117924 35584 118188 35612
rect 117924 35572 117930 35584
rect 117961 35547 118019 35553
rect 117961 35544 117973 35547
rect 117792 35516 117973 35544
rect 115624 35504 115630 35516
rect 117961 35513 117973 35516
rect 118007 35513 118019 35547
rect 117961 35507 118019 35513
rect 109034 35436 109040 35488
rect 109092 35436 109098 35488
rect 109494 35436 109500 35488
rect 109552 35476 109558 35488
rect 109773 35479 109831 35485
rect 109773 35476 109785 35479
rect 109552 35448 109785 35476
rect 109552 35436 109558 35448
rect 109773 35445 109785 35448
rect 109819 35445 109831 35479
rect 109773 35439 109831 35445
rect 115017 35479 115075 35485
rect 115017 35445 115029 35479
rect 115063 35476 115075 35479
rect 115198 35476 115204 35488
rect 115063 35448 115204 35476
rect 115063 35445 115075 35448
rect 115017 35439 115075 35445
rect 115198 35436 115204 35448
rect 115256 35436 115262 35488
rect 117777 35479 117835 35485
rect 117777 35445 117789 35479
rect 117823 35476 117835 35479
rect 118234 35476 118240 35488
rect 117823 35448 118240 35476
rect 117823 35445 117835 35448
rect 117777 35439 117835 35445
rect 118234 35436 118240 35448
rect 118292 35436 118298 35488
rect 1104 35386 7912 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 7912 35386
rect 1104 35312 7912 35334
rect 108008 35386 118864 35408
rect 108008 35334 112914 35386
rect 112966 35334 112978 35386
rect 113030 35334 113042 35386
rect 113094 35334 113106 35386
rect 113158 35334 113170 35386
rect 113222 35334 118864 35386
rect 108008 35312 118864 35334
rect 109034 35232 109040 35284
rect 109092 35272 109098 35284
rect 109221 35275 109279 35281
rect 109221 35272 109233 35275
rect 109092 35244 109233 35272
rect 109092 35232 109098 35244
rect 109221 35241 109233 35244
rect 109267 35241 109279 35275
rect 109221 35235 109279 35241
rect 111610 35232 111616 35284
rect 111668 35232 111674 35284
rect 112257 35275 112315 35281
rect 112257 35241 112269 35275
rect 112303 35272 112315 35275
rect 112438 35272 112444 35284
rect 112303 35244 112444 35272
rect 112303 35241 112315 35244
rect 112257 35235 112315 35241
rect 112438 35232 112444 35244
rect 112496 35232 112502 35284
rect 112530 35232 112536 35284
rect 112588 35272 112594 35284
rect 112809 35275 112867 35281
rect 112809 35272 112821 35275
rect 112588 35244 112821 35272
rect 112588 35232 112594 35244
rect 112809 35241 112821 35244
rect 112855 35241 112867 35275
rect 112809 35235 112867 35241
rect 112990 35232 112996 35284
rect 113048 35272 113054 35284
rect 113048 35244 113772 35272
rect 113048 35232 113054 35244
rect 110325 35207 110383 35213
rect 110325 35173 110337 35207
rect 110371 35204 110383 35207
rect 110874 35204 110880 35216
rect 110371 35176 110880 35204
rect 110371 35173 110383 35176
rect 110325 35167 110383 35173
rect 110874 35164 110880 35176
rect 110932 35164 110938 35216
rect 112070 35164 112076 35216
rect 112128 35204 112134 35216
rect 112625 35207 112683 35213
rect 112625 35204 112637 35207
rect 112128 35176 112637 35204
rect 112128 35164 112134 35176
rect 112625 35173 112637 35176
rect 112671 35173 112683 35207
rect 112625 35167 112683 35173
rect 113266 35164 113272 35216
rect 113324 35204 113330 35216
rect 113634 35204 113640 35216
rect 113324 35176 113640 35204
rect 113324 35164 113330 35176
rect 113634 35164 113640 35176
rect 113692 35164 113698 35216
rect 113744 35204 113772 35244
rect 114094 35232 114100 35284
rect 114152 35232 114158 35284
rect 114925 35275 114983 35281
rect 114925 35241 114937 35275
rect 114971 35272 114983 35275
rect 115106 35272 115112 35284
rect 114971 35244 115112 35272
rect 114971 35241 114983 35244
rect 114925 35235 114983 35241
rect 115106 35232 115112 35244
rect 115164 35232 115170 35284
rect 116489 35275 116547 35281
rect 116489 35241 116501 35275
rect 116535 35272 116547 35275
rect 116578 35272 116584 35284
rect 116535 35244 116584 35272
rect 116535 35241 116547 35244
rect 116489 35235 116547 35241
rect 116578 35232 116584 35244
rect 116636 35232 116642 35284
rect 117314 35232 117320 35284
rect 117372 35232 117378 35284
rect 118234 35232 118240 35284
rect 118292 35272 118298 35284
rect 118513 35275 118571 35281
rect 118513 35272 118525 35275
rect 118292 35244 118525 35272
rect 118292 35232 118298 35244
rect 118513 35241 118525 35244
rect 118559 35241 118571 35275
rect 118513 35235 118571 35241
rect 113744 35176 114324 35204
rect 110049 35139 110107 35145
rect 110049 35105 110061 35139
rect 110095 35136 110107 35139
rect 111242 35136 111248 35148
rect 110095 35108 111248 35136
rect 110095 35105 110107 35108
rect 110049 35099 110107 35105
rect 111242 35096 111248 35108
rect 111300 35096 111306 35148
rect 111429 35139 111487 35145
rect 111429 35105 111441 35139
rect 111475 35105 111487 35139
rect 111429 35099 111487 35105
rect 112548 35108 113220 35136
rect 108758 35028 108764 35080
rect 108816 35068 108822 35080
rect 109313 35071 109371 35077
rect 109313 35068 109325 35071
rect 108816 35040 109325 35068
rect 108816 35028 108822 35040
rect 109313 35037 109325 35040
rect 109359 35037 109371 35071
rect 109313 35031 109371 35037
rect 109957 35071 110015 35077
rect 109957 35037 109969 35071
rect 110003 35068 110015 35071
rect 110598 35068 110604 35080
rect 110003 35040 110604 35068
rect 110003 35037 110015 35040
rect 109957 35031 110015 35037
rect 110598 35028 110604 35040
rect 110656 35028 110662 35080
rect 111337 35071 111395 35077
rect 111337 35037 111349 35071
rect 111383 35037 111395 35071
rect 111444 35068 111472 35099
rect 112548 35077 112576 35108
rect 112533 35071 112591 35077
rect 111444 35040 112484 35068
rect 111337 35031 111395 35037
rect 111352 35000 111380 35031
rect 111978 35000 111984 35012
rect 111352 34972 111984 35000
rect 111978 34960 111984 34972
rect 112036 35000 112042 35012
rect 112257 35003 112315 35009
rect 112257 35000 112269 35003
rect 112036 34972 112269 35000
rect 112036 34960 112042 34972
rect 112257 34969 112269 34972
rect 112303 34969 112315 35003
rect 112456 35000 112484 35040
rect 112533 35037 112545 35071
rect 112579 35037 112591 35071
rect 112533 35031 112591 35037
rect 112898 35028 112904 35080
rect 112956 35028 112962 35080
rect 113192 35077 113220 35108
rect 113450 35096 113456 35148
rect 113508 35136 113514 35148
rect 113729 35139 113787 35145
rect 113729 35136 113741 35139
rect 113508 35108 113741 35136
rect 113508 35096 113514 35108
rect 113729 35105 113741 35108
rect 113775 35105 113787 35139
rect 113729 35099 113787 35105
rect 113821 35139 113879 35145
rect 113821 35105 113833 35139
rect 113867 35136 113879 35139
rect 114186 35136 114192 35148
rect 113867 35108 114192 35136
rect 113867 35105 113879 35108
rect 113821 35099 113879 35105
rect 114186 35096 114192 35108
rect 114244 35096 114250 35148
rect 114296 35136 114324 35176
rect 114554 35164 114560 35216
rect 114612 35204 114618 35216
rect 115017 35207 115075 35213
rect 115017 35204 115029 35207
rect 114612 35176 115029 35204
rect 114612 35164 114618 35176
rect 115017 35173 115029 35176
rect 115063 35173 115075 35207
rect 115017 35167 115075 35173
rect 114646 35136 114652 35148
rect 114296 35108 114652 35136
rect 113177 35071 113235 35077
rect 113177 35037 113189 35071
rect 113223 35068 113235 35071
rect 113358 35068 113364 35080
rect 113223 35040 113364 35068
rect 113223 35037 113235 35040
rect 113177 35031 113235 35037
rect 113358 35028 113364 35040
rect 113416 35028 113422 35080
rect 113545 35071 113603 35077
rect 113545 35037 113557 35071
rect 113591 35037 113603 35071
rect 113545 35031 113603 35037
rect 112806 35000 112812 35012
rect 112456 34972 112812 35000
rect 112257 34963 112315 34969
rect 112806 34960 112812 34972
rect 112864 35000 112870 35012
rect 113560 35000 113588 35031
rect 113634 35028 113640 35080
rect 113692 35028 113698 35080
rect 114296 35077 114324 35108
rect 114646 35096 114652 35108
rect 114704 35096 114710 35148
rect 115569 35139 115627 35145
rect 115569 35136 115581 35139
rect 114756 35108 115581 35136
rect 114005 35071 114063 35077
rect 114005 35037 114017 35071
rect 114051 35068 114063 35071
rect 114097 35071 114155 35077
rect 114097 35068 114109 35071
rect 114051 35040 114109 35068
rect 114051 35037 114063 35040
rect 114005 35031 114063 35037
rect 114097 35037 114109 35040
rect 114143 35037 114155 35071
rect 114097 35031 114155 35037
rect 114281 35071 114339 35077
rect 114281 35037 114293 35071
rect 114327 35037 114339 35071
rect 114281 35031 114339 35037
rect 114112 35000 114140 35031
rect 114462 35028 114468 35080
rect 114520 35028 114526 35080
rect 114756 35077 114784 35108
rect 115569 35105 115581 35108
rect 115615 35105 115627 35139
rect 115569 35099 115627 35105
rect 116118 35096 116124 35148
rect 116176 35096 116182 35148
rect 117590 35096 117596 35148
rect 117648 35096 117654 35148
rect 114741 35071 114799 35077
rect 114741 35037 114753 35071
rect 114787 35037 114799 35071
rect 114741 35031 114799 35037
rect 115198 35028 115204 35080
rect 115256 35028 115262 35080
rect 115290 35028 115296 35080
rect 115348 35028 115354 35080
rect 115474 35028 115480 35080
rect 115532 35028 115538 35080
rect 115661 35071 115719 35077
rect 115661 35037 115673 35071
rect 115707 35037 115719 35071
rect 115661 35031 115719 35037
rect 116213 35071 116271 35077
rect 116213 35037 116225 35071
rect 116259 35068 116271 35071
rect 116302 35068 116308 35080
rect 116259 35040 116308 35068
rect 116259 35037 116271 35040
rect 116213 35031 116271 35037
rect 115216 35000 115244 35028
rect 112864 34972 113404 35000
rect 113560 34972 114048 35000
rect 114112 34972 115244 35000
rect 115676 35000 115704 35031
rect 116302 35028 116308 35040
rect 116360 35028 116366 35080
rect 117409 35071 117467 35077
rect 117409 35037 117421 35071
rect 117455 35068 117467 35071
rect 117608 35068 117636 35096
rect 117455 35040 117636 35068
rect 117685 35071 117743 35077
rect 117455 35037 117467 35040
rect 117409 35031 117467 35037
rect 117685 35037 117697 35071
rect 117731 35037 117743 35071
rect 117685 35031 117743 35037
rect 116486 35000 116492 35012
rect 115676 34972 116492 35000
rect 112864 34960 112870 34972
rect 110598 34892 110604 34944
rect 110656 34932 110662 34944
rect 111058 34932 111064 34944
rect 110656 34904 111064 34932
rect 110656 34892 110662 34904
rect 111058 34892 111064 34904
rect 111116 34892 111122 34944
rect 112441 34935 112499 34941
rect 112441 34901 112453 34935
rect 112487 34932 112499 34935
rect 112990 34932 112996 34944
rect 112487 34904 112996 34932
rect 112487 34901 112499 34904
rect 112441 34895 112499 34901
rect 112990 34892 112996 34904
rect 113048 34892 113054 34944
rect 113376 34941 113404 34972
rect 114020 34944 114048 34972
rect 116486 34960 116492 34972
rect 116544 34960 116550 35012
rect 117130 34960 117136 35012
rect 117188 35000 117194 35012
rect 117700 35000 117728 35031
rect 117958 35000 117964 35012
rect 117188 34972 117964 35000
rect 117188 34960 117194 34972
rect 117958 34960 117964 34972
rect 118016 34960 118022 35012
rect 118142 34960 118148 35012
rect 118200 34960 118206 35012
rect 118326 34960 118332 35012
rect 118384 34960 118390 35012
rect 113361 34935 113419 34941
rect 113361 34901 113373 34935
rect 113407 34901 113419 34935
rect 113361 34895 113419 34901
rect 114002 34892 114008 34944
rect 114060 34892 114066 34944
rect 114094 34892 114100 34944
rect 114152 34932 114158 34944
rect 114370 34932 114376 34944
rect 114152 34904 114376 34932
rect 114152 34892 114158 34904
rect 114370 34892 114376 34904
rect 114428 34932 114434 34944
rect 114557 34935 114615 34941
rect 114557 34932 114569 34935
rect 114428 34904 114569 34932
rect 114428 34892 114434 34904
rect 114557 34901 114569 34904
rect 114603 34901 114615 34935
rect 114557 34895 114615 34901
rect 114646 34892 114652 34944
rect 114704 34932 114710 34944
rect 115290 34932 115296 34944
rect 114704 34904 115296 34932
rect 114704 34892 114710 34904
rect 115290 34892 115296 34904
rect 115348 34892 115354 34944
rect 117222 34892 117228 34944
rect 117280 34932 117286 34944
rect 117866 34932 117872 34944
rect 117280 34904 117872 34932
rect 117280 34892 117286 34904
rect 117866 34892 117872 34904
rect 117924 34932 117930 34944
rect 118053 34935 118111 34941
rect 118053 34932 118065 34935
rect 117924 34904 118065 34932
rect 117924 34892 117930 34904
rect 118053 34901 118065 34904
rect 118099 34901 118111 34935
rect 118053 34895 118111 34901
rect 1104 34842 7912 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 7912 34842
rect 1104 34768 7912 34790
rect 108008 34842 118864 34864
rect 108008 34790 113650 34842
rect 113702 34790 113714 34842
rect 113766 34790 113778 34842
rect 113830 34790 113842 34842
rect 113894 34790 113906 34842
rect 113958 34790 118864 34842
rect 108008 34768 118864 34790
rect 108482 34688 108488 34740
rect 108540 34728 108546 34740
rect 108577 34731 108635 34737
rect 108577 34728 108589 34731
rect 108540 34700 108589 34728
rect 108540 34688 108546 34700
rect 108577 34697 108589 34700
rect 108623 34697 108635 34731
rect 108577 34691 108635 34697
rect 109218 34688 109224 34740
rect 109276 34688 109282 34740
rect 109402 34688 109408 34740
rect 109460 34688 109466 34740
rect 109681 34731 109739 34737
rect 109681 34697 109693 34731
rect 109727 34728 109739 34731
rect 109727 34700 111196 34728
rect 109727 34697 109739 34700
rect 109681 34691 109739 34697
rect 108206 34620 108212 34672
rect 108264 34660 108270 34672
rect 108264 34632 109034 34660
rect 108264 34620 108270 34632
rect 109006 34604 109034 34632
rect 109954 34620 109960 34672
rect 110012 34620 110018 34672
rect 110690 34620 110696 34672
rect 110748 34620 110754 34672
rect 110953 34663 111011 34669
rect 110953 34629 110965 34663
rect 110999 34660 111011 34663
rect 111058 34660 111064 34672
rect 110999 34632 111064 34660
rect 110999 34629 111011 34632
rect 110953 34623 111011 34629
rect 111058 34620 111064 34632
rect 111116 34620 111122 34672
rect 111168 34669 111196 34700
rect 111242 34688 111248 34740
rect 111300 34728 111306 34740
rect 111974 34731 112032 34737
rect 111974 34728 111986 34731
rect 111300 34700 111986 34728
rect 111300 34688 111306 34700
rect 111974 34697 111986 34700
rect 112020 34697 112032 34731
rect 111974 34691 112032 34697
rect 112070 34688 112076 34740
rect 112128 34728 112134 34740
rect 112128 34700 113680 34728
rect 112128 34688 112134 34700
rect 111153 34663 111211 34669
rect 111153 34629 111165 34663
rect 111199 34629 111211 34663
rect 111153 34623 111211 34629
rect 108482 34552 108488 34604
rect 108540 34552 108546 34604
rect 108574 34552 108580 34604
rect 108632 34592 108638 34604
rect 108669 34595 108727 34601
rect 108669 34592 108681 34595
rect 108632 34564 108681 34592
rect 108632 34552 108638 34564
rect 108669 34561 108681 34564
rect 108715 34561 108727 34595
rect 108669 34555 108727 34561
rect 108758 34552 108764 34604
rect 108816 34592 108822 34604
rect 108853 34595 108911 34601
rect 108853 34592 108865 34595
rect 108816 34564 108865 34592
rect 108816 34552 108822 34564
rect 108853 34561 108865 34564
rect 108899 34561 108911 34595
rect 109006 34564 109040 34604
rect 108853 34555 108911 34561
rect 108868 34524 108896 34555
rect 109034 34552 109040 34564
rect 109092 34592 109098 34604
rect 109313 34595 109371 34601
rect 109313 34592 109325 34595
rect 109092 34564 109325 34592
rect 109092 34552 109098 34564
rect 109313 34561 109325 34564
rect 109359 34561 109371 34595
rect 109313 34555 109371 34561
rect 109497 34595 109555 34601
rect 109497 34561 109509 34595
rect 109543 34561 109555 34595
rect 109497 34555 109555 34561
rect 109589 34595 109647 34601
rect 109589 34561 109601 34595
rect 109635 34561 109647 34595
rect 109589 34555 109647 34561
rect 109865 34595 109923 34601
rect 109865 34561 109877 34595
rect 109911 34592 109923 34595
rect 110598 34592 110604 34604
rect 109911 34564 110604 34592
rect 109911 34561 109923 34564
rect 109865 34555 109923 34561
rect 109512 34524 109540 34555
rect 108868 34496 109540 34524
rect 109604 34524 109632 34555
rect 110598 34552 110604 34564
rect 110656 34552 110662 34604
rect 109954 34524 109960 34536
rect 109604 34496 109960 34524
rect 109954 34484 109960 34496
rect 110012 34484 110018 34536
rect 110322 34484 110328 34536
rect 110380 34484 110386 34536
rect 111168 34524 111196 34623
rect 111334 34620 111340 34672
rect 111392 34660 111398 34672
rect 112257 34663 112315 34669
rect 112257 34660 112269 34663
rect 111392 34632 112269 34660
rect 111392 34620 111398 34632
rect 112257 34629 112269 34632
rect 112303 34629 112315 34663
rect 112257 34623 112315 34629
rect 111702 34552 111708 34604
rect 111760 34592 111766 34604
rect 111797 34595 111855 34601
rect 111797 34592 111809 34595
rect 111760 34564 111809 34592
rect 111760 34552 111766 34564
rect 111797 34561 111809 34564
rect 111843 34561 111855 34595
rect 111797 34555 111855 34561
rect 111889 34595 111947 34601
rect 111889 34561 111901 34595
rect 111935 34592 111947 34595
rect 112073 34595 112131 34601
rect 111935 34564 112024 34592
rect 111935 34561 111947 34564
rect 111889 34555 111947 34561
rect 111168 34496 111932 34524
rect 111904 34468 111932 34496
rect 110506 34416 110512 34468
rect 110564 34465 110570 34468
rect 110564 34459 110586 34465
rect 110574 34425 110586 34459
rect 110564 34419 110586 34425
rect 110564 34416 110570 34419
rect 111886 34416 111892 34468
rect 111944 34416 111950 34468
rect 111996 34456 112024 34564
rect 112073 34561 112085 34595
rect 112119 34561 112131 34595
rect 112073 34555 112131 34561
rect 112349 34595 112407 34601
rect 112349 34561 112361 34595
rect 112395 34592 112407 34595
rect 113652 34592 113680 34700
rect 114094 34688 114100 34740
rect 114152 34688 114158 34740
rect 114373 34731 114431 34737
rect 114373 34697 114385 34731
rect 114419 34728 114431 34731
rect 114462 34728 114468 34740
rect 114419 34700 114468 34728
rect 114419 34697 114431 34700
rect 114373 34691 114431 34697
rect 114462 34688 114468 34700
rect 114520 34688 114526 34740
rect 116029 34731 116087 34737
rect 116029 34697 116041 34731
rect 116075 34728 116087 34731
rect 116118 34728 116124 34740
rect 116075 34700 116124 34728
rect 116075 34697 116087 34700
rect 116029 34691 116087 34697
rect 116118 34688 116124 34700
rect 116176 34688 116182 34740
rect 114922 34660 114928 34672
rect 114664 34632 114928 34660
rect 113729 34595 113787 34601
rect 113729 34592 113741 34595
rect 112395 34564 113588 34592
rect 113652 34564 113741 34592
rect 112395 34561 112407 34564
rect 112349 34555 112407 34561
rect 112088 34524 112116 34555
rect 113560 34536 113588 34564
rect 113729 34561 113741 34564
rect 113775 34592 113787 34595
rect 114094 34592 114100 34604
rect 113775 34564 114100 34592
rect 113775 34561 113787 34564
rect 113729 34555 113787 34561
rect 114094 34552 114100 34564
rect 114152 34552 114158 34604
rect 114189 34599 114247 34605
rect 114189 34565 114201 34599
rect 114235 34592 114247 34599
rect 114278 34592 114284 34604
rect 114235 34565 114284 34592
rect 114189 34564 114284 34565
rect 114189 34559 114247 34564
rect 114278 34552 114284 34564
rect 114336 34552 114342 34604
rect 112088 34496 113496 34524
rect 113468 34456 113496 34496
rect 113542 34484 113548 34536
rect 113600 34484 113606 34536
rect 113821 34527 113879 34533
rect 113821 34493 113833 34527
rect 113867 34524 113879 34527
rect 114664 34524 114692 34632
rect 114922 34620 114928 34632
rect 114980 34660 114986 34672
rect 115474 34660 115480 34672
rect 114980 34632 115480 34660
rect 114980 34620 114986 34632
rect 115474 34620 115480 34632
rect 115532 34620 115538 34672
rect 115014 34552 115020 34604
rect 115072 34552 115078 34604
rect 115658 34552 115664 34604
rect 115716 34552 115722 34604
rect 117222 34552 117228 34604
rect 117280 34552 117286 34604
rect 117498 34552 117504 34604
rect 117556 34552 117562 34604
rect 117682 34552 117688 34604
rect 117740 34552 117746 34604
rect 113867 34496 114692 34524
rect 113867 34493 113879 34496
rect 113821 34487 113879 34493
rect 114554 34456 114560 34468
rect 111996 34428 113220 34456
rect 113468 34428 114560 34456
rect 109862 34348 109868 34400
rect 109920 34348 109926 34400
rect 110138 34348 110144 34400
rect 110196 34388 110202 34400
rect 110417 34391 110475 34397
rect 110417 34388 110429 34391
rect 110196 34360 110429 34388
rect 110196 34348 110202 34360
rect 110417 34357 110429 34360
rect 110463 34357 110475 34391
rect 110417 34351 110475 34357
rect 110782 34348 110788 34400
rect 110840 34348 110846 34400
rect 110966 34348 110972 34400
rect 111024 34348 111030 34400
rect 111610 34348 111616 34400
rect 111668 34388 111674 34400
rect 111996 34388 112024 34428
rect 111668 34360 112024 34388
rect 113192 34388 113220 34428
rect 114554 34416 114560 34428
rect 114612 34416 114618 34468
rect 114664 34465 114692 34496
rect 115106 34484 115112 34536
rect 115164 34484 115170 34536
rect 115293 34527 115351 34533
rect 115293 34493 115305 34527
rect 115339 34493 115351 34527
rect 115293 34487 115351 34493
rect 114649 34459 114707 34465
rect 114649 34425 114661 34459
rect 114695 34425 114707 34459
rect 114649 34419 114707 34425
rect 115308 34456 115336 34487
rect 115566 34484 115572 34536
rect 115624 34484 115630 34536
rect 116026 34524 116032 34536
rect 115676 34496 116032 34524
rect 115676 34456 115704 34496
rect 116026 34484 116032 34496
rect 116084 34484 116090 34536
rect 117317 34527 117375 34533
rect 117317 34493 117329 34527
rect 117363 34524 117375 34527
rect 117774 34524 117780 34536
rect 117363 34496 117780 34524
rect 117363 34493 117375 34496
rect 117317 34487 117375 34493
rect 117774 34484 117780 34496
rect 117832 34524 117838 34536
rect 118326 34524 118332 34536
rect 117832 34496 118332 34524
rect 117832 34484 117838 34496
rect 118326 34484 118332 34496
rect 118384 34484 118390 34536
rect 115308 34428 115704 34456
rect 113726 34388 113732 34400
rect 113192 34360 113732 34388
rect 111668 34348 111674 34360
rect 113726 34348 113732 34360
rect 113784 34388 113790 34400
rect 114186 34388 114192 34400
rect 113784 34360 114192 34388
rect 113784 34348 113790 34360
rect 114186 34348 114192 34360
rect 114244 34388 114250 34400
rect 115308 34388 115336 34428
rect 117406 34416 117412 34468
rect 117464 34456 117470 34468
rect 118142 34456 118148 34468
rect 117464 34428 118148 34456
rect 117464 34416 117470 34428
rect 118142 34416 118148 34428
rect 118200 34416 118206 34468
rect 114244 34360 115336 34388
rect 114244 34348 114250 34360
rect 117038 34348 117044 34400
rect 117096 34348 117102 34400
rect 1104 34298 7912 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 7912 34298
rect 1104 34224 7912 34246
rect 108008 34298 118864 34320
rect 108008 34246 112914 34298
rect 112966 34246 112978 34298
rect 113030 34246 113042 34298
rect 113094 34246 113106 34298
rect 113158 34246 113170 34298
rect 113222 34246 118864 34298
rect 108008 34224 118864 34246
rect 108850 34144 108856 34196
rect 108908 34144 108914 34196
rect 109586 34144 109592 34196
rect 109644 34184 109650 34196
rect 109957 34187 110015 34193
rect 109957 34184 109969 34187
rect 109644 34156 109969 34184
rect 109644 34144 109650 34156
rect 109957 34153 109969 34156
rect 110003 34153 110015 34187
rect 109957 34147 110015 34153
rect 110417 34187 110475 34193
rect 110417 34153 110429 34187
rect 110463 34184 110475 34187
rect 110506 34184 110512 34196
rect 110463 34156 110512 34184
rect 110463 34153 110475 34156
rect 110417 34147 110475 34153
rect 110506 34144 110512 34156
rect 110564 34144 110570 34196
rect 113450 34144 113456 34196
rect 113508 34184 113514 34196
rect 113545 34187 113603 34193
rect 113545 34184 113557 34187
rect 113508 34156 113557 34184
rect 113508 34144 113514 34156
rect 113545 34153 113557 34156
rect 113591 34153 113603 34187
rect 113545 34147 113603 34153
rect 113729 34187 113787 34193
rect 113729 34153 113741 34187
rect 113775 34153 113787 34187
rect 113729 34147 113787 34153
rect 110046 34076 110052 34128
rect 110104 34116 110110 34128
rect 110966 34116 110972 34128
rect 110104 34088 110972 34116
rect 110104 34076 110110 34088
rect 110966 34076 110972 34088
rect 111024 34116 111030 34128
rect 111429 34119 111487 34125
rect 111429 34116 111441 34119
rect 111024 34088 111441 34116
rect 111024 34076 111030 34088
rect 111429 34085 111441 34088
rect 111475 34085 111487 34119
rect 111429 34079 111487 34085
rect 112806 34076 112812 34128
rect 112864 34116 112870 34128
rect 113744 34116 113772 34147
rect 114002 34144 114008 34196
rect 114060 34184 114066 34196
rect 114278 34184 114284 34196
rect 114060 34156 114284 34184
rect 114060 34144 114066 34156
rect 114278 34144 114284 34156
rect 114336 34144 114342 34196
rect 115014 34144 115020 34196
rect 115072 34184 115078 34196
rect 115569 34187 115627 34193
rect 115569 34184 115581 34187
rect 115072 34156 115581 34184
rect 115072 34144 115078 34156
rect 115569 34153 115581 34156
rect 115615 34153 115627 34187
rect 115569 34147 115627 34153
rect 116486 34144 116492 34196
rect 116544 34184 116550 34196
rect 117225 34187 117283 34193
rect 116544 34156 117176 34184
rect 116544 34144 116550 34156
rect 117038 34116 117044 34128
rect 112864 34088 114048 34116
rect 112864 34076 112870 34088
rect 110141 34051 110199 34057
rect 108684 34020 109540 34048
rect 108482 33940 108488 33992
rect 108540 33940 108546 33992
rect 108574 33940 108580 33992
rect 108632 33980 108638 33992
rect 108684 33989 108712 34020
rect 108669 33983 108727 33989
rect 108669 33980 108681 33983
rect 108632 33952 108681 33980
rect 108632 33940 108638 33952
rect 108669 33949 108681 33952
rect 108715 33949 108727 33983
rect 108669 33943 108727 33949
rect 109034 33940 109040 33992
rect 109092 33940 109098 33992
rect 109512 33989 109540 34020
rect 110141 34017 110153 34051
rect 110187 34048 110199 34051
rect 110782 34048 110788 34060
rect 110187 34020 110788 34048
rect 110187 34017 110199 34020
rect 110141 34011 110199 34017
rect 110782 34008 110788 34020
rect 110840 34008 110846 34060
rect 111702 34048 111708 34060
rect 111628 34020 111708 34048
rect 109497 33983 109555 33989
rect 109497 33949 109509 33983
rect 109543 33949 109555 33983
rect 109497 33943 109555 33949
rect 109862 33940 109868 33992
rect 109920 33980 109926 33992
rect 109957 33983 110015 33989
rect 109957 33980 109969 33983
rect 109920 33952 109969 33980
rect 109920 33940 109926 33952
rect 109957 33949 109969 33952
rect 110003 33949 110015 33983
rect 109957 33943 110015 33949
rect 110230 33940 110236 33992
rect 110288 33940 110294 33992
rect 110414 33940 110420 33992
rect 110472 33980 110478 33992
rect 110969 33983 111027 33989
rect 110969 33980 110981 33983
rect 110472 33952 110981 33980
rect 110472 33940 110478 33952
rect 110969 33949 110981 33952
rect 111015 33949 111027 33983
rect 110969 33943 111027 33949
rect 111153 33983 111211 33989
rect 111153 33949 111165 33983
rect 111199 33980 111211 33983
rect 111334 33980 111340 33992
rect 111199 33952 111340 33980
rect 111199 33949 111211 33952
rect 111153 33943 111211 33949
rect 108758 33872 108764 33924
rect 108816 33912 108822 33924
rect 110984 33912 111012 33943
rect 111334 33940 111340 33952
rect 111392 33980 111398 33992
rect 111628 33989 111656 34020
rect 111702 34008 111708 34020
rect 111760 34008 111766 34060
rect 114020 33989 114048 34088
rect 114296 34088 117044 34116
rect 111613 33983 111671 33989
rect 111613 33980 111625 33983
rect 111392 33952 111625 33980
rect 111392 33940 111398 33952
rect 111613 33949 111625 33952
rect 111659 33949 111671 33983
rect 111613 33943 111671 33949
rect 114005 33983 114063 33989
rect 114005 33949 114017 33983
rect 114051 33980 114063 33983
rect 114186 33980 114192 33992
rect 114051 33952 114192 33980
rect 114051 33949 114063 33952
rect 114005 33943 114063 33949
rect 114186 33940 114192 33952
rect 114244 33940 114250 33992
rect 114296 33989 114324 34088
rect 117038 34076 117044 34088
rect 117096 34076 117102 34128
rect 115845 34051 115903 34057
rect 115845 34048 115857 34051
rect 115400 34020 115857 34048
rect 114281 33983 114339 33989
rect 114281 33949 114293 33983
rect 114327 33949 114339 33983
rect 114281 33943 114339 33949
rect 114922 33940 114928 33992
rect 114980 33940 114986 33992
rect 115400 33989 115428 34020
rect 115845 34017 115857 34020
rect 115891 34048 115903 34051
rect 116302 34048 116308 34060
rect 115891 34020 116308 34048
rect 115891 34017 115903 34020
rect 115845 34011 115903 34017
rect 116302 34008 116308 34020
rect 116360 34048 116366 34060
rect 117148 34048 117176 34156
rect 117225 34153 117237 34187
rect 117271 34184 117283 34187
rect 117406 34184 117412 34196
rect 117271 34156 117412 34184
rect 117271 34153 117283 34156
rect 117225 34147 117283 34153
rect 117406 34144 117412 34156
rect 117464 34144 117470 34196
rect 117682 34144 117688 34196
rect 117740 34184 117746 34196
rect 118145 34187 118203 34193
rect 118145 34184 118157 34187
rect 117740 34156 118157 34184
rect 117740 34144 117746 34156
rect 118145 34153 118157 34156
rect 118191 34153 118203 34187
rect 118145 34147 118203 34153
rect 117317 34051 117375 34057
rect 117317 34048 117329 34051
rect 116360 34020 117084 34048
rect 117148 34020 117329 34048
rect 116360 34008 116366 34020
rect 115109 33983 115167 33989
rect 115109 33949 115121 33983
rect 115155 33980 115167 33983
rect 115385 33983 115443 33989
rect 115155 33952 115336 33980
rect 115155 33949 115167 33952
rect 115109 33943 115167 33949
rect 111426 33912 111432 33924
rect 108816 33884 109356 33912
rect 110984 33884 111432 33912
rect 108816 33872 108822 33884
rect 109218 33804 109224 33856
rect 109276 33804 109282 33856
rect 109328 33853 109356 33884
rect 111426 33872 111432 33884
rect 111484 33872 111490 33924
rect 113726 33921 113732 33924
rect 111981 33915 112039 33921
rect 111981 33912 111993 33915
rect 111628 33884 111993 33912
rect 111628 33856 111656 33884
rect 111981 33881 111993 33884
rect 112027 33881 112039 33915
rect 111981 33875 112039 33881
rect 113713 33915 113732 33921
rect 113713 33881 113725 33915
rect 113713 33875 113732 33881
rect 113726 33872 113732 33875
rect 113784 33872 113790 33924
rect 113913 33915 113971 33921
rect 113913 33881 113925 33915
rect 113959 33881 113971 33915
rect 113913 33875 113971 33881
rect 115017 33915 115075 33921
rect 115017 33881 115029 33915
rect 115063 33912 115075 33915
rect 115201 33915 115259 33921
rect 115201 33912 115213 33915
rect 115063 33884 115213 33912
rect 115063 33881 115075 33884
rect 115017 33875 115075 33881
rect 115201 33881 115213 33884
rect 115247 33881 115259 33915
rect 115308 33912 115336 33952
rect 115385 33949 115397 33983
rect 115431 33949 115443 33983
rect 115385 33943 115443 33949
rect 116026 33940 116032 33992
rect 116084 33940 116090 33992
rect 116118 33940 116124 33992
rect 116176 33940 116182 33992
rect 116486 33940 116492 33992
rect 116544 33980 116550 33992
rect 117056 33989 117084 34020
rect 117317 34017 117329 34020
rect 117363 34017 117375 34051
rect 117317 34011 117375 34017
rect 117685 34051 117743 34057
rect 117685 34017 117697 34051
rect 117731 34048 117743 34051
rect 117774 34048 117780 34060
rect 117731 34020 117780 34048
rect 117731 34017 117743 34020
rect 117685 34011 117743 34017
rect 117774 34008 117780 34020
rect 117832 34008 117838 34060
rect 116581 33983 116639 33989
rect 116581 33980 116593 33983
rect 116544 33952 116593 33980
rect 116544 33940 116550 33952
rect 116581 33949 116593 33952
rect 116627 33949 116639 33983
rect 116581 33943 116639 33949
rect 116765 33983 116823 33989
rect 116765 33949 116777 33983
rect 116811 33949 116823 33983
rect 116765 33943 116823 33949
rect 117041 33983 117099 33989
rect 117041 33949 117053 33983
rect 117087 33949 117099 33983
rect 117041 33943 117099 33949
rect 117501 33983 117559 33989
rect 117501 33949 117513 33983
rect 117547 33949 117559 33983
rect 117501 33943 117559 33949
rect 116044 33912 116072 33940
rect 115308 33884 116072 33912
rect 116780 33912 116808 33943
rect 117516 33912 117544 33943
rect 117958 33940 117964 33992
rect 118016 33940 118022 33992
rect 116780 33884 117544 33912
rect 115201 33875 115259 33881
rect 109313 33847 109371 33853
rect 109313 33813 109325 33847
rect 109359 33813 109371 33847
rect 109313 33807 109371 33813
rect 110966 33804 110972 33856
rect 111024 33804 111030 33856
rect 111610 33804 111616 33856
rect 111668 33804 111674 33856
rect 111702 33804 111708 33856
rect 111760 33804 111766 33856
rect 111794 33804 111800 33856
rect 111852 33804 111858 33856
rect 113928 33844 113956 33875
rect 114189 33847 114247 33853
rect 114189 33844 114201 33847
rect 113928 33816 114201 33844
rect 114189 33813 114201 33816
rect 114235 33844 114247 33847
rect 114370 33844 114376 33856
rect 114235 33816 114376 33844
rect 114235 33813 114247 33816
rect 114189 33807 114247 33813
rect 114370 33804 114376 33816
rect 114428 33804 114434 33856
rect 115566 33804 115572 33856
rect 115624 33844 115630 33856
rect 116780 33844 116808 33884
rect 117590 33872 117596 33924
rect 117648 33912 117654 33924
rect 117777 33915 117835 33921
rect 117777 33912 117789 33915
rect 117648 33884 117789 33912
rect 117648 33872 117654 33884
rect 117777 33881 117789 33884
rect 117823 33881 117835 33915
rect 117777 33875 117835 33881
rect 115624 33816 116808 33844
rect 115624 33804 115630 33816
rect 1104 33754 7912 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 7912 33754
rect 1104 33680 7912 33702
rect 108008 33754 118864 33776
rect 108008 33702 113650 33754
rect 113702 33702 113714 33754
rect 113766 33702 113778 33754
rect 113830 33702 113842 33754
rect 113894 33702 113906 33754
rect 113958 33702 118864 33754
rect 108008 33680 118864 33702
rect 108482 33600 108488 33652
rect 108540 33640 108546 33652
rect 108577 33643 108635 33649
rect 108577 33640 108589 33643
rect 108540 33612 108589 33640
rect 108540 33600 108546 33612
rect 108577 33609 108589 33612
rect 108623 33609 108635 33643
rect 108577 33603 108635 33609
rect 109678 33600 109684 33652
rect 109736 33640 109742 33652
rect 109773 33643 109831 33649
rect 109773 33640 109785 33643
rect 109736 33612 109785 33640
rect 109736 33600 109742 33612
rect 109773 33609 109785 33612
rect 109819 33640 109831 33643
rect 110693 33643 110751 33649
rect 110693 33640 110705 33643
rect 109819 33612 110705 33640
rect 109819 33609 109831 33612
rect 109773 33603 109831 33609
rect 110693 33609 110705 33612
rect 110739 33609 110751 33643
rect 110693 33603 110751 33609
rect 110877 33643 110935 33649
rect 110877 33609 110889 33643
rect 110923 33640 110935 33643
rect 112993 33643 113051 33649
rect 110923 33612 111564 33640
rect 110923 33609 110935 33612
rect 110877 33603 110935 33609
rect 109218 33532 109224 33584
rect 109276 33572 109282 33584
rect 109589 33575 109647 33581
rect 109589 33572 109601 33575
rect 109276 33544 109601 33572
rect 109276 33532 109282 33544
rect 109589 33541 109601 33544
rect 109635 33541 109647 33575
rect 109589 33535 109647 33541
rect 110969 33575 111027 33581
rect 110969 33541 110981 33575
rect 111015 33572 111027 33575
rect 111015 33544 111472 33572
rect 111015 33541 111027 33544
rect 110969 33535 111027 33541
rect 111444 33516 111472 33544
rect 108298 33464 108304 33516
rect 108356 33464 108362 33516
rect 108666 33464 108672 33516
rect 108724 33504 108730 33516
rect 108761 33507 108819 33513
rect 108761 33504 108773 33507
rect 108724 33476 108773 33504
rect 108724 33464 108730 33476
rect 108761 33473 108773 33476
rect 108807 33473 108819 33507
rect 108761 33467 108819 33473
rect 108945 33507 109003 33513
rect 108945 33473 108957 33507
rect 108991 33504 109003 33507
rect 109126 33504 109132 33516
rect 108991 33476 109132 33504
rect 108991 33473 109003 33476
rect 108945 33467 109003 33473
rect 109126 33464 109132 33476
rect 109184 33464 109190 33516
rect 109770 33464 109776 33516
rect 109828 33504 109834 33516
rect 109865 33507 109923 33513
rect 109865 33504 109877 33507
rect 109828 33476 109877 33504
rect 109828 33464 109834 33476
rect 109865 33473 109877 33476
rect 109911 33504 109923 33507
rect 111061 33507 111119 33513
rect 109911 33476 110828 33504
rect 109911 33473 109923 33476
rect 109865 33467 109923 33473
rect 110598 33396 110604 33448
rect 110656 33436 110662 33448
rect 110693 33439 110751 33445
rect 110693 33436 110705 33439
rect 110656 33408 110705 33436
rect 110656 33396 110662 33408
rect 110693 33405 110705 33408
rect 110739 33405 110751 33439
rect 110800 33436 110828 33476
rect 111061 33473 111073 33507
rect 111107 33504 111119 33507
rect 111334 33504 111340 33516
rect 111107 33476 111340 33504
rect 111107 33473 111119 33476
rect 111061 33467 111119 33473
rect 111334 33464 111340 33476
rect 111392 33464 111398 33516
rect 111426 33464 111432 33516
rect 111484 33464 111490 33516
rect 111536 33513 111564 33612
rect 112993 33609 113005 33643
rect 113039 33640 113051 33643
rect 113821 33643 113879 33649
rect 113821 33640 113833 33643
rect 113039 33612 113833 33640
rect 113039 33609 113051 33612
rect 112993 33603 113051 33609
rect 113821 33609 113833 33612
rect 113867 33609 113879 33643
rect 113821 33603 113879 33609
rect 114189 33643 114247 33649
rect 114189 33609 114201 33643
rect 114235 33609 114247 33643
rect 114189 33603 114247 33609
rect 114833 33643 114891 33649
rect 114833 33609 114845 33643
rect 114879 33640 114891 33643
rect 115106 33640 115112 33652
rect 114879 33612 115112 33640
rect 114879 33609 114891 33612
rect 114833 33603 114891 33609
rect 114204 33572 114232 33603
rect 115106 33600 115112 33612
rect 115164 33600 115170 33652
rect 115198 33600 115204 33652
rect 115256 33640 115262 33652
rect 115385 33643 115443 33649
rect 115385 33640 115397 33643
rect 115256 33612 115397 33640
rect 115256 33600 115262 33612
rect 115385 33609 115397 33612
rect 115431 33609 115443 33643
rect 115385 33603 115443 33609
rect 115566 33600 115572 33652
rect 115624 33600 115630 33652
rect 116302 33640 116308 33652
rect 115676 33612 116308 33640
rect 115676 33572 115704 33612
rect 116302 33600 116308 33612
rect 116360 33640 116366 33652
rect 116360 33612 116532 33640
rect 116360 33600 116366 33612
rect 112272 33544 112760 33572
rect 114204 33544 115704 33572
rect 111521 33507 111579 33513
rect 111521 33473 111533 33507
rect 111567 33504 111579 33507
rect 111794 33504 111800 33516
rect 111567 33476 111800 33504
rect 111567 33473 111579 33476
rect 111521 33467 111579 33473
rect 111153 33439 111211 33445
rect 111153 33436 111165 33439
rect 110800 33408 111165 33436
rect 110693 33399 110751 33405
rect 111153 33405 111165 33408
rect 111199 33405 111211 33439
rect 111153 33399 111211 33405
rect 109586 33328 109592 33380
rect 109644 33328 109650 33380
rect 110708 33368 110736 33399
rect 111610 33396 111616 33448
rect 111668 33396 111674 33448
rect 111628 33368 111656 33396
rect 110708 33340 111656 33368
rect 108485 33303 108543 33309
rect 108485 33269 108497 33303
rect 108531 33300 108543 33303
rect 108942 33300 108948 33312
rect 108531 33272 108948 33300
rect 108531 33269 108543 33272
rect 108485 33263 108543 33269
rect 108942 33260 108948 33272
rect 109000 33260 109006 33312
rect 109221 33303 109279 33309
rect 109221 33269 109233 33303
rect 109267 33300 109279 33303
rect 109402 33300 109408 33312
rect 109267 33272 109408 33300
rect 109267 33269 109279 33272
rect 109221 33263 109279 33269
rect 109402 33260 109408 33272
rect 109460 33260 109466 33312
rect 111720 33300 111748 33476
rect 111794 33464 111800 33476
rect 111852 33464 111858 33516
rect 111978 33464 111984 33516
rect 112036 33464 112042 33516
rect 112073 33439 112131 33445
rect 112073 33405 112085 33439
rect 112119 33436 112131 33439
rect 112272 33436 112300 33544
rect 112732 33516 112760 33544
rect 115750 33532 115756 33584
rect 115808 33581 115814 33584
rect 115808 33575 115871 33581
rect 115808 33541 115825 33575
rect 115859 33541 115871 33575
rect 115808 33535 115871 33541
rect 116029 33575 116087 33581
rect 116029 33541 116041 33575
rect 116075 33572 116087 33575
rect 116210 33572 116216 33584
rect 116075 33544 116216 33572
rect 116075 33541 116087 33544
rect 116029 33535 116087 33541
rect 115808 33532 115814 33535
rect 116210 33532 116216 33544
rect 116268 33532 116274 33584
rect 112622 33464 112628 33516
rect 112680 33464 112686 33516
rect 112714 33464 112720 33516
rect 112772 33504 112778 33516
rect 113729 33507 113787 33513
rect 113729 33504 113741 33507
rect 112772 33476 113741 33504
rect 112772 33464 112778 33476
rect 113729 33473 113741 33476
rect 113775 33473 113787 33507
rect 113729 33467 113787 33473
rect 114554 33464 114560 33516
rect 114612 33504 114618 33516
rect 114649 33507 114707 33513
rect 114649 33504 114661 33507
rect 114612 33476 114661 33504
rect 114612 33464 114618 33476
rect 114649 33473 114661 33476
rect 114695 33473 114707 33507
rect 114649 33467 114707 33473
rect 114830 33464 114836 33516
rect 114888 33464 114894 33516
rect 115444 33507 115502 33513
rect 115444 33473 115456 33507
rect 115490 33504 115502 33507
rect 115658 33504 115664 33516
rect 115490 33476 115664 33504
rect 115490 33473 115502 33476
rect 115444 33467 115502 33473
rect 115658 33464 115664 33476
rect 115716 33464 115722 33516
rect 116397 33507 116455 33513
rect 116397 33473 116409 33507
rect 116443 33473 116455 33507
rect 116504 33504 116532 33612
rect 117498 33600 117504 33652
rect 117556 33640 117562 33652
rect 117685 33643 117743 33649
rect 117685 33640 117697 33643
rect 117556 33612 117697 33640
rect 117556 33600 117562 33612
rect 117685 33609 117697 33612
rect 117731 33609 117743 33643
rect 117685 33603 117743 33609
rect 116581 33507 116639 33513
rect 116581 33504 116593 33507
rect 116504 33476 116593 33504
rect 116397 33467 116455 33473
rect 116581 33473 116593 33476
rect 116627 33504 116639 33507
rect 117317 33507 117375 33513
rect 117317 33504 117329 33507
rect 116627 33476 117329 33504
rect 116627 33473 116639 33476
rect 116581 33467 116639 33473
rect 117317 33473 117329 33476
rect 117363 33473 117375 33507
rect 117317 33467 117375 33473
rect 112533 33439 112591 33445
rect 112533 33436 112545 33439
rect 112119 33408 112300 33436
rect 112364 33408 112545 33436
rect 112119 33405 112131 33408
rect 112073 33399 112131 33405
rect 112364 33377 112392 33408
rect 112533 33405 112545 33408
rect 112579 33405 112591 33439
rect 112533 33399 112591 33405
rect 113637 33439 113695 33445
rect 113637 33405 113649 33439
rect 113683 33436 113695 33439
rect 114002 33436 114008 33448
rect 113683 33408 114008 33436
rect 113683 33405 113695 33408
rect 113637 33399 113695 33405
rect 112349 33371 112407 33377
rect 112349 33337 112361 33371
rect 112395 33337 112407 33371
rect 112349 33331 112407 33337
rect 113652 33300 113680 33399
rect 114002 33396 114008 33408
rect 114060 33436 114066 33448
rect 114925 33439 114983 33445
rect 114925 33436 114937 33439
rect 114060 33408 114937 33436
rect 114060 33396 114066 33408
rect 114925 33405 114937 33408
rect 114971 33405 114983 33439
rect 114925 33399 114983 33405
rect 115017 33439 115075 33445
rect 115017 33405 115029 33439
rect 115063 33436 115075 33439
rect 116026 33436 116032 33448
rect 115063 33408 116032 33436
rect 115063 33405 115075 33408
rect 115017 33399 115075 33405
rect 116026 33396 116032 33408
rect 116084 33396 116090 33448
rect 116118 33396 116124 33448
rect 116176 33436 116182 33448
rect 116412 33436 116440 33467
rect 116176 33408 116532 33436
rect 116176 33396 116182 33408
rect 115474 33328 115480 33380
rect 115532 33368 115538 33380
rect 116504 33368 116532 33408
rect 117130 33396 117136 33448
rect 117188 33396 117194 33448
rect 117225 33439 117283 33445
rect 117225 33405 117237 33439
rect 117271 33436 117283 33439
rect 117682 33436 117688 33448
rect 117271 33408 117688 33436
rect 117271 33405 117283 33408
rect 117225 33399 117283 33405
rect 117682 33396 117688 33408
rect 117740 33396 117746 33448
rect 116670 33368 116676 33380
rect 115532 33340 115888 33368
rect 116504 33340 116676 33368
rect 115532 33328 115538 33340
rect 111720 33272 113680 33300
rect 115382 33260 115388 33312
rect 115440 33300 115446 33312
rect 115860 33309 115888 33340
rect 116670 33328 116676 33340
rect 116728 33368 116734 33380
rect 117958 33368 117964 33380
rect 116728 33340 117964 33368
rect 116728 33328 116734 33340
rect 117958 33328 117964 33340
rect 118016 33328 118022 33380
rect 115661 33303 115719 33309
rect 115661 33300 115673 33303
rect 115440 33272 115673 33300
rect 115440 33260 115446 33272
rect 115661 33269 115673 33272
rect 115707 33269 115719 33303
rect 115661 33263 115719 33269
rect 115845 33303 115903 33309
rect 115845 33269 115857 33303
rect 115891 33269 115903 33303
rect 115845 33263 115903 33269
rect 116581 33303 116639 33309
rect 116581 33269 116593 33303
rect 116627 33300 116639 33303
rect 116946 33300 116952 33312
rect 116627 33272 116952 33300
rect 116627 33269 116639 33272
rect 116581 33263 116639 33269
rect 116946 33260 116952 33272
rect 117004 33300 117010 33312
rect 117774 33300 117780 33312
rect 117004 33272 117780 33300
rect 117004 33260 117010 33272
rect 117774 33260 117780 33272
rect 117832 33260 117838 33312
rect 1104 33210 7912 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 7912 33210
rect 1104 33136 7912 33158
rect 108008 33210 118864 33232
rect 108008 33158 112914 33210
rect 112966 33158 112978 33210
rect 113030 33158 113042 33210
rect 113094 33158 113106 33210
rect 113158 33158 113170 33210
rect 113222 33158 118864 33210
rect 108008 33136 118864 33158
rect 108761 33099 108819 33105
rect 108761 33065 108773 33099
rect 108807 33096 108819 33099
rect 108850 33096 108856 33108
rect 108807 33068 108856 33096
rect 108807 33065 108819 33068
rect 108761 33059 108819 33065
rect 108850 33056 108856 33068
rect 108908 33056 108914 33108
rect 109037 33099 109095 33105
rect 109037 33065 109049 33099
rect 109083 33096 109095 33099
rect 109126 33096 109132 33108
rect 109083 33068 109132 33096
rect 109083 33065 109095 33068
rect 109037 33059 109095 33065
rect 109126 33056 109132 33068
rect 109184 33056 109190 33108
rect 109678 33056 109684 33108
rect 109736 33056 109742 33108
rect 109865 33099 109923 33105
rect 109865 33065 109877 33099
rect 109911 33096 109923 33099
rect 110230 33096 110236 33108
rect 109911 33068 110236 33096
rect 109911 33065 109923 33068
rect 109865 33059 109923 33065
rect 110230 33056 110236 33068
rect 110288 33056 110294 33108
rect 114554 33056 114560 33108
rect 114612 33096 114618 33108
rect 115198 33096 115204 33108
rect 114612 33068 115204 33096
rect 114612 33056 114618 33068
rect 115198 33056 115204 33068
rect 115256 33056 115262 33108
rect 116026 33056 116032 33108
rect 116084 33096 116090 33108
rect 116397 33099 116455 33105
rect 116397 33096 116409 33099
rect 116084 33068 116409 33096
rect 116084 33056 116090 33068
rect 116397 33065 116409 33068
rect 116443 33065 116455 33099
rect 116397 33059 116455 33065
rect 116670 33056 116676 33108
rect 116728 33056 116734 33108
rect 117590 33056 117596 33108
rect 117648 33056 117654 33108
rect 117682 33056 117688 33108
rect 117740 33056 117746 33108
rect 108298 32988 108304 33040
rect 108356 32988 108362 33040
rect 110046 32988 110052 33040
rect 110104 33028 110110 33040
rect 111978 33028 111984 33040
rect 110104 33000 111984 33028
rect 110104 32988 110110 33000
rect 111978 32988 111984 33000
rect 112036 32988 112042 33040
rect 115216 33028 115244 33056
rect 117130 33028 117136 33040
rect 115216 33000 117136 33028
rect 108316 32960 108344 32988
rect 110233 32963 110291 32969
rect 108316 32932 108620 32960
rect 108298 32852 108304 32904
rect 108356 32852 108362 32904
rect 108592 32901 108620 32932
rect 110233 32929 110245 32963
rect 110279 32960 110291 32963
rect 110966 32960 110972 32972
rect 110279 32932 110972 32960
rect 110279 32929 110291 32932
rect 110233 32923 110291 32929
rect 110966 32920 110972 32932
rect 111024 32920 111030 32972
rect 111610 32920 111616 32972
rect 111668 32960 111674 32972
rect 115750 32960 115756 32972
rect 111668 32932 113220 32960
rect 111668 32920 111674 32932
rect 108577 32895 108635 32901
rect 108577 32861 108589 32895
rect 108623 32861 108635 32895
rect 108577 32855 108635 32861
rect 109218 32852 109224 32904
rect 109276 32892 109282 32904
rect 110325 32895 110383 32901
rect 109276 32864 109540 32892
rect 109276 32852 109282 32864
rect 109512 32833 109540 32864
rect 110325 32861 110337 32895
rect 110371 32892 110383 32895
rect 111794 32892 111800 32904
rect 110371 32864 111800 32892
rect 110371 32861 110383 32864
rect 110325 32855 110383 32861
rect 111794 32852 111800 32864
rect 111852 32852 111858 32904
rect 112714 32852 112720 32904
rect 112772 32852 112778 32904
rect 113192 32901 113220 32932
rect 115676 32932 115756 32960
rect 112901 32895 112959 32901
rect 112901 32861 112913 32895
rect 112947 32861 112959 32895
rect 112901 32855 112959 32861
rect 113177 32895 113235 32901
rect 113177 32861 113189 32895
rect 113223 32861 113235 32895
rect 113177 32855 113235 32861
rect 109770 32833 109776 32836
rect 108393 32827 108451 32833
rect 108393 32824 108405 32827
rect 107948 32796 108405 32824
rect 1104 32666 7912 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 7912 32666
rect 1104 32592 7912 32614
rect 107948 32484 107976 32796
rect 108393 32793 108405 32796
rect 108439 32824 108451 32827
rect 109497 32827 109555 32833
rect 108439 32796 109034 32824
rect 108439 32793 108451 32796
rect 108393 32787 108451 32793
rect 109006 32756 109034 32796
rect 109497 32793 109509 32827
rect 109543 32793 109555 32827
rect 109497 32787 109555 32793
rect 109713 32827 109776 32833
rect 109713 32793 109725 32827
rect 109759 32793 109776 32827
rect 109713 32787 109776 32793
rect 109770 32784 109776 32787
rect 109828 32784 109834 32836
rect 112530 32784 112536 32836
rect 112588 32824 112594 32836
rect 112916 32824 112944 32855
rect 115014 32852 115020 32904
rect 115072 32892 115078 32904
rect 115676 32901 115704 32932
rect 115750 32920 115756 32932
rect 115808 32960 115814 32972
rect 117056 32969 117084 33000
rect 117130 32988 117136 33000
rect 117188 32988 117194 33040
rect 117041 32963 117099 32969
rect 115808 32932 116256 32960
rect 115808 32920 115814 32932
rect 116228 32904 116256 32932
rect 117041 32929 117053 32963
rect 117087 32929 117099 32963
rect 117041 32923 117099 32929
rect 118142 32920 118148 32972
rect 118200 32920 118206 32972
rect 115385 32895 115443 32901
rect 115385 32892 115397 32895
rect 115072 32864 115397 32892
rect 115072 32852 115078 32864
rect 115385 32861 115397 32864
rect 115431 32861 115443 32895
rect 115385 32855 115443 32861
rect 115661 32895 115719 32901
rect 115661 32861 115673 32895
rect 115707 32861 115719 32895
rect 115661 32855 115719 32861
rect 112990 32824 112996 32836
rect 112588 32796 112996 32824
rect 112588 32784 112594 32796
rect 112990 32784 112996 32796
rect 113048 32824 113054 32836
rect 115290 32824 115296 32836
rect 113048 32796 115296 32824
rect 113048 32784 113054 32796
rect 115290 32784 115296 32796
rect 115348 32784 115354 32836
rect 115400 32824 115428 32855
rect 115842 32852 115848 32904
rect 115900 32852 115906 32904
rect 115934 32852 115940 32904
rect 115992 32852 115998 32904
rect 116121 32895 116179 32901
rect 116121 32892 116133 32895
rect 116044 32864 116133 32892
rect 115860 32824 115888 32852
rect 115400 32796 115888 32824
rect 109402 32756 109408 32768
rect 109006 32728 109408 32756
rect 109402 32716 109408 32728
rect 109460 32716 109466 32768
rect 109862 32716 109868 32768
rect 109920 32756 109926 32768
rect 109957 32759 110015 32765
rect 109957 32756 109969 32759
rect 109920 32728 109969 32756
rect 109920 32716 109926 32728
rect 109957 32725 109969 32728
rect 110003 32725 110015 32759
rect 109957 32719 110015 32725
rect 112901 32759 112959 32765
rect 112901 32725 112913 32759
rect 112947 32756 112959 32759
rect 113174 32756 113180 32768
rect 112947 32728 113180 32756
rect 112947 32725 112959 32728
rect 112901 32719 112959 32725
rect 113174 32716 113180 32728
rect 113232 32716 113238 32768
rect 113269 32759 113327 32765
rect 113269 32725 113281 32759
rect 113315 32756 113327 32759
rect 114278 32756 114284 32768
rect 113315 32728 114284 32756
rect 113315 32725 113327 32728
rect 113269 32719 113327 32725
rect 114278 32716 114284 32728
rect 114336 32716 114342 32768
rect 115474 32716 115480 32768
rect 115532 32756 115538 32768
rect 115569 32759 115627 32765
rect 115569 32756 115581 32759
rect 115532 32728 115581 32756
rect 115532 32716 115538 32728
rect 115569 32725 115581 32728
rect 115615 32756 115627 32759
rect 115842 32756 115848 32768
rect 115615 32728 115848 32756
rect 115615 32725 115627 32728
rect 115569 32719 115627 32725
rect 115842 32716 115848 32728
rect 115900 32756 115906 32768
rect 116044 32756 116072 32864
rect 116121 32861 116133 32864
rect 116167 32861 116179 32895
rect 116121 32855 116179 32861
rect 116210 32852 116216 32904
rect 116268 32852 116274 32904
rect 116394 32852 116400 32904
rect 116452 32892 116458 32904
rect 116489 32895 116547 32901
rect 116489 32892 116501 32895
rect 116452 32864 116501 32892
rect 116452 32852 116458 32864
rect 116489 32861 116501 32864
rect 116535 32861 116547 32895
rect 116489 32855 116547 32861
rect 117682 32852 117688 32904
rect 117740 32892 117746 32904
rect 118053 32895 118111 32901
rect 118053 32892 118065 32895
rect 117740 32864 118065 32892
rect 117740 32852 117746 32864
rect 118053 32861 118065 32864
rect 118099 32861 118111 32895
rect 118053 32855 118111 32861
rect 115900 32728 116072 32756
rect 115900 32716 115906 32728
rect 117130 32716 117136 32768
rect 117188 32716 117194 32768
rect 117222 32716 117228 32768
rect 117280 32716 117286 32768
rect 108008 32666 118864 32688
rect 108008 32614 113650 32666
rect 113702 32614 113714 32666
rect 113766 32614 113778 32666
rect 113830 32614 113842 32666
rect 113894 32614 113906 32666
rect 113958 32614 118864 32666
rect 108008 32592 118864 32614
rect 108390 32512 108396 32564
rect 108448 32552 108454 32564
rect 108501 32555 108559 32561
rect 108501 32552 108513 32555
rect 108448 32524 108513 32552
rect 108448 32512 108454 32524
rect 108501 32521 108513 32524
rect 108547 32521 108559 32555
rect 108501 32515 108559 32521
rect 108666 32512 108672 32564
rect 108724 32512 108730 32564
rect 109313 32555 109371 32561
rect 109313 32521 109325 32555
rect 109359 32552 109371 32555
rect 110138 32552 110144 32564
rect 109359 32524 110144 32552
rect 109359 32521 109371 32524
rect 109313 32515 109371 32521
rect 110138 32512 110144 32524
rect 110196 32512 110202 32564
rect 112622 32512 112628 32564
rect 112680 32512 112686 32564
rect 114281 32555 114339 32561
rect 114281 32521 114293 32555
rect 114327 32552 114339 32555
rect 114462 32552 114468 32564
rect 114327 32524 114468 32552
rect 114327 32521 114339 32524
rect 114281 32515 114339 32521
rect 114462 32512 114468 32524
rect 114520 32512 114526 32564
rect 115658 32512 115664 32564
rect 115716 32512 115722 32564
rect 116118 32512 116124 32564
rect 116176 32512 116182 32564
rect 116210 32512 116216 32564
rect 116268 32552 116274 32564
rect 116581 32555 116639 32561
rect 116581 32552 116593 32555
rect 116268 32524 116593 32552
rect 116268 32512 116274 32524
rect 116581 32521 116593 32524
rect 116627 32521 116639 32555
rect 116581 32515 116639 32521
rect 117317 32555 117375 32561
rect 117317 32521 117329 32555
rect 117363 32552 117375 32555
rect 117590 32552 117596 32564
rect 117363 32524 117596 32552
rect 117363 32521 117375 32524
rect 117317 32515 117375 32521
rect 117590 32512 117596 32524
rect 117648 32512 117654 32564
rect 117682 32512 117688 32564
rect 117740 32512 117746 32564
rect 118142 32512 118148 32564
rect 118200 32512 118206 32564
rect 108301 32487 108359 32493
rect 108301 32484 108313 32487
rect 107948 32456 108313 32484
rect 108301 32453 108313 32456
rect 108347 32453 108359 32487
rect 112640 32484 112668 32512
rect 116136 32484 116164 32512
rect 108301 32447 108359 32453
rect 109006 32456 110000 32484
rect 109006 32428 109034 32456
rect 108942 32376 108948 32428
rect 109000 32388 109034 32428
rect 109000 32376 109006 32388
rect 109494 32376 109500 32428
rect 109552 32416 109558 32428
rect 109972 32425 110000 32456
rect 112180 32456 113312 32484
rect 112180 32428 112208 32456
rect 109589 32419 109647 32425
rect 109589 32416 109601 32419
rect 109552 32388 109601 32416
rect 109552 32376 109558 32388
rect 109589 32385 109601 32388
rect 109635 32385 109647 32419
rect 109589 32379 109647 32385
rect 109957 32419 110015 32425
rect 109957 32385 109969 32419
rect 110003 32385 110015 32419
rect 109957 32379 110015 32385
rect 110966 32376 110972 32428
rect 111024 32376 111030 32428
rect 111153 32419 111211 32425
rect 111153 32385 111165 32419
rect 111199 32416 111211 32419
rect 111426 32416 111432 32428
rect 111199 32388 111432 32416
rect 111199 32385 111211 32388
rect 111153 32379 111211 32385
rect 111426 32376 111432 32388
rect 111484 32376 111490 32428
rect 111613 32419 111671 32425
rect 111613 32385 111625 32419
rect 111659 32385 111671 32419
rect 111613 32379 111671 32385
rect 111889 32419 111947 32425
rect 111889 32385 111901 32419
rect 111935 32385 111947 32419
rect 111889 32379 111947 32385
rect 109037 32351 109095 32357
rect 109037 32317 109049 32351
rect 109083 32348 109095 32351
rect 109862 32348 109868 32360
rect 109083 32320 109868 32348
rect 109083 32317 109095 32320
rect 109037 32311 109095 32317
rect 109862 32308 109868 32320
rect 109920 32308 109926 32360
rect 111334 32308 111340 32360
rect 111392 32348 111398 32360
rect 111628 32348 111656 32379
rect 111392 32320 111656 32348
rect 111392 32308 111398 32320
rect 109773 32283 109831 32289
rect 109773 32280 109785 32283
rect 108500 32252 109785 32280
rect 108500 32224 108528 32252
rect 109773 32249 109785 32252
rect 109819 32249 109831 32283
rect 109773 32243 109831 32249
rect 108482 32172 108488 32224
rect 108540 32172 108546 32224
rect 109402 32172 109408 32224
rect 109460 32212 109466 32224
rect 109497 32215 109555 32221
rect 109497 32212 109509 32215
rect 109460 32184 109509 32212
rect 109460 32172 109466 32184
rect 109497 32181 109509 32184
rect 109543 32212 109555 32215
rect 110049 32215 110107 32221
rect 110049 32212 110061 32215
rect 109543 32184 110061 32212
rect 109543 32181 109555 32184
rect 109497 32175 109555 32181
rect 110049 32181 110061 32184
rect 110095 32181 110107 32215
rect 110049 32175 110107 32181
rect 110874 32172 110880 32224
rect 110932 32212 110938 32224
rect 111337 32215 111395 32221
rect 111337 32212 111349 32215
rect 110932 32184 111349 32212
rect 110932 32172 110938 32184
rect 111337 32181 111349 32184
rect 111383 32181 111395 32215
rect 111337 32175 111395 32181
rect 111797 32215 111855 32221
rect 111797 32181 111809 32215
rect 111843 32212 111855 32215
rect 111904 32212 111932 32379
rect 112162 32376 112168 32428
rect 112220 32376 112226 32428
rect 112714 32416 112720 32428
rect 112272 32388 112720 32416
rect 112070 32308 112076 32360
rect 112128 32348 112134 32360
rect 112272 32348 112300 32388
rect 112714 32376 112720 32388
rect 112772 32376 112778 32428
rect 112901 32419 112959 32425
rect 112901 32385 112913 32419
rect 112947 32416 112959 32419
rect 112990 32416 112996 32428
rect 112947 32388 112996 32416
rect 112947 32385 112959 32388
rect 112901 32379 112959 32385
rect 112990 32376 112996 32388
rect 113048 32376 113054 32428
rect 113284 32425 113312 32456
rect 116044 32456 116164 32484
rect 116412 32456 116808 32484
rect 113269 32419 113327 32425
rect 113269 32385 113281 32419
rect 113315 32385 113327 32419
rect 113269 32379 113327 32385
rect 113362 32419 113420 32425
rect 113362 32385 113374 32419
rect 113408 32385 113420 32419
rect 113362 32379 113420 32385
rect 112128 32320 112300 32348
rect 112128 32308 112134 32320
rect 112438 32308 112444 32360
rect 112496 32348 112502 32360
rect 113376 32348 113404 32379
rect 114278 32376 114284 32428
rect 114336 32416 114342 32428
rect 114833 32419 114891 32425
rect 114336 32388 114381 32416
rect 114336 32376 114342 32388
rect 114833 32385 114845 32419
rect 114879 32385 114891 32419
rect 114833 32379 114891 32385
rect 115293 32419 115351 32425
rect 115293 32385 115305 32419
rect 115339 32385 115351 32419
rect 115293 32379 115351 32385
rect 112496 32320 113404 32348
rect 113637 32351 113695 32357
rect 112496 32308 112502 32320
rect 113637 32317 113649 32351
rect 113683 32348 113695 32351
rect 113821 32351 113879 32357
rect 113821 32348 113833 32351
rect 113683 32320 113833 32348
rect 113683 32317 113695 32320
rect 113637 32311 113695 32317
rect 113821 32317 113833 32320
rect 113867 32317 113879 32351
rect 114848 32348 114876 32379
rect 115198 32348 115204 32360
rect 113821 32311 113879 32317
rect 114388 32320 115204 32348
rect 112625 32283 112683 32289
rect 112625 32249 112637 32283
rect 112671 32280 112683 32283
rect 113450 32280 113456 32292
rect 112671 32252 113456 32280
rect 112671 32249 112683 32252
rect 112625 32243 112683 32249
rect 113450 32240 113456 32252
rect 113508 32240 113514 32292
rect 114186 32280 114192 32292
rect 113836 32252 114192 32280
rect 111978 32212 111984 32224
rect 111843 32184 111984 32212
rect 111843 32181 111855 32184
rect 111797 32175 111855 32181
rect 111978 32172 111984 32184
rect 112036 32172 112042 32224
rect 112073 32215 112131 32221
rect 112073 32181 112085 32215
rect 112119 32212 112131 32215
rect 112254 32212 112260 32224
rect 112119 32184 112260 32212
rect 112119 32181 112131 32184
rect 112073 32175 112131 32181
rect 112254 32172 112260 32184
rect 112312 32172 112318 32224
rect 112346 32172 112352 32224
rect 112404 32212 112410 32224
rect 113836 32212 113864 32252
rect 114186 32240 114192 32252
rect 114244 32280 114250 32292
rect 114388 32280 114416 32320
rect 115198 32308 115204 32320
rect 115256 32308 115262 32360
rect 115308 32348 115336 32379
rect 115382 32376 115388 32428
rect 115440 32416 115446 32428
rect 115569 32419 115627 32425
rect 115569 32416 115581 32419
rect 115440 32388 115581 32416
rect 115440 32376 115446 32388
rect 115569 32385 115581 32388
rect 115615 32385 115627 32419
rect 115569 32379 115627 32385
rect 115753 32419 115811 32425
rect 115753 32385 115765 32419
rect 115799 32385 115811 32419
rect 115753 32379 115811 32385
rect 115937 32419 115995 32425
rect 115937 32385 115949 32419
rect 115983 32416 115995 32419
rect 116044 32416 116072 32456
rect 115983 32388 116072 32416
rect 116121 32419 116179 32425
rect 115983 32385 115995 32388
rect 115937 32379 115995 32385
rect 116121 32385 116133 32419
rect 116167 32416 116179 32419
rect 116302 32416 116308 32428
rect 116167 32388 116308 32416
rect 116167 32385 116179 32388
rect 116121 32379 116179 32385
rect 115474 32348 115480 32360
rect 115308 32320 115480 32348
rect 115474 32308 115480 32320
rect 115532 32348 115538 32360
rect 115768 32348 115796 32379
rect 116302 32376 116308 32388
rect 116360 32376 116366 32428
rect 115532 32320 115796 32348
rect 115532 32308 115538 32320
rect 115842 32308 115848 32360
rect 115900 32348 115906 32360
rect 115900 32320 116072 32348
rect 115900 32308 115906 32320
rect 114244 32252 114416 32280
rect 114465 32283 114523 32289
rect 114244 32240 114250 32252
rect 114465 32249 114477 32283
rect 114511 32280 114523 32283
rect 115934 32280 115940 32292
rect 114511 32252 115940 32280
rect 114511 32249 114523 32252
rect 114465 32243 114523 32249
rect 115934 32240 115940 32252
rect 115992 32240 115998 32292
rect 116044 32289 116072 32320
rect 116210 32308 116216 32360
rect 116268 32348 116274 32360
rect 116412 32348 116440 32456
rect 116780 32428 116808 32456
rect 116489 32419 116547 32425
rect 116489 32385 116501 32419
rect 116535 32385 116547 32419
rect 116489 32379 116547 32385
rect 116268 32320 116440 32348
rect 116268 32308 116274 32320
rect 116029 32283 116087 32289
rect 116029 32249 116041 32283
rect 116075 32280 116087 32283
rect 116504 32280 116532 32379
rect 116762 32376 116768 32428
rect 116820 32376 116826 32428
rect 116854 32376 116860 32428
rect 116912 32376 116918 32428
rect 116946 32376 116952 32428
rect 117004 32425 117010 32428
rect 117004 32419 117058 32425
rect 117004 32385 117012 32419
rect 117046 32385 117058 32419
rect 117004 32379 117058 32385
rect 117133 32419 117191 32425
rect 117133 32385 117145 32419
rect 117179 32385 117191 32419
rect 117133 32379 117191 32385
rect 117225 32422 117283 32425
rect 117314 32422 117320 32428
rect 117225 32419 117320 32422
rect 117225 32385 117237 32419
rect 117271 32394 117320 32419
rect 117271 32385 117283 32394
rect 117225 32379 117283 32385
rect 117004 32376 117010 32379
rect 116578 32308 116584 32360
rect 116636 32348 116642 32360
rect 117147 32348 117175 32379
rect 117314 32376 117320 32394
rect 117372 32376 117378 32428
rect 117498 32376 117504 32428
rect 117556 32376 117562 32428
rect 117774 32376 117780 32428
rect 117832 32376 117838 32428
rect 117870 32419 117928 32425
rect 117870 32385 117882 32419
rect 117916 32385 117928 32419
rect 117870 32379 117928 32385
rect 116636 32320 117175 32348
rect 116636 32308 116642 32320
rect 117406 32280 117412 32292
rect 116075 32252 116440 32280
rect 116504 32252 117412 32280
rect 116075 32249 116087 32252
rect 116029 32243 116087 32249
rect 112404 32184 113864 32212
rect 112404 32172 112410 32184
rect 113910 32172 113916 32224
rect 113968 32172 113974 32224
rect 114922 32172 114928 32224
rect 114980 32212 114986 32224
rect 115106 32212 115112 32224
rect 114980 32184 115112 32212
rect 114980 32172 114986 32184
rect 115106 32172 115112 32184
rect 115164 32172 115170 32224
rect 115477 32215 115535 32221
rect 115477 32181 115489 32215
rect 115523 32212 115535 32215
rect 116210 32212 116216 32224
rect 115523 32184 116216 32212
rect 115523 32181 115535 32184
rect 115477 32175 115535 32181
rect 116210 32172 116216 32184
rect 116268 32172 116274 32224
rect 116302 32172 116308 32224
rect 116360 32172 116366 32224
rect 116412 32212 116440 32252
rect 117406 32240 117412 32252
rect 117464 32240 117470 32292
rect 117884 32212 117912 32379
rect 116412 32184 117912 32212
rect 1104 32122 7912 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 7912 32122
rect 1104 32048 7912 32070
rect 108008 32122 118864 32144
rect 108008 32070 112914 32122
rect 112966 32070 112978 32122
rect 113030 32070 113042 32122
rect 113094 32070 113106 32122
rect 113158 32070 113170 32122
rect 113222 32070 118864 32122
rect 108008 32048 118864 32070
rect 109497 32011 109555 32017
rect 109497 32008 109509 32011
rect 109006 31980 109509 32008
rect 109006 31940 109034 31980
rect 109497 31977 109509 31980
rect 109543 31977 109555 32011
rect 109497 31971 109555 31977
rect 111521 32011 111579 32017
rect 111521 31977 111533 32011
rect 111567 32008 111579 32011
rect 112070 32008 112076 32020
rect 111567 31980 112076 32008
rect 111567 31977 111579 31980
rect 111521 31971 111579 31977
rect 112070 31968 112076 31980
rect 112128 31968 112134 32020
rect 115382 31968 115388 32020
rect 115440 31968 115446 32020
rect 115474 31968 115480 32020
rect 115532 31968 115538 32020
rect 116026 32008 116032 32020
rect 115584 31980 116032 32008
rect 108960 31912 109034 31940
rect 109221 31943 109279 31949
rect 108758 31832 108764 31884
rect 108816 31872 108822 31884
rect 108960 31881 108988 31912
rect 109221 31909 109233 31943
rect 109267 31940 109279 31943
rect 110322 31940 110328 31952
rect 109267 31912 110328 31940
rect 109267 31909 109279 31912
rect 109221 31903 109279 31909
rect 110322 31900 110328 31912
rect 110380 31900 110386 31952
rect 110598 31900 110604 31952
rect 110656 31940 110662 31952
rect 110969 31943 111027 31949
rect 110969 31940 110981 31943
rect 110656 31912 110981 31940
rect 110656 31900 110662 31912
rect 110969 31909 110981 31912
rect 111015 31940 111027 31943
rect 111702 31940 111708 31952
rect 111015 31912 111708 31940
rect 111015 31909 111027 31912
rect 110969 31903 111027 31909
rect 111702 31900 111708 31912
rect 111760 31900 111766 31952
rect 112717 31943 112775 31949
rect 112717 31909 112729 31943
rect 112763 31940 112775 31943
rect 113174 31940 113180 31952
rect 112763 31912 113180 31940
rect 112763 31909 112775 31912
rect 112717 31903 112775 31909
rect 113174 31900 113180 31912
rect 113232 31900 113238 31952
rect 114094 31900 114100 31952
rect 114152 31940 114158 31952
rect 114152 31912 114416 31940
rect 114152 31900 114158 31912
rect 108945 31875 109003 31881
rect 108816 31844 108896 31872
rect 108816 31832 108822 31844
rect 108868 31816 108896 31844
rect 108945 31841 108957 31875
rect 108991 31841 109003 31875
rect 108945 31835 109003 31841
rect 109865 31875 109923 31881
rect 109865 31841 109877 31875
rect 109911 31872 109923 31875
rect 109954 31872 109960 31884
rect 109911 31844 109960 31872
rect 109911 31841 109923 31844
rect 109865 31835 109923 31841
rect 109954 31832 109960 31844
rect 110012 31832 110018 31884
rect 110874 31832 110880 31884
rect 110932 31832 110938 31884
rect 111613 31875 111671 31881
rect 111613 31841 111625 31875
rect 111659 31872 111671 31875
rect 111886 31872 111892 31884
rect 111659 31844 111892 31872
rect 111659 31841 111671 31844
rect 111613 31835 111671 31841
rect 111886 31832 111892 31844
rect 111944 31832 111950 31884
rect 114388 31881 114416 31912
rect 115198 31900 115204 31952
rect 115256 31940 115262 31952
rect 115584 31940 115612 31980
rect 116026 31968 116032 31980
rect 116084 31968 116090 32020
rect 116305 32011 116363 32017
rect 116305 31977 116317 32011
rect 116351 32008 116363 32011
rect 116351 31980 116716 32008
rect 116351 31977 116363 31980
rect 116305 31971 116363 31977
rect 115256 31912 115612 31940
rect 116044 31940 116072 31968
rect 116581 31943 116639 31949
rect 116581 31940 116593 31943
rect 116044 31912 116593 31940
rect 115256 31900 115262 31912
rect 112349 31875 112407 31881
rect 112349 31841 112361 31875
rect 112395 31872 112407 31875
rect 114373 31875 114431 31881
rect 112395 31844 113312 31872
rect 112395 31841 112407 31844
rect 112349 31835 112407 31841
rect 113284 31816 113312 31844
rect 114373 31841 114385 31875
rect 114419 31841 114431 31875
rect 114373 31835 114431 31841
rect 114462 31832 114468 31884
rect 114520 31872 114526 31884
rect 114520 31844 115244 31872
rect 114520 31832 114526 31844
rect 108298 31764 108304 31816
rect 108356 31764 108362 31816
rect 108482 31764 108488 31816
rect 108540 31764 108546 31816
rect 108850 31764 108856 31816
rect 108908 31764 108914 31816
rect 109773 31807 109831 31813
rect 109773 31773 109785 31807
rect 109819 31804 109831 31807
rect 110414 31804 110420 31816
rect 109819 31776 110420 31804
rect 109819 31773 109831 31776
rect 109773 31767 109831 31773
rect 110414 31764 110420 31776
rect 110472 31804 110478 31816
rect 111340 31807 111398 31813
rect 111340 31804 111352 31807
rect 110472 31776 110920 31804
rect 110472 31764 110478 31776
rect 110892 31736 110920 31776
rect 111076 31776 111352 31804
rect 111076 31736 111104 31776
rect 111340 31773 111352 31776
rect 111386 31773 111398 31807
rect 111340 31767 111398 31773
rect 111794 31764 111800 31816
rect 111852 31804 111858 31816
rect 112165 31807 112223 31813
rect 111852 31776 112116 31804
rect 111852 31764 111858 31776
rect 110892 31708 111104 31736
rect 111337 31671 111395 31677
rect 111337 31637 111349 31671
rect 111383 31668 111395 31671
rect 111426 31668 111432 31680
rect 111383 31640 111432 31668
rect 111383 31637 111395 31640
rect 111337 31631 111395 31637
rect 111426 31628 111432 31640
rect 111484 31628 111490 31680
rect 111518 31628 111524 31680
rect 111576 31668 111582 31680
rect 111797 31671 111855 31677
rect 111797 31668 111809 31671
rect 111576 31640 111809 31668
rect 111576 31628 111582 31640
rect 111797 31637 111809 31640
rect 111843 31637 111855 31671
rect 112088 31668 112116 31776
rect 112165 31773 112177 31807
rect 112211 31773 112223 31807
rect 112165 31767 112223 31773
rect 112533 31807 112591 31813
rect 112533 31773 112545 31807
rect 112579 31804 112591 31807
rect 112993 31807 113051 31813
rect 112993 31804 113005 31807
rect 112579 31776 113005 31804
rect 112579 31773 112591 31776
rect 112533 31767 112591 31773
rect 112993 31773 113005 31776
rect 113039 31804 113051 31807
rect 113039 31776 113128 31804
rect 113039 31773 113051 31776
rect 112993 31767 113051 31773
rect 112180 31736 112208 31767
rect 112346 31736 112352 31748
rect 112180 31708 112352 31736
rect 112346 31696 112352 31708
rect 112404 31696 112410 31748
rect 113100 31736 113128 31776
rect 113266 31764 113272 31816
rect 113324 31764 113330 31816
rect 113821 31807 113879 31813
rect 113821 31773 113833 31807
rect 113867 31804 113879 31807
rect 114002 31804 114008 31816
rect 113867 31776 114008 31804
rect 113867 31773 113879 31776
rect 113821 31767 113879 31773
rect 114002 31764 114008 31776
rect 114060 31764 114066 31816
rect 114094 31764 114100 31816
rect 114152 31764 114158 31816
rect 114833 31807 114891 31813
rect 114833 31773 114845 31807
rect 114879 31804 114891 31807
rect 114922 31804 114928 31816
rect 114879 31776 114928 31804
rect 114879 31773 114891 31776
rect 114833 31767 114891 31773
rect 114922 31764 114928 31776
rect 114980 31764 114986 31816
rect 115216 31813 115244 31844
rect 115109 31807 115167 31813
rect 115109 31773 115121 31807
rect 115155 31773 115167 31807
rect 115109 31767 115167 31773
rect 115201 31807 115259 31813
rect 115201 31773 115213 31807
rect 115247 31804 115259 31807
rect 115477 31807 115535 31813
rect 115477 31804 115489 31807
rect 115247 31776 115489 31804
rect 115247 31773 115259 31776
rect 115201 31767 115259 31773
rect 115477 31773 115489 31776
rect 115523 31773 115535 31807
rect 115584 31804 115612 31912
rect 116581 31909 116593 31912
rect 116627 31909 116639 31943
rect 116688 31940 116716 31980
rect 117130 31968 117136 32020
rect 117188 32008 117194 32020
rect 117317 32011 117375 32017
rect 117317 32008 117329 32011
rect 117188 31980 117329 32008
rect 117188 31968 117194 31980
rect 117317 31977 117329 31980
rect 117363 31977 117375 32011
rect 117317 31971 117375 31977
rect 117424 31980 118096 32008
rect 116854 31940 116860 31952
rect 116688 31912 116860 31940
rect 116581 31903 116639 31909
rect 116854 31900 116860 31912
rect 116912 31940 116918 31952
rect 117424 31940 117452 31980
rect 116912 31912 117452 31940
rect 116912 31900 116918 31912
rect 117590 31900 117596 31952
rect 117648 31940 117654 31952
rect 117869 31943 117927 31949
rect 117869 31940 117881 31943
rect 117648 31912 117881 31940
rect 117648 31900 117654 31912
rect 117869 31909 117881 31912
rect 117915 31909 117927 31943
rect 117869 31903 117927 31909
rect 115934 31832 115940 31884
rect 115992 31832 115998 31884
rect 116394 31832 116400 31884
rect 116452 31872 116458 31884
rect 116452 31844 116900 31872
rect 116452 31832 116458 31844
rect 115661 31807 115719 31813
rect 115661 31804 115673 31807
rect 115584 31776 115673 31804
rect 115477 31767 115535 31773
rect 115661 31773 115673 31776
rect 115707 31773 115719 31807
rect 115661 31767 115719 31773
rect 113450 31736 113456 31748
rect 113100 31708 113456 31736
rect 113450 31696 113456 31708
rect 113508 31696 113514 31748
rect 113910 31696 113916 31748
rect 113968 31736 113974 31748
rect 114189 31739 114247 31745
rect 114189 31736 114201 31739
rect 113968 31708 114201 31736
rect 113968 31696 113974 31708
rect 114189 31705 114201 31708
rect 114235 31736 114247 31739
rect 114278 31736 114284 31748
rect 114235 31708 114284 31736
rect 114235 31705 114247 31708
rect 114189 31699 114247 31705
rect 114278 31696 114284 31708
rect 114336 31696 114342 31748
rect 115124 31736 115152 31767
rect 115750 31764 115756 31816
rect 115808 31804 115814 31816
rect 116872 31813 116900 31844
rect 117314 31832 117320 31884
rect 117372 31872 117378 31884
rect 117501 31875 117559 31881
rect 117501 31872 117513 31875
rect 117372 31844 117513 31872
rect 117372 31832 117378 31844
rect 117501 31841 117513 31844
rect 117547 31841 117559 31875
rect 117501 31835 117559 31841
rect 116029 31807 116087 31813
rect 116029 31804 116041 31807
rect 115808 31776 116041 31804
rect 115808 31764 115814 31776
rect 116029 31773 116041 31776
rect 116075 31773 116087 31807
rect 116765 31807 116823 31813
rect 116765 31804 116777 31807
rect 116029 31767 116087 31773
rect 116228 31776 116777 31804
rect 116228 31748 116256 31776
rect 116765 31773 116777 31776
rect 116811 31773 116823 31807
rect 116765 31767 116823 31773
rect 116857 31807 116915 31813
rect 116857 31773 116869 31807
rect 116903 31804 116915 31807
rect 116946 31804 116952 31816
rect 116903 31776 116952 31804
rect 116903 31773 116915 31776
rect 116857 31767 116915 31773
rect 116946 31764 116952 31776
rect 117004 31764 117010 31816
rect 117041 31807 117099 31813
rect 117041 31773 117053 31807
rect 117087 31804 117099 31807
rect 117087 31776 117268 31804
rect 117087 31773 117099 31776
rect 117041 31767 117099 31773
rect 116210 31736 116216 31748
rect 115124 31708 116216 31736
rect 116210 31696 116216 31708
rect 116268 31696 116274 31748
rect 117240 31736 117268 31776
rect 117590 31764 117596 31816
rect 117648 31764 117654 31816
rect 118068 31813 118096 31980
rect 118053 31807 118111 31813
rect 118053 31773 118065 31807
rect 118099 31773 118111 31807
rect 118053 31767 118111 31773
rect 118237 31807 118295 31813
rect 118237 31773 118249 31807
rect 118283 31804 118295 31807
rect 118510 31804 118516 31816
rect 118283 31776 118516 31804
rect 118283 31773 118295 31776
rect 118237 31767 118295 31773
rect 118510 31764 118516 31776
rect 118568 31764 118574 31816
rect 117958 31736 117964 31748
rect 117240 31708 117964 31736
rect 117958 31696 117964 31708
rect 118016 31696 118022 31748
rect 114370 31668 114376 31680
rect 112088 31640 114376 31668
rect 111797 31631 111855 31637
rect 114370 31628 114376 31640
rect 114428 31668 114434 31680
rect 115842 31668 115848 31680
rect 114428 31640 115848 31668
rect 114428 31628 114434 31640
rect 115842 31628 115848 31640
rect 115900 31628 115906 31680
rect 115934 31628 115940 31680
rect 115992 31668 115998 31680
rect 116670 31668 116676 31680
rect 115992 31640 116676 31668
rect 115992 31628 115998 31640
rect 116670 31628 116676 31640
rect 116728 31668 116734 31680
rect 117222 31668 117228 31680
rect 116728 31640 117228 31668
rect 116728 31628 116734 31640
rect 117222 31628 117228 31640
rect 117280 31628 117286 31680
rect 118326 31628 118332 31680
rect 118384 31628 118390 31680
rect 1104 31578 7912 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 7912 31578
rect 1104 31504 7912 31526
rect 108008 31578 118864 31600
rect 108008 31526 113650 31578
rect 113702 31526 113714 31578
rect 113766 31526 113778 31578
rect 113830 31526 113842 31578
rect 113894 31526 113906 31578
rect 113958 31526 118864 31578
rect 108008 31504 118864 31526
rect 110966 31424 110972 31476
rect 111024 31464 111030 31476
rect 111153 31467 111211 31473
rect 111153 31464 111165 31467
rect 111024 31436 111165 31464
rect 111024 31424 111030 31436
rect 111153 31433 111165 31436
rect 111199 31433 111211 31467
rect 111886 31464 111892 31476
rect 111153 31427 111211 31433
rect 111444 31436 111892 31464
rect 108850 31356 108856 31408
rect 108908 31356 108914 31408
rect 110046 31356 110052 31408
rect 110104 31396 110110 31408
rect 111305 31399 111363 31405
rect 111305 31396 111317 31399
rect 110104 31368 111317 31396
rect 110104 31356 110110 31368
rect 111305 31365 111317 31368
rect 111351 31396 111363 31399
rect 111444 31396 111472 31436
rect 111886 31424 111892 31436
rect 111944 31424 111950 31476
rect 111981 31467 112039 31473
rect 111981 31433 111993 31467
rect 112027 31464 112039 31467
rect 112162 31464 112168 31476
rect 112027 31436 112168 31464
rect 112027 31433 112039 31436
rect 111981 31427 112039 31433
rect 112162 31424 112168 31436
rect 112220 31424 112226 31476
rect 112438 31424 112444 31476
rect 112496 31424 112502 31476
rect 114462 31424 114468 31476
rect 114520 31424 114526 31476
rect 115477 31467 115535 31473
rect 115477 31464 115489 31467
rect 114572 31436 115489 31464
rect 111351 31368 111472 31396
rect 111521 31399 111579 31405
rect 111351 31365 111363 31368
rect 111305 31359 111363 31365
rect 111521 31365 111533 31399
rect 111567 31396 111579 31399
rect 111794 31396 111800 31408
rect 111567 31368 111800 31396
rect 111567 31365 111579 31368
rect 111521 31359 111579 31365
rect 111794 31356 111800 31368
rect 111852 31356 111858 31408
rect 113266 31356 113272 31408
rect 113324 31396 113330 31408
rect 113324 31368 113680 31396
rect 113324 31356 113330 31368
rect 109586 31288 109592 31340
rect 109644 31328 109650 31340
rect 110601 31331 110659 31337
rect 110601 31328 110613 31331
rect 109644 31300 110613 31328
rect 109644 31288 109650 31300
rect 110601 31297 110613 31300
rect 110647 31297 110659 31331
rect 110601 31291 110659 31297
rect 111260 31300 111840 31328
rect 110417 31263 110475 31269
rect 110417 31229 110429 31263
rect 110463 31229 110475 31263
rect 110417 31223 110475 31229
rect 108298 31152 108304 31204
rect 108356 31192 108362 31204
rect 109037 31195 109095 31201
rect 109037 31192 109049 31195
rect 108356 31164 109049 31192
rect 108356 31152 108362 31164
rect 109037 31161 109049 31164
rect 109083 31161 109095 31195
rect 110432 31192 110460 31223
rect 110506 31220 110512 31272
rect 110564 31220 110570 31272
rect 110598 31192 110604 31204
rect 110432 31164 110604 31192
rect 109037 31155 109095 31161
rect 110598 31152 110604 31164
rect 110656 31152 110662 31204
rect 110969 31195 111027 31201
rect 110969 31161 110981 31195
rect 111015 31192 111027 31195
rect 111260 31192 111288 31300
rect 111015 31164 111288 31192
rect 111812 31192 111840 31300
rect 111886 31288 111892 31340
rect 111944 31288 111950 31340
rect 111978 31288 111984 31340
rect 112036 31328 112042 31340
rect 112073 31331 112131 31337
rect 112073 31328 112085 31331
rect 112036 31300 112085 31328
rect 112036 31288 112042 31300
rect 112073 31297 112085 31300
rect 112119 31297 112131 31331
rect 112073 31291 112131 31297
rect 112254 31288 112260 31340
rect 112312 31288 112318 31340
rect 112441 31331 112499 31337
rect 112441 31297 112453 31331
rect 112487 31297 112499 31331
rect 112441 31291 112499 31297
rect 112717 31331 112775 31337
rect 112717 31297 112729 31331
rect 112763 31297 112775 31331
rect 112717 31291 112775 31297
rect 111904 31260 111932 31288
rect 112346 31260 112352 31272
rect 111904 31232 112352 31260
rect 112346 31220 112352 31232
rect 112404 31260 112410 31272
rect 112456 31260 112484 31291
rect 112404 31232 112484 31260
rect 112404 31220 112410 31232
rect 112530 31220 112536 31272
rect 112588 31220 112594 31272
rect 112732 31192 112760 31291
rect 112806 31288 112812 31340
rect 112864 31328 112870 31340
rect 113085 31331 113143 31337
rect 113085 31328 113097 31331
rect 112864 31300 113097 31328
rect 112864 31288 112870 31300
rect 113085 31297 113097 31300
rect 113131 31297 113143 31331
rect 113085 31291 113143 31297
rect 113450 31288 113456 31340
rect 113508 31288 113514 31340
rect 113652 31337 113680 31368
rect 113637 31331 113695 31337
rect 113637 31297 113649 31331
rect 113683 31297 113695 31331
rect 113637 31291 113695 31297
rect 113818 31288 113824 31340
rect 113876 31288 113882 31340
rect 114094 31288 114100 31340
rect 114152 31288 114158 31340
rect 114278 31288 114284 31340
rect 114336 31328 114342 31340
rect 114373 31331 114431 31337
rect 114373 31328 114385 31331
rect 114336 31300 114385 31328
rect 114336 31288 114342 31300
rect 114373 31297 114385 31300
rect 114419 31328 114431 31331
rect 114572 31328 114600 31436
rect 115477 31433 115489 31436
rect 115523 31464 115535 31467
rect 116118 31464 116124 31476
rect 115523 31436 116124 31464
rect 115523 31433 115535 31436
rect 115477 31427 115535 31433
rect 116118 31424 116124 31436
rect 116176 31424 116182 31476
rect 116578 31424 116584 31476
rect 116636 31424 116642 31476
rect 117774 31464 117780 31476
rect 116688 31436 117780 31464
rect 115106 31356 115112 31408
rect 115164 31396 115170 31408
rect 116688 31396 116716 31436
rect 117774 31424 117780 31436
rect 117832 31424 117838 31476
rect 117958 31424 117964 31476
rect 118016 31464 118022 31476
rect 118053 31467 118111 31473
rect 118053 31464 118065 31467
rect 118016 31436 118065 31464
rect 118016 31424 118022 31436
rect 118053 31433 118065 31436
rect 118099 31433 118111 31467
rect 118053 31427 118111 31433
rect 115164 31368 116716 31396
rect 115164 31356 115170 31368
rect 116762 31356 116768 31408
rect 116820 31396 116826 31408
rect 116946 31396 116952 31408
rect 116820 31368 116952 31396
rect 116820 31356 116826 31368
rect 116946 31356 116952 31368
rect 117004 31356 117010 31408
rect 117317 31399 117375 31405
rect 117317 31365 117329 31399
rect 117363 31396 117375 31399
rect 117593 31399 117651 31405
rect 117593 31396 117605 31399
rect 117363 31368 117605 31396
rect 117363 31365 117375 31368
rect 117317 31359 117375 31365
rect 117593 31365 117605 31368
rect 117639 31365 117651 31399
rect 117593 31359 117651 31365
rect 114419 31300 114600 31328
rect 114419 31297 114431 31300
rect 114373 31291 114431 31297
rect 114646 31288 114652 31340
rect 114704 31328 114710 31340
rect 114925 31331 114983 31337
rect 114925 31328 114937 31331
rect 114704 31300 114937 31328
rect 114704 31288 114710 31300
rect 114925 31297 114937 31300
rect 114971 31297 114983 31331
rect 114925 31291 114983 31297
rect 115385 31331 115443 31337
rect 115385 31297 115397 31331
rect 115431 31328 115443 31331
rect 115934 31328 115940 31340
rect 115431 31300 115940 31328
rect 115431 31297 115443 31300
rect 115385 31291 115443 31297
rect 115934 31288 115940 31300
rect 115992 31328 115998 31340
rect 116213 31331 116271 31337
rect 116213 31328 116225 31331
rect 115992 31300 116225 31328
rect 115992 31288 115998 31300
rect 116213 31297 116225 31300
rect 116259 31297 116271 31331
rect 116213 31291 116271 31297
rect 116394 31288 116400 31340
rect 116452 31288 116458 31340
rect 116486 31288 116492 31340
rect 116544 31288 116550 31340
rect 116670 31288 116676 31340
rect 116728 31288 116734 31340
rect 112993 31263 113051 31269
rect 112993 31229 113005 31263
rect 113039 31260 113051 31263
rect 114112 31260 114140 31288
rect 115017 31263 115075 31269
rect 115017 31260 115029 31263
rect 113039 31232 114140 31260
rect 114204 31232 115029 31260
rect 113039 31229 113051 31232
rect 112993 31223 113051 31229
rect 113358 31192 113364 31204
rect 111812 31164 113364 31192
rect 111015 31161 111027 31164
rect 110969 31155 111027 31161
rect 113358 31152 113364 31164
rect 113416 31192 113422 31204
rect 114204 31192 114232 31232
rect 115017 31229 115029 31232
rect 115063 31229 115075 31263
rect 115017 31223 115075 31229
rect 115109 31263 115167 31269
rect 115109 31229 115121 31263
rect 115155 31229 115167 31263
rect 115109 31223 115167 31229
rect 113416 31164 114232 31192
rect 113416 31152 113422 31164
rect 114370 31152 114376 31204
rect 114428 31192 114434 31204
rect 115124 31192 115152 31223
rect 116578 31220 116584 31272
rect 116636 31260 116642 31272
rect 117332 31260 117360 31359
rect 117406 31288 117412 31340
rect 117464 31288 117470 31340
rect 118237 31331 118295 31337
rect 118237 31297 118249 31331
rect 118283 31328 118295 31331
rect 118510 31328 118516 31340
rect 118283 31300 118516 31328
rect 118283 31297 118295 31300
rect 118237 31291 118295 31297
rect 118510 31288 118516 31300
rect 118568 31288 118574 31340
rect 116636 31232 117360 31260
rect 116636 31220 116642 31232
rect 117958 31192 117964 31204
rect 114428 31164 115152 31192
rect 115400 31164 117964 31192
rect 114428 31152 114434 31164
rect 108758 31084 108764 31136
rect 108816 31124 108822 31136
rect 109221 31127 109279 31133
rect 109221 31124 109233 31127
rect 108816 31096 109233 31124
rect 108816 31084 108822 31096
rect 109221 31093 109233 31096
rect 109267 31093 109279 31127
rect 109221 31087 109279 31093
rect 111334 31084 111340 31136
rect 111392 31084 111398 31136
rect 111610 31084 111616 31136
rect 111668 31124 111674 31136
rect 114186 31124 114192 31136
rect 111668 31096 114192 31124
rect 111668 31084 111674 31096
rect 114186 31084 114192 31096
rect 114244 31084 114250 31136
rect 114554 31084 114560 31136
rect 114612 31084 114618 31136
rect 114830 31084 114836 31136
rect 114888 31124 114894 31136
rect 115400 31124 115428 31164
rect 117958 31152 117964 31164
rect 118016 31152 118022 31204
rect 114888 31096 115428 31124
rect 114888 31084 114894 31096
rect 116302 31084 116308 31136
rect 116360 31084 116366 31136
rect 117130 31084 117136 31136
rect 117188 31124 117194 31136
rect 117777 31127 117835 31133
rect 117777 31124 117789 31127
rect 117188 31096 117789 31124
rect 117188 31084 117194 31096
rect 117777 31093 117789 31096
rect 117823 31093 117835 31127
rect 117777 31087 117835 31093
rect 1104 31034 7912 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 7912 31034
rect 1104 30960 7912 30982
rect 108008 31034 118864 31056
rect 108008 30982 112914 31034
rect 112966 30982 112978 31034
rect 113030 30982 113042 31034
rect 113094 30982 113106 31034
rect 113158 30982 113170 31034
rect 113222 30982 118864 31034
rect 108008 30960 118864 30982
rect 109497 30923 109555 30929
rect 109497 30889 109509 30923
rect 109543 30920 109555 30923
rect 109586 30920 109592 30932
rect 109543 30892 109592 30920
rect 109543 30889 109555 30892
rect 109497 30883 109555 30889
rect 109586 30880 109592 30892
rect 109644 30880 109650 30932
rect 109773 30923 109831 30929
rect 109773 30889 109785 30923
rect 109819 30920 109831 30923
rect 110506 30920 110512 30932
rect 109819 30892 110512 30920
rect 109819 30889 109831 30892
rect 109773 30883 109831 30889
rect 110506 30880 110512 30892
rect 110564 30880 110570 30932
rect 111426 30880 111432 30932
rect 111484 30880 111490 30932
rect 111702 30880 111708 30932
rect 111760 30920 111766 30932
rect 112533 30923 112591 30929
rect 112533 30920 112545 30923
rect 111760 30892 112545 30920
rect 111760 30880 111766 30892
rect 112533 30889 112545 30892
rect 112579 30889 112591 30923
rect 112533 30883 112591 30889
rect 114281 30923 114339 30929
rect 114281 30889 114293 30923
rect 114327 30920 114339 30923
rect 114646 30920 114652 30932
rect 114327 30892 114652 30920
rect 114327 30889 114339 30892
rect 114281 30883 114339 30889
rect 114646 30880 114652 30892
rect 114704 30880 114710 30932
rect 116026 30880 116032 30932
rect 116084 30880 116090 30932
rect 116578 30920 116584 30932
rect 116320 30892 116584 30920
rect 110046 30812 110052 30864
rect 110104 30812 110110 30864
rect 112257 30855 112315 30861
rect 112257 30821 112269 30855
rect 112303 30821 112315 30855
rect 112257 30815 112315 30821
rect 109313 30787 109371 30793
rect 109313 30753 109325 30787
rect 109359 30784 109371 30787
rect 110874 30784 110880 30796
rect 109359 30756 110880 30784
rect 109359 30753 109371 30756
rect 109313 30747 109371 30753
rect 110874 30744 110880 30756
rect 110932 30744 110938 30796
rect 111521 30787 111579 30793
rect 111521 30753 111533 30787
rect 111567 30784 111579 30787
rect 111886 30784 111892 30796
rect 111567 30756 111892 30784
rect 111567 30753 111579 30756
rect 111521 30747 111579 30753
rect 111886 30744 111892 30756
rect 111944 30784 111950 30796
rect 111944 30756 112116 30784
rect 111944 30744 111950 30756
rect 109218 30676 109224 30728
rect 109276 30676 109282 30728
rect 109678 30676 109684 30728
rect 109736 30676 109742 30728
rect 110233 30719 110291 30725
rect 110233 30685 110245 30719
rect 110279 30716 110291 30719
rect 110322 30716 110328 30728
rect 110279 30688 110328 30716
rect 110279 30685 110291 30688
rect 110233 30679 110291 30685
rect 110322 30676 110328 30688
rect 110380 30676 110386 30728
rect 110417 30719 110475 30725
rect 110417 30685 110429 30719
rect 110463 30716 110475 30719
rect 110506 30716 110512 30728
rect 110463 30688 110512 30716
rect 110463 30685 110475 30688
rect 110417 30679 110475 30685
rect 110506 30676 110512 30688
rect 110564 30676 110570 30728
rect 111334 30676 111340 30728
rect 111392 30716 111398 30728
rect 111610 30716 111616 30728
rect 111392 30688 111616 30716
rect 111392 30676 111398 30688
rect 111610 30676 111616 30688
rect 111668 30676 111674 30728
rect 111981 30719 112039 30725
rect 111981 30716 111993 30719
rect 111904 30688 111993 30716
rect 111904 30660 111932 30688
rect 111981 30685 111993 30688
rect 112027 30685 112039 30719
rect 111981 30679 112039 30685
rect 111886 30608 111892 30660
rect 111944 30608 111950 30660
rect 112088 30648 112116 30756
rect 112272 30716 112300 30815
rect 115106 30812 115112 30864
rect 115164 30852 115170 30864
rect 116320 30852 116348 30892
rect 116578 30880 116584 30892
rect 116636 30880 116642 30932
rect 117130 30880 117136 30932
rect 117188 30880 117194 30932
rect 117314 30880 117320 30932
rect 117372 30880 117378 30932
rect 115164 30824 116348 30852
rect 115164 30812 115170 30824
rect 113266 30744 113272 30796
rect 113324 30784 113330 30796
rect 114005 30787 114063 30793
rect 113324 30756 113956 30784
rect 113324 30744 113330 30756
rect 112441 30719 112499 30725
rect 112441 30716 112453 30719
rect 112272 30688 112453 30716
rect 112441 30685 112453 30688
rect 112487 30685 112499 30719
rect 112441 30679 112499 30685
rect 112901 30719 112959 30725
rect 112901 30685 112913 30719
rect 112947 30685 112959 30719
rect 112901 30679 112959 30685
rect 112257 30651 112315 30657
rect 112257 30648 112269 30651
rect 112088 30620 112269 30648
rect 112257 30617 112269 30620
rect 112303 30617 112315 30651
rect 112916 30648 112944 30679
rect 113082 30676 113088 30728
rect 113140 30676 113146 30728
rect 113177 30719 113235 30725
rect 113177 30685 113189 30719
rect 113223 30716 113235 30719
rect 113818 30716 113824 30728
rect 113223 30688 113824 30716
rect 113223 30685 113235 30688
rect 113177 30679 113235 30685
rect 113818 30676 113824 30688
rect 113876 30676 113882 30728
rect 113928 30725 113956 30756
rect 114005 30753 114017 30787
rect 114051 30784 114063 30787
rect 114278 30784 114284 30796
rect 114051 30756 114284 30784
rect 114051 30753 114063 30756
rect 114005 30747 114063 30753
rect 114278 30744 114284 30756
rect 114336 30744 114342 30796
rect 114462 30744 114468 30796
rect 114520 30784 114526 30796
rect 114741 30787 114799 30793
rect 114741 30784 114753 30787
rect 114520 30756 114753 30784
rect 114520 30744 114526 30756
rect 114741 30753 114753 30756
rect 114787 30753 114799 30787
rect 114741 30747 114799 30753
rect 114922 30744 114928 30796
rect 114980 30784 114986 30796
rect 115474 30784 115480 30796
rect 114980 30756 115480 30784
rect 114980 30744 114986 30756
rect 115474 30744 115480 30756
rect 115532 30784 115538 30796
rect 116121 30787 116179 30793
rect 116121 30784 116133 30787
rect 115532 30756 116133 30784
rect 115532 30744 115538 30756
rect 116121 30753 116133 30756
rect 116167 30753 116179 30787
rect 116121 30747 116179 30753
rect 113913 30719 113971 30725
rect 113913 30685 113925 30719
rect 113959 30716 113971 30719
rect 114373 30719 114431 30725
rect 114373 30716 114385 30719
rect 113959 30688 114385 30716
rect 113959 30685 113971 30688
rect 113913 30679 113971 30685
rect 114373 30685 114385 30688
rect 114419 30685 114431 30719
rect 114373 30679 114431 30685
rect 114557 30719 114615 30725
rect 114557 30685 114569 30719
rect 114603 30716 114615 30719
rect 114646 30716 114652 30728
rect 114603 30688 114652 30716
rect 114603 30685 114615 30688
rect 114557 30679 114615 30685
rect 114646 30676 114652 30688
rect 114704 30676 114710 30728
rect 114833 30719 114891 30725
rect 114833 30685 114845 30719
rect 114879 30685 114891 30719
rect 114833 30679 114891 30685
rect 115845 30719 115903 30725
rect 115845 30685 115857 30719
rect 115891 30716 115903 30719
rect 116026 30716 116032 30728
rect 115891 30688 116032 30716
rect 115891 30685 115903 30688
rect 115845 30679 115903 30685
rect 113269 30651 113327 30657
rect 113269 30648 113281 30651
rect 112916 30620 113281 30648
rect 112257 30611 112315 30617
rect 113269 30617 113281 30620
rect 113315 30648 113327 30651
rect 113358 30648 113364 30660
rect 113315 30620 113364 30648
rect 113315 30617 113327 30620
rect 113269 30611 113327 30617
rect 113358 30608 113364 30620
rect 113416 30608 113422 30660
rect 113453 30651 113511 30657
rect 113453 30617 113465 30651
rect 113499 30617 113511 30651
rect 113453 30611 113511 30617
rect 111797 30583 111855 30589
rect 111797 30549 111809 30583
rect 111843 30580 111855 30583
rect 112070 30580 112076 30592
rect 111843 30552 112076 30580
rect 111843 30549 111855 30552
rect 111797 30543 111855 30549
rect 112070 30540 112076 30552
rect 112128 30540 112134 30592
rect 113082 30540 113088 30592
rect 113140 30580 113146 30592
rect 113468 30580 113496 30611
rect 113542 30608 113548 30660
rect 113600 30648 113606 30660
rect 114465 30651 114523 30657
rect 114465 30648 114477 30651
rect 113600 30620 114477 30648
rect 113600 30608 113606 30620
rect 114465 30617 114477 30620
rect 114511 30617 114523 30651
rect 114465 30611 114523 30617
rect 113140 30552 113496 30580
rect 113637 30583 113695 30589
rect 113140 30540 113146 30552
rect 113637 30549 113649 30583
rect 113683 30580 113695 30583
rect 114002 30580 114008 30592
rect 113683 30552 114008 30580
rect 113683 30549 113695 30552
rect 113637 30543 113695 30549
rect 114002 30540 114008 30552
rect 114060 30580 114066 30592
rect 114848 30580 114876 30679
rect 116026 30676 116032 30688
rect 116084 30676 116090 30728
rect 116320 30725 116348 30824
rect 116394 30812 116400 30864
rect 116452 30852 116458 30864
rect 116854 30852 116860 30864
rect 116452 30824 116860 30852
rect 116452 30812 116458 30824
rect 116854 30812 116860 30824
rect 116912 30852 116918 30864
rect 117225 30855 117283 30861
rect 117225 30852 117237 30855
rect 116912 30824 117237 30852
rect 116912 30812 116918 30824
rect 117225 30821 117237 30824
rect 117271 30821 117283 30855
rect 117225 30815 117283 30821
rect 118053 30787 118111 30793
rect 118053 30784 118065 30787
rect 116964 30756 118065 30784
rect 116964 30728 116992 30756
rect 118053 30753 118065 30756
rect 118099 30753 118111 30787
rect 118053 30747 118111 30753
rect 116305 30719 116363 30725
rect 116305 30685 116317 30719
rect 116351 30685 116363 30719
rect 116305 30679 116363 30685
rect 116394 30676 116400 30728
rect 116452 30716 116458 30728
rect 116581 30719 116639 30725
rect 116581 30716 116593 30719
rect 116452 30688 116593 30716
rect 116452 30676 116458 30688
rect 116581 30685 116593 30688
rect 116627 30685 116639 30719
rect 116581 30679 116639 30685
rect 116765 30719 116823 30725
rect 116765 30685 116777 30719
rect 116811 30716 116823 30719
rect 116857 30719 116915 30725
rect 116857 30716 116869 30719
rect 116811 30688 116869 30716
rect 116811 30685 116823 30688
rect 116765 30679 116823 30685
rect 116857 30685 116869 30688
rect 116903 30716 116915 30719
rect 116946 30716 116952 30728
rect 116903 30688 116952 30716
rect 116903 30685 116915 30688
rect 116857 30679 116915 30685
rect 116946 30676 116952 30688
rect 117004 30676 117010 30728
rect 117958 30676 117964 30728
rect 118016 30676 118022 30728
rect 118237 30719 118295 30725
rect 118237 30685 118249 30719
rect 118283 30716 118295 30719
rect 118326 30716 118332 30728
rect 118283 30688 118332 30716
rect 118283 30685 118295 30688
rect 118237 30679 118295 30685
rect 118326 30676 118332 30688
rect 118384 30676 118390 30728
rect 115934 30608 115940 30660
rect 115992 30648 115998 30660
rect 116673 30651 116731 30657
rect 116673 30648 116685 30651
rect 115992 30620 116685 30648
rect 115992 30608 115998 30620
rect 116673 30617 116685 30620
rect 116719 30617 116731 30651
rect 116673 30611 116731 30617
rect 116780 30620 117820 30648
rect 114060 30552 114876 30580
rect 114060 30540 114066 30552
rect 116486 30540 116492 30592
rect 116544 30540 116550 30592
rect 116578 30540 116584 30592
rect 116636 30580 116642 30592
rect 116780 30580 116808 30620
rect 116636 30552 116808 30580
rect 116949 30583 117007 30589
rect 116636 30540 116642 30552
rect 116949 30549 116961 30583
rect 116995 30580 117007 30583
rect 117130 30580 117136 30592
rect 116995 30552 117136 30580
rect 116995 30549 117007 30552
rect 116949 30543 117007 30549
rect 117130 30540 117136 30552
rect 117188 30540 117194 30592
rect 117590 30540 117596 30592
rect 117648 30540 117654 30592
rect 117792 30589 117820 30620
rect 117777 30583 117835 30589
rect 117777 30549 117789 30583
rect 117823 30549 117835 30583
rect 117777 30543 117835 30549
rect 1104 30490 7912 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 7912 30490
rect 1104 30416 7912 30438
rect 108008 30490 118864 30512
rect 108008 30438 113650 30490
rect 113702 30438 113714 30490
rect 113766 30438 113778 30490
rect 113830 30438 113842 30490
rect 113894 30438 113906 30490
rect 113958 30438 118864 30490
rect 108008 30416 118864 30438
rect 109218 30336 109224 30388
rect 109276 30336 109282 30388
rect 110874 30336 110880 30388
rect 110932 30376 110938 30388
rect 111518 30376 111524 30388
rect 110932 30348 111524 30376
rect 110932 30336 110938 30348
rect 109586 30268 109592 30320
rect 109644 30308 109650 30320
rect 110414 30308 110420 30320
rect 109644 30280 110420 30308
rect 109644 30268 109650 30280
rect 109770 30200 109776 30252
rect 109828 30200 109834 30252
rect 109862 30200 109868 30252
rect 109920 30240 109926 30252
rect 110064 30249 110092 30280
rect 110414 30268 110420 30280
rect 110472 30268 110478 30320
rect 111153 30311 111211 30317
rect 111153 30308 111165 30311
rect 110524 30280 111165 30308
rect 109957 30243 110015 30249
rect 109957 30240 109969 30243
rect 109920 30212 109969 30240
rect 109920 30200 109926 30212
rect 109957 30209 109969 30212
rect 110003 30209 110015 30243
rect 109957 30203 110015 30209
rect 110049 30243 110107 30249
rect 110049 30209 110061 30243
rect 110095 30209 110107 30243
rect 110049 30203 110107 30209
rect 110138 30200 110144 30252
rect 110196 30200 110202 30252
rect 110524 30249 110552 30280
rect 111153 30277 111165 30280
rect 111199 30277 111211 30311
rect 111153 30271 111211 30277
rect 110509 30243 110567 30249
rect 110509 30240 110521 30243
rect 110432 30212 110521 30240
rect 110432 30181 110460 30212
rect 110509 30209 110521 30212
rect 110555 30209 110567 30243
rect 110509 30203 110567 30209
rect 110598 30200 110604 30252
rect 110656 30200 110662 30252
rect 110785 30243 110843 30249
rect 110785 30209 110797 30243
rect 110831 30209 110843 30243
rect 110785 30203 110843 30209
rect 109681 30175 109739 30181
rect 109681 30141 109693 30175
rect 109727 30172 109739 30175
rect 110417 30175 110475 30181
rect 110417 30172 110429 30175
rect 109727 30144 110429 30172
rect 109727 30141 109739 30144
rect 109681 30135 109739 30141
rect 110417 30141 110429 30144
rect 110463 30141 110475 30175
rect 110417 30135 110475 30141
rect 110800 30172 110828 30203
rect 110874 30200 110880 30252
rect 110932 30200 110938 30252
rect 111242 30240 111248 30252
rect 110984 30212 111248 30240
rect 110984 30172 111012 30212
rect 111242 30200 111248 30212
rect 111300 30240 111306 30252
rect 111444 30249 111472 30348
rect 111518 30336 111524 30348
rect 111576 30336 111582 30388
rect 112070 30336 112076 30388
rect 112128 30336 112134 30388
rect 113542 30336 113548 30388
rect 113600 30376 113606 30388
rect 113637 30379 113695 30385
rect 113637 30376 113649 30379
rect 113600 30348 113649 30376
rect 113600 30336 113606 30348
rect 113637 30345 113649 30348
rect 113683 30345 113695 30379
rect 113637 30339 113695 30345
rect 114922 30336 114928 30388
rect 114980 30376 114986 30388
rect 117130 30376 117136 30388
rect 114980 30348 117136 30376
rect 114980 30336 114986 30348
rect 111889 30311 111947 30317
rect 111889 30277 111901 30311
rect 111935 30308 111947 30311
rect 112088 30308 112116 30336
rect 112530 30308 112536 30320
rect 111935 30280 112116 30308
rect 112180 30280 112536 30308
rect 111935 30277 111947 30280
rect 111889 30271 111947 30277
rect 111337 30243 111395 30249
rect 111337 30240 111349 30243
rect 111300 30212 111349 30240
rect 111300 30200 111306 30212
rect 111337 30209 111349 30212
rect 111383 30209 111395 30243
rect 111337 30203 111395 30209
rect 111429 30243 111487 30249
rect 111429 30209 111441 30243
rect 111475 30209 111487 30243
rect 111429 30203 111487 30209
rect 111705 30243 111763 30249
rect 111705 30209 111717 30243
rect 111751 30209 111763 30243
rect 111705 30203 111763 30209
rect 110800 30144 111012 30172
rect 111061 30175 111119 30181
rect 109405 30107 109463 30113
rect 109405 30073 109417 30107
rect 109451 30104 109463 30107
rect 110800 30104 110828 30144
rect 111061 30141 111073 30175
rect 111107 30172 111119 30175
rect 111720 30172 111748 30203
rect 111978 30200 111984 30252
rect 112036 30200 112042 30252
rect 112070 30200 112076 30252
rect 112128 30240 112134 30252
rect 112180 30240 112208 30280
rect 112530 30268 112536 30280
rect 112588 30268 112594 30320
rect 113269 30311 113327 30317
rect 113269 30277 113281 30311
rect 113315 30308 113327 30311
rect 113913 30311 113971 30317
rect 113913 30308 113925 30311
rect 113315 30280 113925 30308
rect 113315 30277 113327 30280
rect 113269 30271 113327 30277
rect 113913 30277 113925 30280
rect 113959 30277 113971 30311
rect 113913 30271 113971 30277
rect 114024 30311 114082 30317
rect 114024 30277 114036 30311
rect 114070 30308 114082 30311
rect 114554 30308 114560 30320
rect 114070 30280 114560 30308
rect 114070 30277 114082 30280
rect 114024 30271 114082 30277
rect 114554 30268 114560 30280
rect 114612 30268 114618 30320
rect 115477 30311 115535 30317
rect 115477 30308 115489 30311
rect 115308 30280 115489 30308
rect 112128 30212 112208 30240
rect 112128 30200 112134 30212
rect 112254 30200 112260 30252
rect 112312 30200 112318 30252
rect 112806 30200 112812 30252
rect 112864 30240 112870 30252
rect 113453 30243 113511 30249
rect 113453 30240 113465 30243
rect 112864 30212 113465 30240
rect 112864 30200 112870 30212
rect 113453 30209 113465 30212
rect 113499 30209 113511 30243
rect 113453 30203 113511 30209
rect 113726 30200 113732 30252
rect 113784 30200 113790 30252
rect 113821 30243 113879 30249
rect 113821 30209 113833 30243
rect 113867 30209 113879 30243
rect 113821 30203 113879 30209
rect 115109 30243 115167 30249
rect 115109 30209 115121 30243
rect 115155 30209 115167 30243
rect 115109 30203 115167 30209
rect 115201 30243 115259 30249
rect 115201 30209 115213 30243
rect 115247 30240 115259 30243
rect 115308 30240 115336 30280
rect 115477 30277 115489 30280
rect 115523 30277 115535 30311
rect 115693 30311 115751 30317
rect 115693 30308 115705 30311
rect 115477 30271 115535 30277
rect 115676 30277 115705 30308
rect 115739 30308 115751 30311
rect 116302 30308 116308 30320
rect 115739 30280 116308 30308
rect 115739 30277 115751 30280
rect 115676 30271 115751 30277
rect 115247 30212 115336 30240
rect 115247 30209 115259 30212
rect 115201 30203 115259 30209
rect 111886 30172 111892 30184
rect 111107 30144 111892 30172
rect 111107 30141 111119 30144
rect 111061 30135 111119 30141
rect 111886 30132 111892 30144
rect 111944 30132 111950 30184
rect 113836 30172 113864 30203
rect 111996 30144 113864 30172
rect 111996 30113 112024 30144
rect 114186 30132 114192 30184
rect 114244 30132 114250 30184
rect 109451 30076 110828 30104
rect 111981 30107 112039 30113
rect 109451 30073 109463 30076
rect 109405 30067 109463 30073
rect 111981 30073 111993 30107
rect 112027 30073 112039 30107
rect 111981 30067 112039 30073
rect 114097 30107 114155 30113
rect 114097 30073 114109 30107
rect 114143 30104 114155 30107
rect 115014 30104 115020 30116
rect 114143 30076 115020 30104
rect 114143 30073 114155 30076
rect 114097 30067 114155 30073
rect 115014 30064 115020 30076
rect 115072 30064 115078 30116
rect 115124 30104 115152 30203
rect 115308 30172 115336 30212
rect 115385 30243 115443 30249
rect 115385 30209 115397 30243
rect 115431 30240 115443 30243
rect 115676 30240 115704 30271
rect 116302 30268 116308 30280
rect 116360 30268 116366 30320
rect 116412 30252 116440 30348
rect 117130 30336 117136 30348
rect 117188 30376 117194 30388
rect 117866 30376 117872 30388
rect 117188 30348 117872 30376
rect 117188 30336 117194 30348
rect 117866 30336 117872 30348
rect 117924 30336 117930 30388
rect 116854 30268 116860 30320
rect 116912 30268 116918 30320
rect 115431 30212 115704 30240
rect 116213 30243 116271 30249
rect 115431 30209 115443 30212
rect 115385 30203 115443 30209
rect 116213 30209 116225 30243
rect 116259 30240 116271 30243
rect 116394 30240 116400 30252
rect 116259 30212 116400 30240
rect 116259 30209 116271 30212
rect 116213 30203 116271 30209
rect 116394 30200 116400 30212
rect 116452 30200 116458 30252
rect 116486 30200 116492 30252
rect 116544 30200 116550 30252
rect 116578 30200 116584 30252
rect 116636 30240 116642 30252
rect 116719 30243 116777 30249
rect 116719 30240 116731 30243
rect 116636 30212 116731 30240
rect 116636 30200 116642 30212
rect 116719 30209 116731 30212
rect 116765 30209 116777 30243
rect 116719 30203 116777 30209
rect 116946 30200 116952 30252
rect 117004 30200 117010 30252
rect 117147 30249 117175 30336
rect 117590 30268 117596 30320
rect 117648 30308 117654 30320
rect 117648 30280 118004 30308
rect 117648 30268 117654 30280
rect 117132 30243 117190 30249
rect 117132 30209 117144 30243
rect 117178 30209 117190 30243
rect 117132 30203 117190 30209
rect 117222 30200 117228 30252
rect 117280 30200 117286 30252
rect 117685 30243 117743 30249
rect 117685 30209 117697 30243
rect 117731 30240 117743 30243
rect 117774 30240 117780 30252
rect 117731 30212 117780 30240
rect 117731 30209 117743 30212
rect 117685 30203 117743 30209
rect 117774 30200 117780 30212
rect 117832 30200 117838 30252
rect 117976 30249 118004 30280
rect 118510 30268 118516 30320
rect 118568 30268 118574 30320
rect 117869 30243 117927 30249
rect 117869 30209 117881 30243
rect 117915 30209 117927 30243
rect 117869 30203 117927 30209
rect 117961 30243 118019 30249
rect 117961 30209 117973 30243
rect 118007 30209 118019 30243
rect 117961 30203 118019 30209
rect 115308 30144 115980 30172
rect 115952 30113 115980 30144
rect 116026 30132 116032 30184
rect 116084 30172 116090 30184
rect 116596 30172 116624 30200
rect 116964 30172 116992 30200
rect 116084 30144 116624 30172
rect 116780 30144 116992 30172
rect 117884 30172 117912 30203
rect 118050 30200 118056 30252
rect 118108 30240 118114 30252
rect 118237 30243 118295 30249
rect 118237 30240 118249 30243
rect 118108 30212 118249 30240
rect 118108 30200 118114 30212
rect 118237 30209 118249 30212
rect 118283 30209 118295 30243
rect 118237 30203 118295 30209
rect 118068 30172 118096 30200
rect 117884 30144 118096 30172
rect 116084 30132 116090 30144
rect 115937 30107 115995 30113
rect 115124 30076 115704 30104
rect 111150 29996 111156 30048
rect 111208 29996 111214 30048
rect 115382 29996 115388 30048
rect 115440 29996 115446 30048
rect 115676 30045 115704 30076
rect 115937 30073 115949 30107
rect 115983 30073 115995 30107
rect 116780 30104 116808 30144
rect 115937 30067 115995 30073
rect 116136 30076 116808 30104
rect 116136 30048 116164 30076
rect 116854 30064 116860 30116
rect 116912 30104 116918 30116
rect 118145 30107 118203 30113
rect 118145 30104 118157 30107
rect 116912 30076 118157 30104
rect 116912 30064 116918 30076
rect 118145 30073 118157 30076
rect 118191 30073 118203 30107
rect 118145 30067 118203 30073
rect 115661 30039 115719 30045
rect 115661 30005 115673 30039
rect 115707 30036 115719 30039
rect 115750 30036 115756 30048
rect 115707 30008 115756 30036
rect 115707 30005 115719 30008
rect 115661 29999 115719 30005
rect 115750 29996 115756 30008
rect 115808 29996 115814 30048
rect 115842 29996 115848 30048
rect 115900 29996 115906 30048
rect 116118 29996 116124 30048
rect 116176 29996 116182 30048
rect 116578 29996 116584 30048
rect 116636 29996 116642 30048
rect 117406 29996 117412 30048
rect 117464 30036 117470 30048
rect 117501 30039 117559 30045
rect 117501 30036 117513 30039
rect 117464 30008 117513 30036
rect 117464 29996 117470 30008
rect 117501 30005 117513 30008
rect 117547 30005 117559 30039
rect 117501 29999 117559 30005
rect 1104 29946 7912 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 7912 29946
rect 1104 29872 7912 29894
rect 108008 29946 118864 29968
rect 108008 29894 112914 29946
rect 112966 29894 112978 29946
rect 113030 29894 113042 29946
rect 113094 29894 113106 29946
rect 113158 29894 113170 29946
rect 113222 29894 118864 29946
rect 108008 29872 118864 29894
rect 109313 29835 109371 29841
rect 109313 29801 109325 29835
rect 109359 29832 109371 29835
rect 109678 29832 109684 29844
rect 109359 29804 109684 29832
rect 109359 29801 109371 29804
rect 109313 29795 109371 29801
rect 109678 29792 109684 29804
rect 109736 29792 109742 29844
rect 109770 29792 109776 29844
rect 109828 29832 109834 29844
rect 110138 29832 110144 29844
rect 109828 29804 110144 29832
rect 109828 29792 109834 29804
rect 110138 29792 110144 29804
rect 110196 29792 110202 29844
rect 110233 29835 110291 29841
rect 110233 29801 110245 29835
rect 110279 29832 110291 29835
rect 110598 29832 110604 29844
rect 110279 29804 110604 29832
rect 110279 29801 110291 29804
rect 110233 29795 110291 29801
rect 110598 29792 110604 29804
rect 110656 29792 110662 29844
rect 111150 29792 111156 29844
rect 111208 29832 111214 29844
rect 111208 29804 113312 29832
rect 111208 29792 111214 29804
rect 110414 29724 110420 29776
rect 110472 29764 110478 29776
rect 110966 29764 110972 29776
rect 110472 29736 110972 29764
rect 110472 29724 110478 29736
rect 110966 29724 110972 29736
rect 111024 29724 111030 29776
rect 111242 29724 111248 29776
rect 111300 29724 111306 29776
rect 112993 29767 113051 29773
rect 112993 29764 113005 29767
rect 112364 29736 113005 29764
rect 109862 29696 109868 29708
rect 109512 29668 109868 29696
rect 109512 29637 109540 29668
rect 109862 29656 109868 29668
rect 109920 29656 109926 29708
rect 110046 29656 110052 29708
rect 110104 29696 110110 29708
rect 112070 29696 112076 29708
rect 110104 29668 110736 29696
rect 110104 29656 110110 29668
rect 109497 29631 109555 29637
rect 109497 29597 109509 29631
rect 109543 29597 109555 29631
rect 109497 29591 109555 29597
rect 109586 29588 109592 29640
rect 109644 29628 109650 29640
rect 109681 29631 109739 29637
rect 109681 29628 109693 29631
rect 109644 29600 109693 29628
rect 109644 29588 109650 29600
rect 109681 29597 109693 29600
rect 109727 29597 109739 29631
rect 109681 29591 109739 29597
rect 109770 29588 109776 29640
rect 109828 29588 109834 29640
rect 109957 29631 110015 29637
rect 109957 29597 109969 29631
rect 110003 29628 110015 29631
rect 110138 29628 110144 29640
rect 110003 29600 110144 29628
rect 110003 29597 110015 29600
rect 109957 29591 110015 29597
rect 110138 29588 110144 29600
rect 110196 29588 110202 29640
rect 110708 29637 110736 29668
rect 111628 29668 112076 29696
rect 110693 29631 110751 29637
rect 110693 29597 110705 29631
rect 110739 29597 110751 29631
rect 110693 29591 110751 29597
rect 110782 29588 110788 29640
rect 110840 29588 110846 29640
rect 110966 29588 110972 29640
rect 111024 29588 111030 29640
rect 111058 29588 111064 29640
rect 111116 29588 111122 29640
rect 110233 29563 110291 29569
rect 110233 29529 110245 29563
rect 110279 29560 110291 29563
rect 111628 29560 111656 29668
rect 112070 29656 112076 29668
rect 112128 29656 112134 29708
rect 112364 29705 112392 29736
rect 112993 29733 113005 29736
rect 113039 29733 113051 29767
rect 112993 29727 113051 29733
rect 113284 29705 113312 29804
rect 114186 29792 114192 29844
rect 114244 29832 114250 29844
rect 115293 29835 115351 29841
rect 115293 29832 115305 29835
rect 114244 29804 115305 29832
rect 114244 29792 114250 29804
rect 115293 29801 115305 29804
rect 115339 29801 115351 29835
rect 115293 29795 115351 29801
rect 115661 29835 115719 29841
rect 115661 29801 115673 29835
rect 115707 29832 115719 29835
rect 115707 29804 116348 29832
rect 115707 29801 115719 29804
rect 115661 29795 115719 29801
rect 115124 29736 116256 29764
rect 112349 29699 112407 29705
rect 112349 29665 112361 29699
rect 112395 29665 112407 29699
rect 112349 29659 112407 29665
rect 113269 29699 113327 29705
rect 113269 29665 113281 29699
rect 113315 29665 113327 29699
rect 113269 29659 113327 29665
rect 114094 29656 114100 29708
rect 114152 29696 114158 29708
rect 114152 29668 114232 29696
rect 114152 29656 114158 29668
rect 111702 29588 111708 29640
rect 111760 29588 111766 29640
rect 111886 29588 111892 29640
rect 111944 29588 111950 29640
rect 114204 29637 114232 29668
rect 113361 29631 113419 29637
rect 113361 29597 113373 29631
rect 113407 29630 113419 29631
rect 114189 29631 114247 29637
rect 113407 29628 113496 29630
rect 113407 29602 114140 29628
rect 113407 29597 113419 29602
rect 113468 29600 114140 29602
rect 113361 29591 113419 29597
rect 110279 29532 111656 29560
rect 111720 29560 111748 29588
rect 112254 29560 112260 29572
rect 111720 29532 112260 29560
rect 110279 29529 110291 29532
rect 110233 29523 110291 29529
rect 112254 29520 112260 29532
rect 112312 29560 112318 29572
rect 114112 29569 114140 29600
rect 114189 29597 114201 29631
rect 114235 29597 114247 29631
rect 114189 29591 114247 29597
rect 114922 29588 114928 29640
rect 114980 29588 114986 29640
rect 115124 29637 115152 29736
rect 115569 29699 115627 29705
rect 115569 29665 115581 29699
rect 115615 29696 115627 29699
rect 115615 29668 115888 29696
rect 115615 29665 115627 29668
rect 115569 29659 115627 29665
rect 115860 29640 115888 29668
rect 115109 29631 115167 29637
rect 115109 29597 115121 29631
rect 115155 29628 115167 29631
rect 115290 29628 115296 29640
rect 115155 29600 115296 29628
rect 115155 29597 115167 29600
rect 115109 29591 115167 29597
rect 115290 29588 115296 29600
rect 115348 29588 115354 29640
rect 115382 29588 115388 29640
rect 115440 29628 115446 29640
rect 115661 29631 115719 29637
rect 115661 29628 115673 29631
rect 115440 29600 115673 29628
rect 115440 29588 115446 29600
rect 115661 29597 115673 29600
rect 115707 29597 115719 29631
rect 115661 29591 115719 29597
rect 112533 29563 112591 29569
rect 112533 29560 112545 29563
rect 112312 29532 112545 29560
rect 112312 29520 112318 29532
rect 112533 29529 112545 29532
rect 112579 29529 112591 29563
rect 112533 29523 112591 29529
rect 114097 29563 114155 29569
rect 114097 29529 114109 29563
rect 114143 29560 114155 29563
rect 115676 29560 115704 29591
rect 115842 29588 115848 29640
rect 115900 29588 115906 29640
rect 116029 29631 116087 29637
rect 116029 29597 116041 29631
rect 116075 29597 116087 29631
rect 116029 29591 116087 29597
rect 116044 29560 116072 29591
rect 114143 29532 115152 29560
rect 115676 29532 116072 29560
rect 116228 29560 116256 29736
rect 116320 29637 116348 29804
rect 117774 29792 117780 29844
rect 117832 29792 117838 29844
rect 117866 29792 117872 29844
rect 117924 29832 117930 29844
rect 118145 29835 118203 29841
rect 118145 29832 118157 29835
rect 117924 29804 118157 29832
rect 117924 29792 117930 29804
rect 118145 29801 118157 29804
rect 118191 29801 118203 29835
rect 118145 29795 118203 29801
rect 117498 29764 117504 29776
rect 117148 29736 117504 29764
rect 116486 29656 116492 29708
rect 116544 29696 116550 29708
rect 116544 29668 117084 29696
rect 116544 29656 116550 29668
rect 116305 29631 116363 29637
rect 116305 29597 116317 29631
rect 116351 29628 116363 29631
rect 116578 29628 116584 29640
rect 116351 29600 116584 29628
rect 116351 29597 116363 29600
rect 116305 29591 116363 29597
rect 116578 29588 116584 29600
rect 116636 29588 116642 29640
rect 117056 29637 117084 29668
rect 117148 29637 117176 29736
rect 117498 29724 117504 29736
rect 117556 29764 117562 29776
rect 118326 29764 118332 29776
rect 117556 29736 118332 29764
rect 117556 29724 117562 29736
rect 118326 29724 118332 29736
rect 118384 29724 118390 29776
rect 117516 29668 118096 29696
rect 117041 29631 117099 29637
rect 117041 29597 117053 29631
rect 117087 29597 117099 29631
rect 117041 29591 117099 29597
rect 117133 29631 117191 29637
rect 117133 29597 117145 29631
rect 117179 29597 117191 29631
rect 117133 29591 117191 29597
rect 116762 29560 116768 29572
rect 116228 29532 116768 29560
rect 114143 29529 114155 29532
rect 114097 29523 114155 29529
rect 115124 29504 115152 29532
rect 116762 29520 116768 29532
rect 116820 29520 116826 29572
rect 116949 29563 117007 29569
rect 116949 29529 116961 29563
rect 116995 29560 117007 29563
rect 117516 29560 117544 29668
rect 118068 29640 118096 29668
rect 117590 29588 117596 29640
rect 117648 29588 117654 29640
rect 118050 29588 118056 29640
rect 118108 29588 118114 29640
rect 118510 29588 118516 29640
rect 118568 29588 118574 29640
rect 116995 29532 117544 29560
rect 117608 29560 117636 29588
rect 117774 29569 117780 29572
rect 117745 29563 117780 29569
rect 117745 29560 117757 29563
rect 117608 29532 117757 29560
rect 116995 29529 117007 29532
rect 116949 29523 117007 29529
rect 117745 29529 117757 29532
rect 117745 29523 117780 29529
rect 117774 29520 117780 29523
rect 117832 29520 117838 29572
rect 117958 29520 117964 29572
rect 118016 29520 118022 29572
rect 110046 29452 110052 29504
rect 110104 29452 110110 29504
rect 111889 29495 111947 29501
rect 111889 29461 111901 29495
rect 111935 29492 111947 29495
rect 112441 29495 112499 29501
rect 112441 29492 112453 29495
rect 111935 29464 112453 29492
rect 111935 29461 111947 29464
rect 111889 29455 111947 29461
rect 112441 29461 112453 29464
rect 112487 29461 112499 29495
rect 112441 29455 112499 29461
rect 112806 29452 112812 29504
rect 112864 29492 112870 29504
rect 112901 29495 112959 29501
rect 112901 29492 112913 29495
rect 112864 29464 112913 29492
rect 112864 29452 112870 29464
rect 112901 29461 112913 29464
rect 112947 29461 112959 29495
rect 112901 29455 112959 29461
rect 114738 29452 114744 29504
rect 114796 29492 114802 29504
rect 114925 29495 114983 29501
rect 114925 29492 114937 29495
rect 114796 29464 114937 29492
rect 114796 29452 114802 29464
rect 114925 29461 114937 29464
rect 114971 29461 114983 29495
rect 114925 29455 114983 29461
rect 115106 29452 115112 29504
rect 115164 29452 115170 29504
rect 115934 29452 115940 29504
rect 115992 29492 115998 29504
rect 116489 29495 116547 29501
rect 116489 29492 116501 29495
rect 115992 29464 116501 29492
rect 115992 29452 115998 29464
rect 116489 29461 116501 29464
rect 116535 29461 116547 29495
rect 116489 29455 116547 29461
rect 116854 29452 116860 29504
rect 116912 29452 116918 29504
rect 117314 29452 117320 29504
rect 117372 29492 117378 29504
rect 117498 29492 117504 29504
rect 117372 29464 117504 29492
rect 117372 29452 117378 29464
rect 117498 29452 117504 29464
rect 117556 29452 117562 29504
rect 117590 29452 117596 29504
rect 117648 29452 117654 29504
rect 118142 29452 118148 29504
rect 118200 29492 118206 29504
rect 118329 29495 118387 29501
rect 118329 29492 118341 29495
rect 118200 29464 118341 29492
rect 118200 29452 118206 29464
rect 118329 29461 118341 29464
rect 118375 29461 118387 29495
rect 118329 29455 118387 29461
rect 1104 29402 7912 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 7912 29402
rect 1104 29328 7912 29350
rect 108008 29402 118864 29424
rect 108008 29350 113650 29402
rect 113702 29350 113714 29402
rect 113766 29350 113778 29402
rect 113830 29350 113842 29402
rect 113894 29350 113906 29402
rect 113958 29350 118864 29402
rect 108008 29328 118864 29350
rect 109586 29248 109592 29300
rect 109644 29248 109650 29300
rect 109681 29291 109739 29297
rect 109681 29257 109693 29291
rect 109727 29288 109739 29291
rect 109862 29288 109868 29300
rect 109727 29260 109868 29288
rect 109727 29257 109739 29260
rect 109681 29251 109739 29257
rect 109862 29248 109868 29260
rect 109920 29248 109926 29300
rect 110138 29248 110144 29300
rect 110196 29288 110202 29300
rect 110322 29288 110328 29300
rect 110196 29260 110328 29288
rect 110196 29248 110202 29260
rect 110322 29248 110328 29260
rect 110380 29248 110386 29300
rect 110601 29291 110659 29297
rect 110601 29257 110613 29291
rect 110647 29288 110659 29291
rect 110782 29288 110788 29300
rect 110647 29260 110788 29288
rect 110647 29257 110659 29260
rect 110601 29251 110659 29257
rect 110782 29248 110788 29260
rect 110840 29248 110846 29300
rect 113358 29248 113364 29300
rect 113416 29288 113422 29300
rect 116210 29288 116216 29300
rect 113416 29260 113956 29288
rect 113416 29248 113422 29260
rect 109770 29180 109776 29232
rect 109828 29220 109834 29232
rect 110233 29223 110291 29229
rect 110233 29220 110245 29223
rect 109828 29192 110245 29220
rect 109828 29180 109834 29192
rect 110233 29189 110245 29192
rect 110279 29189 110291 29223
rect 110340 29220 110368 29248
rect 110449 29223 110507 29229
rect 110449 29220 110461 29223
rect 110340 29192 110461 29220
rect 110233 29183 110291 29189
rect 110449 29189 110461 29192
rect 110495 29220 110507 29223
rect 110495 29192 111196 29220
rect 110495 29189 110507 29192
rect 110449 29183 110507 29189
rect 109405 29155 109463 29161
rect 109405 29121 109417 29155
rect 109451 29121 109463 29155
rect 109405 29115 109463 29121
rect 109589 29155 109647 29161
rect 109589 29121 109601 29155
rect 109635 29152 109647 29155
rect 109865 29155 109923 29161
rect 109635 29124 109816 29152
rect 109635 29121 109647 29124
rect 109589 29115 109647 29121
rect 109420 29084 109448 29115
rect 109678 29084 109684 29096
rect 109420 29056 109684 29084
rect 109678 29044 109684 29056
rect 109736 29044 109742 29096
rect 109788 28948 109816 29124
rect 109865 29121 109877 29155
rect 109911 29121 109923 29155
rect 109865 29115 109923 29121
rect 110049 29155 110107 29161
rect 110049 29121 110061 29155
rect 110095 29121 110107 29155
rect 110049 29115 110107 29121
rect 109880 29016 109908 29115
rect 110064 29084 110092 29115
rect 110138 29112 110144 29164
rect 110196 29112 110202 29164
rect 110248 29152 110276 29183
rect 110598 29152 110604 29164
rect 110248 29124 110604 29152
rect 110598 29112 110604 29124
rect 110656 29112 110662 29164
rect 110414 29084 110420 29096
rect 110064 29056 110420 29084
rect 110414 29044 110420 29056
rect 110472 29044 110478 29096
rect 110969 29019 111027 29025
rect 110969 29016 110981 29019
rect 109880 28988 110981 29016
rect 110969 28985 110981 28988
rect 111015 29016 111027 29019
rect 111058 29016 111064 29028
rect 111015 28988 111064 29016
rect 111015 28985 111027 28988
rect 110969 28979 111027 28985
rect 111058 28976 111064 28988
rect 111116 28976 111122 29028
rect 111168 29016 111196 29192
rect 113450 29180 113456 29232
rect 113508 29220 113514 29232
rect 113508 29192 113772 29220
rect 113508 29180 113514 29192
rect 113744 29164 113772 29192
rect 113928 29167 113956 29260
rect 115952 29260 116216 29288
rect 115017 29223 115075 29229
rect 115017 29189 115029 29223
rect 115063 29220 115075 29223
rect 115569 29223 115627 29229
rect 115569 29220 115581 29223
rect 115063 29192 115581 29220
rect 115063 29189 115075 29192
rect 115017 29183 115075 29189
rect 115569 29189 115581 29192
rect 115615 29189 115627 29223
rect 115952 29220 115980 29260
rect 116210 29248 116216 29260
rect 116268 29288 116274 29300
rect 116946 29288 116952 29300
rect 116268 29260 116952 29288
rect 116268 29248 116274 29260
rect 116946 29248 116952 29260
rect 117004 29248 117010 29300
rect 117406 29248 117412 29300
rect 117464 29288 117470 29300
rect 117464 29260 117820 29288
rect 117464 29248 117470 29260
rect 116854 29220 116860 29232
rect 115569 29183 115627 29189
rect 115860 29192 115980 29220
rect 116044 29192 116860 29220
rect 111334 29112 111340 29164
rect 111392 29112 111398 29164
rect 113545 29155 113603 29161
rect 113545 29121 113557 29155
rect 113591 29121 113603 29155
rect 113545 29115 113603 29121
rect 111429 29087 111487 29093
rect 111429 29053 111441 29087
rect 111475 29084 111487 29087
rect 111978 29084 111984 29096
rect 111475 29056 111984 29084
rect 111475 29053 111487 29056
rect 111429 29047 111487 29053
rect 111978 29044 111984 29056
rect 112036 29044 112042 29096
rect 111794 29016 111800 29028
rect 111168 28988 111800 29016
rect 111794 28976 111800 28988
rect 111852 29016 111858 29028
rect 113361 29019 113419 29025
rect 113361 29016 113373 29019
rect 111852 28988 113373 29016
rect 111852 28976 111858 28988
rect 113361 28985 113373 28988
rect 113407 28985 113419 29019
rect 113560 29016 113588 29115
rect 113726 29112 113732 29164
rect 113784 29112 113790 29164
rect 113914 29161 113972 29167
rect 113914 29127 113926 29161
rect 113960 29127 113972 29161
rect 113914 29121 113972 29127
rect 114097 29155 114155 29161
rect 114097 29121 114109 29155
rect 114143 29152 114155 29155
rect 114186 29152 114192 29164
rect 114143 29124 114192 29152
rect 114143 29121 114155 29124
rect 114097 29115 114155 29121
rect 114186 29112 114192 29124
rect 114244 29112 114250 29164
rect 114922 29112 114928 29164
rect 114980 29112 114986 29164
rect 115106 29112 115112 29164
rect 115164 29112 115170 29164
rect 115293 29155 115351 29161
rect 115293 29121 115305 29155
rect 115339 29121 115351 29155
rect 115293 29115 115351 29121
rect 115385 29155 115443 29161
rect 115385 29121 115397 29155
rect 115431 29121 115443 29155
rect 115385 29115 115443 29121
rect 113821 29087 113879 29093
rect 113821 29053 113833 29087
rect 113867 29084 113879 29087
rect 114002 29084 114008 29096
rect 113867 29056 114008 29084
rect 113867 29053 113879 29056
rect 113821 29047 113879 29053
rect 114002 29044 114008 29056
rect 114060 29044 114066 29096
rect 114741 29019 114799 29025
rect 114741 29016 114753 29019
rect 113560 28988 114753 29016
rect 113361 28979 113419 28985
rect 114741 28985 114753 28988
rect 114787 29016 114799 29019
rect 115106 29016 115112 29028
rect 114787 28988 115112 29016
rect 114787 28985 114799 28988
rect 114741 28979 114799 28985
rect 115106 28976 115112 28988
rect 115164 28976 115170 29028
rect 115308 29016 115336 29115
rect 115400 29084 115428 29115
rect 115474 29112 115480 29164
rect 115532 29112 115538 29164
rect 115860 29161 115888 29192
rect 115661 29155 115719 29161
rect 115661 29121 115673 29155
rect 115707 29152 115719 29155
rect 115845 29155 115903 29161
rect 115845 29152 115857 29155
rect 115707 29124 115857 29152
rect 115707 29121 115719 29124
rect 115661 29115 115719 29121
rect 115845 29121 115857 29124
rect 115891 29121 115903 29155
rect 115845 29115 115903 29121
rect 115934 29112 115940 29164
rect 115992 29112 115998 29164
rect 116044 29161 116072 29192
rect 116854 29180 116860 29192
rect 116912 29180 116918 29232
rect 117225 29223 117283 29229
rect 117225 29189 117237 29223
rect 117271 29220 117283 29223
rect 117590 29220 117596 29232
rect 117271 29192 117596 29220
rect 117271 29189 117283 29192
rect 117225 29183 117283 29189
rect 117590 29180 117596 29192
rect 117648 29220 117654 29232
rect 117685 29223 117743 29229
rect 117685 29220 117697 29223
rect 117648 29192 117697 29220
rect 117648 29180 117654 29192
rect 117685 29189 117697 29192
rect 117731 29189 117743 29223
rect 117685 29183 117743 29189
rect 116029 29155 116087 29161
rect 116029 29121 116041 29155
rect 116075 29121 116087 29155
rect 116029 29115 116087 29121
rect 116121 29155 116179 29161
rect 116121 29121 116133 29155
rect 116167 29152 116179 29155
rect 116397 29155 116455 29161
rect 116397 29152 116409 29155
rect 116167 29124 116409 29152
rect 116167 29121 116179 29124
rect 116121 29115 116179 29121
rect 116397 29121 116409 29124
rect 116443 29121 116455 29155
rect 116397 29115 116455 29121
rect 115952 29084 115980 29112
rect 115400 29056 115980 29084
rect 116044 29016 116072 29115
rect 115308 28988 116072 29016
rect 110414 28948 110420 28960
rect 109788 28920 110420 28948
rect 110414 28908 110420 28920
rect 110472 28908 110478 28960
rect 115474 28908 115480 28960
rect 115532 28948 115538 28960
rect 116136 28948 116164 29115
rect 116412 29084 116440 29115
rect 116486 29112 116492 29164
rect 116544 29112 116550 29164
rect 116673 29155 116731 29161
rect 116673 29121 116685 29155
rect 116719 29152 116731 29155
rect 116762 29152 116768 29164
rect 116719 29124 116768 29152
rect 116719 29121 116731 29124
rect 116673 29115 116731 29121
rect 116762 29112 116768 29124
rect 116820 29112 116826 29164
rect 116949 29155 117007 29161
rect 116949 29121 116961 29155
rect 116995 29152 117007 29155
rect 117314 29152 117320 29164
rect 116995 29124 117320 29152
rect 116995 29121 117007 29124
rect 116949 29115 117007 29121
rect 117314 29112 117320 29124
rect 117372 29112 117378 29164
rect 117501 29155 117559 29161
rect 117501 29121 117513 29155
rect 117547 29152 117559 29155
rect 117547 29124 117636 29152
rect 117547 29121 117559 29124
rect 117501 29115 117559 29121
rect 117608 29096 117636 29124
rect 117406 29084 117412 29096
rect 116412 29056 117412 29084
rect 117406 29044 117412 29056
rect 117464 29044 117470 29096
rect 117590 29044 117596 29096
rect 117648 29044 117654 29096
rect 117133 29019 117191 29025
rect 117133 28985 117145 29019
rect 117179 29016 117191 29019
rect 117682 29016 117688 29028
rect 117179 28988 117688 29016
rect 117179 28985 117191 28988
rect 117133 28979 117191 28985
rect 117682 28976 117688 28988
rect 117740 28976 117746 29028
rect 117792 29016 117820 29260
rect 117961 29019 118019 29025
rect 117961 29016 117973 29019
rect 117792 28988 117973 29016
rect 117961 28985 117973 28988
rect 118007 28985 118019 29019
rect 117961 28979 118019 28985
rect 118142 28976 118148 29028
rect 118200 28976 118206 29028
rect 118510 28976 118516 29028
rect 118568 28976 118574 29028
rect 115532 28920 116164 28948
rect 116305 28951 116363 28957
rect 115532 28908 115538 28920
rect 116305 28917 116317 28951
rect 116351 28948 116363 28951
rect 116670 28948 116676 28960
rect 116351 28920 116676 28948
rect 116351 28917 116363 28920
rect 116305 28911 116363 28917
rect 116670 28908 116676 28920
rect 116728 28908 116734 28960
rect 116854 28908 116860 28960
rect 116912 28908 116918 28960
rect 116946 28908 116952 28960
rect 117004 28948 117010 28960
rect 117225 28951 117283 28957
rect 117225 28948 117237 28951
rect 117004 28920 117237 28948
rect 117004 28908 117010 28920
rect 117225 28917 117237 28920
rect 117271 28917 117283 28951
rect 117225 28911 117283 28917
rect 1104 28858 7912 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 7912 28858
rect 1104 28784 7912 28806
rect 108008 28858 118864 28880
rect 108008 28806 112914 28858
rect 112966 28806 112978 28858
rect 113030 28806 113042 28858
rect 113094 28806 113106 28858
rect 113158 28806 113170 28858
rect 113222 28806 118864 28858
rect 108008 28784 118864 28806
rect 110046 28704 110052 28756
rect 110104 28744 110110 28756
rect 110233 28747 110291 28753
rect 110233 28744 110245 28747
rect 110104 28716 110245 28744
rect 110104 28704 110110 28716
rect 110233 28713 110245 28716
rect 110279 28713 110291 28747
rect 110233 28707 110291 28713
rect 111061 28747 111119 28753
rect 111061 28713 111073 28747
rect 111107 28744 111119 28747
rect 111702 28744 111708 28756
rect 111107 28716 111708 28744
rect 111107 28713 111119 28716
rect 111061 28707 111119 28713
rect 109770 28568 109776 28620
rect 109828 28608 109834 28620
rect 110138 28608 110144 28620
rect 109828 28580 110144 28608
rect 109828 28568 109834 28580
rect 109862 28500 109868 28552
rect 109920 28500 109926 28552
rect 109972 28549 110000 28580
rect 110138 28568 110144 28580
rect 110196 28568 110202 28620
rect 110248 28608 110276 28707
rect 111702 28704 111708 28716
rect 111760 28704 111766 28756
rect 111978 28704 111984 28756
rect 112036 28704 112042 28756
rect 112438 28704 112444 28756
rect 112496 28744 112502 28756
rect 112993 28747 113051 28753
rect 112993 28744 113005 28747
rect 112496 28716 113005 28744
rect 112496 28704 112502 28716
rect 112993 28713 113005 28716
rect 113039 28744 113051 28747
rect 113450 28744 113456 28756
rect 113039 28716 113456 28744
rect 113039 28713 113051 28716
rect 112993 28707 113051 28713
rect 113450 28704 113456 28716
rect 113508 28704 113514 28756
rect 113726 28704 113732 28756
rect 113784 28744 113790 28756
rect 114005 28747 114063 28753
rect 114005 28744 114017 28747
rect 113784 28716 114017 28744
rect 113784 28704 113790 28716
rect 114005 28713 114017 28716
rect 114051 28744 114063 28747
rect 114094 28744 114100 28756
rect 114051 28716 114100 28744
rect 114051 28713 114063 28716
rect 114005 28707 114063 28713
rect 114094 28704 114100 28716
rect 114152 28704 114158 28756
rect 114922 28704 114928 28756
rect 114980 28744 114986 28756
rect 115845 28747 115903 28753
rect 115845 28744 115857 28747
rect 114980 28716 115857 28744
rect 114980 28704 114986 28716
rect 115845 28713 115857 28716
rect 115891 28713 115903 28747
rect 115845 28707 115903 28713
rect 118050 28704 118056 28756
rect 118108 28704 118114 28756
rect 110598 28636 110604 28688
rect 110656 28676 110662 28688
rect 112533 28679 112591 28685
rect 112533 28676 112545 28679
rect 110656 28648 112545 28676
rect 110656 28636 110662 28648
rect 112533 28645 112545 28648
rect 112579 28645 112591 28679
rect 112533 28639 112591 28645
rect 113269 28679 113327 28685
rect 113269 28645 113281 28679
rect 113315 28645 113327 28679
rect 115934 28676 115940 28688
rect 113269 28639 113327 28645
rect 113376 28648 115940 28676
rect 110693 28611 110751 28617
rect 110693 28608 110705 28611
rect 110248 28580 110705 28608
rect 110693 28577 110705 28580
rect 110739 28577 110751 28611
rect 113284 28608 113312 28639
rect 110693 28571 110751 28577
rect 112180 28580 113312 28608
rect 109957 28543 110015 28549
rect 109957 28509 109969 28543
rect 110003 28509 110015 28543
rect 109957 28503 110015 28509
rect 110049 28543 110107 28549
rect 110049 28509 110061 28543
rect 110095 28509 110107 28543
rect 110049 28503 110107 28509
rect 110064 28472 110092 28503
rect 110230 28500 110236 28552
rect 110288 28540 110294 28552
rect 112180 28549 112208 28580
rect 110877 28543 110935 28549
rect 110877 28540 110889 28543
rect 110288 28512 110889 28540
rect 110288 28500 110294 28512
rect 110877 28509 110889 28512
rect 110923 28509 110935 28543
rect 110877 28503 110935 28509
rect 112165 28543 112223 28549
rect 112165 28509 112177 28543
rect 112211 28540 112223 28543
rect 112254 28540 112260 28552
rect 112211 28512 112260 28540
rect 112211 28509 112223 28512
rect 112165 28503 112223 28509
rect 112254 28500 112260 28512
rect 112312 28500 112318 28552
rect 112438 28500 112444 28552
rect 112496 28500 112502 28552
rect 112625 28543 112683 28549
rect 112625 28509 112637 28543
rect 112671 28540 112683 28543
rect 113376 28540 113404 28648
rect 115934 28636 115940 28648
rect 115992 28676 115998 28688
rect 116118 28676 116124 28688
rect 115992 28648 116124 28676
rect 115992 28636 115998 28648
rect 116118 28636 116124 28648
rect 116176 28636 116182 28688
rect 114204 28580 114508 28608
rect 112671 28512 112944 28540
rect 112671 28509 112683 28512
rect 112625 28503 112683 28509
rect 110414 28472 110420 28484
rect 110064 28444 110420 28472
rect 110414 28432 110420 28444
rect 110472 28472 110478 28484
rect 110782 28472 110788 28484
rect 110472 28444 110788 28472
rect 110472 28432 110478 28444
rect 110782 28432 110788 28444
rect 110840 28432 110846 28484
rect 112349 28475 112407 28481
rect 112349 28441 112361 28475
rect 112395 28472 112407 28475
rect 112395 28444 112852 28472
rect 112395 28441 112407 28444
rect 112349 28435 112407 28441
rect 112622 28364 112628 28416
rect 112680 28404 112686 28416
rect 112824 28413 112852 28444
rect 112809 28407 112867 28413
rect 112809 28404 112821 28407
rect 112680 28376 112821 28404
rect 112680 28364 112686 28376
rect 112809 28373 112821 28376
rect 112855 28373 112867 28407
rect 112916 28404 112944 28512
rect 113284 28512 113404 28540
rect 113284 28481 113312 28512
rect 113542 28500 113548 28552
rect 113600 28500 113606 28552
rect 114204 28549 114232 28580
rect 114480 28552 114508 28580
rect 114738 28568 114744 28620
rect 114796 28568 114802 28620
rect 114830 28568 114836 28620
rect 114888 28568 114894 28620
rect 115014 28568 115020 28620
rect 115072 28608 115078 28620
rect 115474 28608 115480 28620
rect 115072 28580 115480 28608
rect 115072 28568 115078 28580
rect 115474 28568 115480 28580
rect 115532 28608 115538 28620
rect 117041 28611 117099 28617
rect 115532 28580 116072 28608
rect 115532 28568 115538 28580
rect 114189 28543 114247 28549
rect 114189 28509 114201 28543
rect 114235 28509 114247 28543
rect 114189 28503 114247 28509
rect 114370 28500 114376 28552
rect 114428 28500 114434 28552
rect 114462 28500 114468 28552
rect 114520 28540 114526 28552
rect 114649 28543 114707 28549
rect 114649 28540 114661 28543
rect 114520 28512 114661 28540
rect 114520 28500 114526 28512
rect 114649 28509 114661 28512
rect 114695 28509 114707 28543
rect 114649 28503 114707 28509
rect 114925 28543 114983 28549
rect 114925 28509 114937 28543
rect 114971 28509 114983 28543
rect 114925 28503 114983 28509
rect 113177 28475 113235 28481
rect 113177 28441 113189 28475
rect 113223 28472 113235 28475
rect 113269 28475 113327 28481
rect 113269 28472 113281 28475
rect 113223 28444 113281 28472
rect 113223 28441 113235 28444
rect 113177 28435 113235 28441
rect 113269 28441 113281 28444
rect 113315 28441 113327 28475
rect 113269 28435 113327 28441
rect 113450 28432 113456 28484
rect 113508 28472 113514 28484
rect 114940 28472 114968 28503
rect 115106 28500 115112 28552
rect 115164 28500 115170 28552
rect 115290 28500 115296 28552
rect 115348 28500 115354 28552
rect 116044 28549 116072 28580
rect 117041 28577 117053 28611
rect 117087 28608 117099 28611
rect 117087 28580 118556 28608
rect 117087 28577 117099 28580
rect 117041 28571 117099 28577
rect 116029 28543 116087 28549
rect 116029 28509 116041 28543
rect 116075 28509 116087 28543
rect 116029 28503 116087 28509
rect 116210 28500 116216 28552
rect 116268 28500 116274 28552
rect 117130 28500 117136 28552
rect 117188 28540 117194 28552
rect 117409 28543 117467 28549
rect 117409 28540 117421 28543
rect 117188 28512 117421 28540
rect 117188 28500 117194 28512
rect 117409 28509 117421 28512
rect 117455 28509 117467 28543
rect 117409 28503 117467 28509
rect 117685 28543 117743 28549
rect 117685 28509 117697 28543
rect 117731 28540 117743 28543
rect 117774 28540 117780 28552
rect 117731 28512 117780 28540
rect 117731 28509 117743 28512
rect 117685 28503 117743 28509
rect 117774 28500 117780 28512
rect 117832 28500 117838 28552
rect 117869 28543 117927 28549
rect 117869 28509 117881 28543
rect 117915 28509 117927 28543
rect 117869 28503 117927 28509
rect 113508 28444 114508 28472
rect 114940 28444 115612 28472
rect 113508 28432 113514 28444
rect 112977 28407 113035 28413
rect 112977 28404 112989 28407
rect 112916 28376 112989 28404
rect 112809 28367 112867 28373
rect 112977 28373 112989 28376
rect 113023 28404 113035 28407
rect 113542 28404 113548 28416
rect 113023 28376 113548 28404
rect 113023 28373 113035 28376
rect 112977 28367 113035 28373
rect 113542 28364 113548 28376
rect 113600 28364 113606 28416
rect 114480 28413 114508 28444
rect 115584 28416 115612 28444
rect 117038 28432 117044 28484
rect 117096 28472 117102 28484
rect 117225 28475 117283 28481
rect 117225 28472 117237 28475
rect 117096 28444 117237 28472
rect 117096 28432 117102 28444
rect 117225 28441 117237 28444
rect 117271 28441 117283 28475
rect 117884 28472 117912 28503
rect 118234 28500 118240 28552
rect 118292 28500 118298 28552
rect 118528 28549 118556 28580
rect 118513 28543 118571 28549
rect 118513 28509 118525 28543
rect 118559 28540 118571 28543
rect 118602 28540 118608 28552
rect 118559 28512 118608 28540
rect 118559 28509 118571 28512
rect 118513 28503 118571 28509
rect 118602 28500 118608 28512
rect 118660 28500 118666 28552
rect 117958 28472 117964 28484
rect 117884 28444 117964 28472
rect 117225 28435 117283 28441
rect 117958 28432 117964 28444
rect 118016 28472 118022 28484
rect 118016 28444 118372 28472
rect 118016 28432 118022 28444
rect 114465 28407 114523 28413
rect 114465 28373 114477 28407
rect 114511 28373 114523 28407
rect 114465 28367 114523 28373
rect 114922 28364 114928 28416
rect 114980 28404 114986 28416
rect 115201 28407 115259 28413
rect 115201 28404 115213 28407
rect 114980 28376 115213 28404
rect 114980 28364 114986 28376
rect 115201 28373 115213 28376
rect 115247 28373 115259 28407
rect 115201 28367 115259 28373
rect 115566 28364 115572 28416
rect 115624 28404 115630 28416
rect 116946 28404 116952 28416
rect 115624 28376 116952 28404
rect 115624 28364 115630 28376
rect 116946 28364 116952 28376
rect 117004 28364 117010 28416
rect 117590 28364 117596 28416
rect 117648 28364 117654 28416
rect 117774 28364 117780 28416
rect 117832 28364 117838 28416
rect 118344 28413 118372 28444
rect 118329 28407 118387 28413
rect 118329 28373 118341 28407
rect 118375 28373 118387 28407
rect 118329 28367 118387 28373
rect 1104 28314 7912 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 7912 28314
rect 1104 28240 7912 28262
rect 108008 28314 118864 28336
rect 108008 28262 113650 28314
rect 113702 28262 113714 28314
rect 113766 28262 113778 28314
rect 113830 28262 113842 28314
rect 113894 28262 113906 28314
rect 113958 28262 118864 28314
rect 108008 28240 118864 28262
rect 109589 28203 109647 28209
rect 109589 28169 109601 28203
rect 109635 28200 109647 28203
rect 110230 28200 110236 28212
rect 109635 28172 110236 28200
rect 109635 28169 109647 28172
rect 109589 28163 109647 28169
rect 110230 28160 110236 28172
rect 110288 28160 110294 28212
rect 113358 28160 113364 28212
rect 113416 28200 113422 28212
rect 113453 28203 113511 28209
rect 113453 28200 113465 28203
rect 113416 28172 113465 28200
rect 113416 28160 113422 28172
rect 113453 28169 113465 28172
rect 113499 28169 113511 28203
rect 113453 28163 113511 28169
rect 113542 28160 113548 28212
rect 113600 28200 113606 28212
rect 114281 28203 114339 28209
rect 114281 28200 114293 28203
rect 113600 28172 114293 28200
rect 113600 28160 113606 28172
rect 114281 28169 114293 28172
rect 114327 28169 114339 28203
rect 114281 28163 114339 28169
rect 114370 28160 114376 28212
rect 114428 28200 114434 28212
rect 116026 28200 116032 28212
rect 114428 28172 116032 28200
rect 114428 28160 114434 28172
rect 112346 28132 112352 28144
rect 111628 28104 112352 28132
rect 109770 28024 109776 28076
rect 109828 28024 109834 28076
rect 109865 28067 109923 28073
rect 109865 28033 109877 28067
rect 109911 28033 109923 28067
rect 109865 28027 109923 28033
rect 109880 27996 109908 28027
rect 109954 28024 109960 28076
rect 110012 28024 110018 28076
rect 110141 28067 110199 28073
rect 110141 28033 110153 28067
rect 110187 28064 110199 28067
rect 111058 28064 111064 28076
rect 110187 28036 111064 28064
rect 110187 28033 110199 28036
rect 110141 28027 110199 28033
rect 111058 28024 111064 28036
rect 111116 28024 111122 28076
rect 111628 28073 111656 28104
rect 112346 28092 112352 28104
rect 112404 28132 112410 28144
rect 113376 28132 113404 28160
rect 112404 28104 113404 28132
rect 113913 28135 113971 28141
rect 112404 28092 112410 28104
rect 113913 28101 113925 28135
rect 113959 28132 113971 28135
rect 114002 28132 114008 28144
rect 113959 28104 114008 28132
rect 113959 28101 113971 28104
rect 113913 28095 113971 28101
rect 114002 28092 114008 28104
rect 114060 28092 114066 28144
rect 114738 28132 114744 28144
rect 114664 28104 114744 28132
rect 111613 28067 111671 28073
rect 111613 28033 111625 28067
rect 111659 28033 111671 28067
rect 111613 28027 111671 28033
rect 111702 28024 111708 28076
rect 111760 28024 111766 28076
rect 112254 28024 112260 28076
rect 112312 28024 112318 28076
rect 112533 28067 112591 28073
rect 112533 28033 112545 28067
rect 112579 28064 112591 28067
rect 112622 28064 112628 28076
rect 112579 28036 112628 28064
rect 112579 28033 112591 28036
rect 112533 28027 112591 28033
rect 112622 28024 112628 28036
rect 112680 28024 112686 28076
rect 112717 28067 112775 28073
rect 112717 28033 112729 28067
rect 112763 28033 112775 28067
rect 112717 28027 112775 28033
rect 110782 27996 110788 28008
rect 109880 27968 110788 27996
rect 110782 27956 110788 27968
rect 110840 27996 110846 28008
rect 111245 27999 111303 28005
rect 111245 27996 111257 27999
rect 110840 27968 111257 27996
rect 110840 27956 110846 27968
rect 111245 27965 111257 27968
rect 111291 27965 111303 27999
rect 111245 27959 111303 27965
rect 112732 27928 112760 28027
rect 113266 28024 113272 28076
rect 113324 28064 113330 28076
rect 113821 28067 113879 28073
rect 113821 28064 113833 28067
rect 113324 28036 113833 28064
rect 113324 28024 113330 28036
rect 113821 28033 113833 28036
rect 113867 28064 113879 28067
rect 113867 28036 114416 28064
rect 113867 28033 113879 28036
rect 113821 28027 113879 28033
rect 114094 27956 114100 28008
rect 114152 27956 114158 28008
rect 114388 27996 114416 28036
rect 114462 28024 114468 28076
rect 114520 28024 114526 28076
rect 114554 28024 114560 28076
rect 114612 28024 114618 28076
rect 114664 28073 114692 28104
rect 114738 28092 114744 28104
rect 114796 28132 114802 28144
rect 115661 28135 115719 28141
rect 115661 28132 115673 28135
rect 114796 28104 115673 28132
rect 114796 28092 114802 28104
rect 115661 28101 115673 28104
rect 115707 28101 115719 28135
rect 115661 28095 115719 28101
rect 114649 28067 114707 28073
rect 114649 28033 114661 28067
rect 114695 28033 114707 28067
rect 114649 28027 114707 28033
rect 114830 28024 114836 28076
rect 114888 28024 114894 28076
rect 115017 28067 115075 28073
rect 115017 28033 115029 28067
rect 115063 28033 115075 28067
rect 115017 28027 115075 28033
rect 115032 27996 115060 28027
rect 115566 28024 115572 28076
rect 115624 28024 115630 28076
rect 115768 28073 115796 28172
rect 116026 28160 116032 28172
rect 116084 28160 116090 28212
rect 116578 28160 116584 28212
rect 116636 28200 116642 28212
rect 117317 28203 117375 28209
rect 116636 28172 117176 28200
rect 116636 28160 116642 28172
rect 117148 28144 117176 28172
rect 117317 28169 117329 28203
rect 117363 28200 117375 28203
rect 117774 28200 117780 28212
rect 117363 28172 117780 28200
rect 117363 28169 117375 28172
rect 117317 28163 117375 28169
rect 117774 28160 117780 28172
rect 117832 28160 117838 28212
rect 118053 28203 118111 28209
rect 118053 28169 118065 28203
rect 118099 28169 118111 28203
rect 118053 28163 118111 28169
rect 116412 28104 116900 28132
rect 115753 28067 115811 28073
rect 115753 28033 115765 28067
rect 115799 28033 115811 28067
rect 115753 28027 115811 28033
rect 116118 28024 116124 28076
rect 116176 28024 116182 28076
rect 116412 28073 116440 28104
rect 116872 28076 116900 28104
rect 117130 28092 117136 28144
rect 117188 28132 117194 28144
rect 118068 28132 118096 28163
rect 118234 28160 118240 28212
rect 118292 28200 118298 28212
rect 118421 28203 118479 28209
rect 118421 28200 118433 28203
rect 118292 28172 118433 28200
rect 118292 28160 118298 28172
rect 118421 28169 118433 28172
rect 118467 28169 118479 28203
rect 118421 28163 118479 28169
rect 117188 28104 118096 28132
rect 117188 28092 117194 28104
rect 116397 28067 116455 28073
rect 116397 28033 116409 28067
rect 116443 28033 116455 28067
rect 116397 28027 116455 28033
rect 116578 28024 116584 28076
rect 116636 28024 116642 28076
rect 116670 28024 116676 28076
rect 116728 28024 116734 28076
rect 116854 28024 116860 28076
rect 116912 28024 116918 28076
rect 116946 28024 116952 28076
rect 117004 28064 117010 28076
rect 117004 28036 117636 28064
rect 117004 28024 117010 28036
rect 114388 27968 115060 27996
rect 114370 27928 114376 27940
rect 112732 27900 114376 27928
rect 114370 27888 114376 27900
rect 114428 27888 114434 27940
rect 115032 27928 115060 27968
rect 116259 27999 116317 28005
rect 116259 27965 116271 27999
rect 116305 27996 116317 27999
rect 116688 27996 116716 28024
rect 116305 27968 116716 27996
rect 116305 27965 116317 27968
rect 116259 27959 116317 27965
rect 117406 27956 117412 28008
rect 117464 27956 117470 28008
rect 117501 27999 117559 28005
rect 117501 27965 117513 27999
rect 117547 27965 117559 27999
rect 117608 27996 117636 28036
rect 117682 28024 117688 28076
rect 117740 28064 117746 28076
rect 117777 28067 117835 28073
rect 117777 28064 117789 28067
rect 117740 28036 117789 28064
rect 117740 28024 117746 28036
rect 117777 28033 117789 28036
rect 117823 28033 117835 28067
rect 117777 28027 117835 28033
rect 118234 28024 118240 28076
rect 118292 28024 118298 28076
rect 117869 27999 117927 28005
rect 117869 27996 117881 27999
rect 117608 27968 117881 27996
rect 117501 27959 117559 27965
rect 117869 27965 117881 27968
rect 117915 27965 117927 27999
rect 117869 27959 117927 27965
rect 116857 27931 116915 27937
rect 115032 27900 116624 27928
rect 111886 27820 111892 27872
rect 111944 27820 111950 27872
rect 112073 27863 112131 27869
rect 112073 27829 112085 27863
rect 112119 27860 112131 27863
rect 112254 27860 112260 27872
rect 112119 27832 112260 27860
rect 112119 27829 112131 27832
rect 112073 27823 112131 27829
rect 112254 27820 112260 27832
rect 112312 27820 112318 27872
rect 115014 27820 115020 27872
rect 115072 27820 115078 27872
rect 116486 27820 116492 27872
rect 116544 27820 116550 27872
rect 116596 27860 116624 27900
rect 116857 27897 116869 27931
rect 116903 27928 116915 27931
rect 117516 27928 117544 27959
rect 116903 27900 117544 27928
rect 116903 27897 116915 27900
rect 116857 27891 116915 27897
rect 116949 27863 117007 27869
rect 116949 27860 116961 27863
rect 116596 27832 116961 27860
rect 116949 27829 116961 27832
rect 116995 27829 117007 27863
rect 116949 27823 117007 27829
rect 1104 27770 7912 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 7912 27770
rect 1104 27696 7912 27718
rect 108008 27770 118864 27792
rect 108008 27718 112914 27770
rect 112966 27718 112978 27770
rect 113030 27718 113042 27770
rect 113094 27718 113106 27770
rect 113158 27718 113170 27770
rect 113222 27718 118864 27770
rect 108008 27696 118864 27718
rect 109954 27616 109960 27668
rect 110012 27656 110018 27668
rect 110325 27659 110383 27665
rect 110325 27656 110337 27659
rect 110012 27628 110337 27656
rect 110012 27616 110018 27628
rect 110325 27625 110337 27628
rect 110371 27625 110383 27659
rect 110325 27619 110383 27625
rect 110984 27628 112392 27656
rect 110046 27588 110052 27600
rect 109788 27560 110052 27588
rect 109788 27461 109816 27560
rect 110046 27548 110052 27560
rect 110104 27588 110110 27600
rect 110984 27588 111012 27628
rect 110104 27560 111012 27588
rect 110104 27548 110110 27560
rect 111058 27548 111064 27600
rect 111116 27548 111122 27600
rect 112254 27588 112260 27600
rect 111168 27560 112260 27588
rect 109862 27480 109868 27532
rect 109920 27480 109926 27532
rect 111168 27520 111196 27560
rect 112254 27548 112260 27560
rect 112312 27548 112318 27600
rect 112364 27588 112392 27628
rect 114462 27616 114468 27668
rect 114520 27616 114526 27668
rect 116118 27616 116124 27668
rect 116176 27656 116182 27668
rect 116949 27659 117007 27665
rect 116949 27656 116961 27659
rect 116176 27628 116961 27656
rect 116176 27616 116182 27628
rect 116949 27625 116961 27628
rect 116995 27656 117007 27659
rect 117038 27656 117044 27668
rect 116995 27628 117044 27656
rect 116995 27625 117007 27628
rect 116949 27619 117007 27625
rect 117038 27616 117044 27628
rect 117096 27616 117102 27668
rect 118234 27616 118240 27668
rect 118292 27616 118298 27668
rect 112364 27560 113220 27588
rect 110892 27492 111196 27520
rect 110892 27461 110920 27492
rect 111242 27480 111248 27532
rect 111300 27520 111306 27532
rect 111705 27523 111763 27529
rect 111300 27492 111472 27520
rect 111300 27480 111306 27492
rect 109773 27455 109831 27461
rect 109773 27421 109785 27455
rect 109819 27421 109831 27455
rect 110233 27455 110291 27461
rect 110233 27452 110245 27455
rect 109773 27415 109831 27421
rect 110156 27424 110245 27452
rect 110156 27384 110184 27424
rect 110233 27421 110245 27424
rect 110279 27421 110291 27455
rect 110233 27415 110291 27421
rect 110417 27455 110475 27461
rect 110417 27421 110429 27455
rect 110463 27452 110475 27455
rect 110877 27455 110935 27461
rect 110877 27452 110889 27455
rect 110463 27424 110889 27452
rect 110463 27421 110475 27424
rect 110417 27415 110475 27421
rect 110877 27421 110889 27424
rect 110923 27452 110935 27455
rect 110966 27452 110972 27464
rect 110923 27424 110972 27452
rect 110923 27421 110935 27424
rect 110877 27415 110935 27421
rect 110966 27412 110972 27424
rect 111024 27412 111030 27464
rect 111153 27455 111211 27461
rect 111153 27421 111165 27455
rect 111199 27421 111211 27455
rect 111153 27415 111211 27421
rect 110693 27387 110751 27393
rect 110693 27384 110705 27387
rect 110156 27356 110705 27384
rect 110156 27325 110184 27356
rect 110693 27353 110705 27356
rect 110739 27353 110751 27387
rect 111168 27384 111196 27415
rect 111334 27412 111340 27464
rect 111392 27412 111398 27464
rect 111444 27452 111472 27492
rect 111705 27489 111717 27523
rect 111751 27520 111763 27523
rect 111886 27520 111892 27532
rect 111751 27492 111892 27520
rect 111751 27489 111763 27492
rect 111705 27483 111763 27489
rect 111886 27480 111892 27492
rect 111944 27480 111950 27532
rect 111981 27455 112039 27461
rect 111981 27452 111993 27455
rect 111444 27424 111993 27452
rect 111981 27421 111993 27424
rect 112027 27421 112039 27455
rect 111981 27415 112039 27421
rect 112254 27412 112260 27464
rect 112312 27412 112318 27464
rect 113192 27461 113220 27560
rect 113542 27548 113548 27600
rect 113600 27588 113606 27600
rect 116489 27591 116547 27597
rect 113600 27560 114784 27588
rect 113600 27548 113606 27560
rect 113266 27480 113272 27532
rect 113324 27480 113330 27532
rect 114094 27480 114100 27532
rect 114152 27520 114158 27532
rect 114189 27523 114247 27529
rect 114189 27520 114201 27523
rect 114152 27492 114201 27520
rect 114152 27480 114158 27492
rect 114189 27489 114201 27492
rect 114235 27489 114247 27523
rect 114189 27483 114247 27489
rect 113177 27455 113235 27461
rect 113177 27421 113189 27455
rect 113223 27421 113235 27455
rect 113177 27415 113235 27421
rect 114646 27412 114652 27464
rect 114704 27412 114710 27464
rect 114756 27461 114784 27560
rect 116489 27557 116501 27591
rect 116535 27557 116547 27591
rect 116489 27551 116547 27557
rect 115290 27480 115296 27532
rect 115348 27520 115354 27532
rect 115845 27523 115903 27529
rect 115845 27520 115857 27523
rect 115348 27492 115857 27520
rect 115348 27480 115354 27492
rect 115845 27489 115857 27492
rect 115891 27489 115903 27523
rect 115845 27483 115903 27489
rect 114741 27455 114799 27461
rect 114741 27421 114753 27455
rect 114787 27421 114799 27455
rect 114741 27415 114799 27421
rect 114922 27412 114928 27464
rect 114980 27412 114986 27464
rect 115014 27412 115020 27464
rect 115072 27412 115078 27464
rect 115477 27455 115535 27461
rect 115477 27421 115489 27455
rect 115523 27421 115535 27455
rect 115477 27415 115535 27421
rect 111797 27387 111855 27393
rect 111797 27384 111809 27387
rect 111168 27356 111809 27384
rect 110693 27347 110751 27353
rect 111797 27353 111809 27356
rect 111843 27353 111855 27387
rect 111797 27347 111855 27353
rect 112530 27344 112536 27396
rect 112588 27344 112594 27396
rect 112714 27344 112720 27396
rect 112772 27384 112778 27396
rect 114005 27387 114063 27393
rect 112772 27356 113680 27384
rect 112772 27344 112778 27356
rect 110141 27319 110199 27325
rect 110141 27285 110153 27319
rect 110187 27285 110199 27319
rect 110141 27279 110199 27285
rect 111613 27319 111671 27325
rect 111613 27285 111625 27319
rect 111659 27316 111671 27319
rect 111978 27316 111984 27328
rect 111659 27288 111984 27316
rect 111659 27285 111671 27288
rect 111613 27279 111671 27285
rect 111978 27276 111984 27288
rect 112036 27276 112042 27328
rect 112162 27276 112168 27328
rect 112220 27316 112226 27328
rect 113652 27325 113680 27356
rect 114005 27353 114017 27387
rect 114051 27384 114063 27387
rect 115382 27384 115388 27396
rect 114051 27356 115388 27384
rect 114051 27353 114063 27356
rect 114005 27347 114063 27353
rect 115382 27344 115388 27356
rect 115440 27344 115446 27396
rect 115492 27384 115520 27415
rect 115934 27412 115940 27464
rect 115992 27452 115998 27464
rect 116029 27455 116087 27461
rect 116029 27452 116041 27455
rect 115992 27424 116041 27452
rect 115992 27412 115998 27424
rect 116029 27421 116041 27424
rect 116075 27421 116087 27455
rect 116029 27415 116087 27421
rect 116118 27412 116124 27464
rect 116176 27452 116182 27464
rect 116305 27455 116363 27461
rect 116305 27452 116317 27455
rect 116176 27424 116317 27452
rect 116176 27412 116182 27424
rect 116305 27421 116317 27424
rect 116351 27452 116363 27455
rect 116504 27452 116532 27551
rect 117406 27548 117412 27600
rect 117464 27588 117470 27600
rect 117501 27591 117559 27597
rect 117501 27588 117513 27591
rect 117464 27560 117513 27588
rect 117464 27548 117470 27560
rect 117501 27557 117513 27560
rect 117547 27557 117559 27591
rect 117501 27551 117559 27557
rect 118326 27548 118332 27600
rect 118384 27548 118390 27600
rect 116762 27480 116768 27532
rect 116820 27480 116826 27532
rect 117590 27480 117596 27532
rect 117648 27520 117654 27532
rect 117777 27523 117835 27529
rect 117777 27520 117789 27523
rect 117648 27492 117789 27520
rect 117648 27480 117654 27492
rect 117777 27489 117789 27492
rect 117823 27489 117835 27523
rect 117777 27483 117835 27489
rect 116351 27424 116532 27452
rect 116351 27421 116363 27424
rect 116305 27415 116363 27421
rect 116578 27412 116584 27464
rect 116636 27452 116642 27464
rect 116673 27455 116731 27461
rect 116673 27452 116685 27455
rect 116636 27424 116685 27452
rect 116636 27412 116642 27424
rect 116673 27421 116685 27424
rect 116719 27421 116731 27455
rect 116673 27415 116731 27421
rect 116854 27412 116860 27464
rect 116912 27452 116918 27464
rect 116949 27455 117007 27461
rect 116949 27452 116961 27455
rect 116912 27424 116961 27452
rect 116912 27412 116918 27424
rect 116949 27421 116961 27424
rect 116995 27421 117007 27455
rect 116949 27415 117007 27421
rect 117869 27455 117927 27461
rect 117869 27421 117881 27455
rect 117915 27452 117927 27455
rect 118142 27452 118148 27464
rect 117915 27424 118148 27452
rect 117915 27421 117927 27424
rect 117869 27415 117927 27421
rect 118142 27412 118148 27424
rect 118200 27412 118206 27464
rect 118510 27412 118516 27464
rect 118568 27412 118574 27464
rect 116213 27387 116271 27393
rect 116213 27384 116225 27387
rect 115492 27356 116225 27384
rect 116213 27353 116225 27356
rect 116259 27384 116271 27387
rect 116486 27384 116492 27396
rect 116259 27356 116492 27384
rect 116259 27353 116271 27356
rect 116213 27347 116271 27353
rect 116486 27344 116492 27356
rect 116544 27344 116550 27396
rect 112349 27319 112407 27325
rect 112349 27316 112361 27319
rect 112220 27288 112361 27316
rect 112220 27276 112226 27288
rect 112349 27285 112361 27288
rect 112395 27285 112407 27319
rect 112349 27279 112407 27285
rect 113637 27319 113695 27325
rect 113637 27285 113649 27319
rect 113683 27285 113695 27319
rect 113637 27279 113695 27285
rect 114094 27276 114100 27328
rect 114152 27276 114158 27328
rect 115658 27276 115664 27328
rect 115716 27276 115722 27328
rect 1104 27226 7912 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 7912 27226
rect 1104 27152 7912 27174
rect 108008 27226 118864 27248
rect 108008 27174 113650 27226
rect 113702 27174 113714 27226
rect 113766 27174 113778 27226
rect 113830 27174 113842 27226
rect 113894 27174 113906 27226
rect 113958 27174 118864 27226
rect 108008 27152 118864 27174
rect 110782 27072 110788 27124
rect 110840 27072 110846 27124
rect 113913 27115 113971 27121
rect 113913 27081 113925 27115
rect 113959 27112 113971 27115
rect 114002 27112 114008 27124
rect 113959 27084 114008 27112
rect 113959 27081 113971 27084
rect 113913 27075 113971 27081
rect 114002 27072 114008 27084
rect 114060 27072 114066 27124
rect 114830 27072 114836 27124
rect 114888 27072 114894 27124
rect 115290 27072 115296 27124
rect 115348 27072 115354 27124
rect 115382 27072 115388 27124
rect 115440 27072 115446 27124
rect 118510 27072 118516 27124
rect 118568 27072 118574 27124
rect 112162 27044 112168 27056
rect 111076 27016 112168 27044
rect 110966 26936 110972 26988
rect 111024 26936 111030 26988
rect 111076 26985 111104 27016
rect 112162 27004 112168 27016
rect 112220 27004 112226 27056
rect 112530 27004 112536 27056
rect 112588 27044 112594 27056
rect 114848 27044 114876 27072
rect 115937 27047 115995 27053
rect 115937 27044 115949 27047
rect 112588 27016 114876 27044
rect 115676 27016 115949 27044
rect 112588 27004 112594 27016
rect 115676 26988 115704 27016
rect 115937 27013 115949 27016
rect 115983 27013 115995 27047
rect 115937 27007 115995 27013
rect 116118 27004 116124 27056
rect 116176 27004 116182 27056
rect 111061 26979 111119 26985
rect 111061 26945 111073 26979
rect 111107 26945 111119 26979
rect 111061 26939 111119 26945
rect 111242 26936 111248 26988
rect 111300 26936 111306 26988
rect 111334 26936 111340 26988
rect 111392 26976 111398 26988
rect 111392 26948 111748 26976
rect 111392 26936 111398 26948
rect 111720 26849 111748 26948
rect 112070 26936 112076 26988
rect 112128 26936 112134 26988
rect 113542 26936 113548 26988
rect 113600 26936 113606 26988
rect 114738 26936 114744 26988
rect 114796 26976 114802 26988
rect 114833 26979 114891 26985
rect 114833 26976 114845 26979
rect 114796 26948 114845 26976
rect 114796 26936 114802 26948
rect 114833 26945 114845 26948
rect 114879 26945 114891 26979
rect 114833 26939 114891 26945
rect 115569 26979 115627 26985
rect 115569 26945 115581 26979
rect 115615 26945 115627 26979
rect 115569 26939 115627 26945
rect 112165 26911 112223 26917
rect 112165 26877 112177 26911
rect 112211 26908 112223 26911
rect 112346 26908 112352 26920
rect 112211 26880 112352 26908
rect 112211 26877 112223 26880
rect 112165 26871 112223 26877
rect 112346 26868 112352 26880
rect 112404 26868 112410 26920
rect 113637 26911 113695 26917
rect 113637 26877 113649 26911
rect 113683 26908 113695 26911
rect 114646 26908 114652 26920
rect 113683 26880 114652 26908
rect 113683 26877 113695 26880
rect 113637 26871 113695 26877
rect 114646 26868 114652 26880
rect 114704 26868 114710 26920
rect 114925 26911 114983 26917
rect 114925 26877 114937 26911
rect 114971 26877 114983 26911
rect 115584 26908 115612 26939
rect 115658 26936 115664 26988
rect 115716 26936 115722 26988
rect 115842 26936 115848 26988
rect 115900 26936 115906 26988
rect 116136 26908 116164 27004
rect 115584 26880 116164 26908
rect 114925 26871 114983 26877
rect 111705 26843 111763 26849
rect 111705 26809 111717 26843
rect 111751 26809 111763 26843
rect 114940 26840 114968 26871
rect 114940 26812 115888 26840
rect 111705 26803 111763 26809
rect 115860 26784 115888 26812
rect 115842 26732 115848 26784
rect 115900 26732 115906 26784
rect 1104 26682 7912 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 7912 26682
rect 1104 26608 7912 26630
rect 108008 26682 118864 26704
rect 108008 26630 112914 26682
rect 112966 26630 112978 26682
rect 113030 26630 113042 26682
rect 113094 26630 113106 26682
rect 113158 26630 113170 26682
rect 113222 26630 118864 26682
rect 108008 26608 118864 26630
rect 111242 26528 111248 26580
rect 111300 26568 111306 26580
rect 111429 26571 111487 26577
rect 111429 26568 111441 26571
rect 111300 26540 111441 26568
rect 111300 26528 111306 26540
rect 111429 26537 111441 26540
rect 111475 26537 111487 26571
rect 111429 26531 111487 26537
rect 114094 26528 114100 26580
rect 114152 26568 114158 26580
rect 114649 26571 114707 26577
rect 114649 26568 114661 26571
rect 114152 26540 114661 26568
rect 114152 26528 114158 26540
rect 114649 26537 114661 26540
rect 114695 26537 114707 26571
rect 114649 26531 114707 26537
rect 115290 26528 115296 26580
rect 115348 26568 115354 26580
rect 115842 26568 115848 26580
rect 115348 26540 115848 26568
rect 115348 26528 115354 26540
rect 115842 26528 115848 26540
rect 115900 26528 115906 26580
rect 115109 26503 115167 26509
rect 115109 26469 115121 26503
rect 115155 26469 115167 26503
rect 115109 26463 115167 26469
rect 112714 26432 112720 26444
rect 111628 26404 112720 26432
rect 109862 26324 109868 26376
rect 109920 26364 109926 26376
rect 111628 26373 111656 26404
rect 112714 26392 112720 26404
rect 112772 26392 112778 26444
rect 111613 26367 111671 26373
rect 111613 26364 111625 26367
rect 109920 26336 111625 26364
rect 109920 26324 109926 26336
rect 111613 26333 111625 26336
rect 111659 26333 111671 26367
rect 111613 26327 111671 26333
rect 111797 26367 111855 26373
rect 111797 26333 111809 26367
rect 111843 26364 111855 26367
rect 112530 26364 112536 26376
rect 111843 26336 112536 26364
rect 111843 26333 111855 26336
rect 111797 26327 111855 26333
rect 112530 26324 112536 26336
rect 112588 26324 112594 26376
rect 114833 26367 114891 26373
rect 114833 26333 114845 26367
rect 114879 26364 114891 26367
rect 115124 26364 115152 26463
rect 114879 26336 115152 26364
rect 114879 26333 114891 26336
rect 114833 26327 114891 26333
rect 115014 26256 115020 26308
rect 115072 26256 115078 26308
rect 115382 26256 115388 26308
rect 115440 26296 115446 26308
rect 115477 26299 115535 26305
rect 115477 26296 115489 26299
rect 115440 26268 115489 26296
rect 115440 26256 115446 26268
rect 115477 26265 115489 26268
rect 115523 26265 115535 26299
rect 115477 26259 115535 26265
rect 114738 26188 114744 26240
rect 114796 26228 114802 26240
rect 115267 26231 115325 26237
rect 115267 26228 115279 26231
rect 114796 26200 115279 26228
rect 114796 26188 114802 26200
rect 115267 26197 115279 26200
rect 115313 26197 115325 26231
rect 115267 26191 115325 26197
rect 1104 26138 7912 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 7912 26138
rect 1104 26064 7912 26086
rect 108008 26138 118864 26160
rect 108008 26086 113650 26138
rect 113702 26086 113714 26138
rect 113766 26086 113778 26138
rect 113830 26086 113842 26138
rect 113894 26086 113906 26138
rect 113958 26086 118864 26138
rect 108008 26064 118864 26086
rect 115017 26027 115075 26033
rect 115017 25993 115029 26027
rect 115063 26024 115075 26027
rect 115382 26024 115388 26036
rect 115063 25996 115388 26024
rect 115063 25993 115075 25996
rect 115017 25987 115075 25993
rect 115382 25984 115388 25996
rect 115440 25984 115446 26036
rect 114738 25916 114744 25968
rect 114796 25956 114802 25968
rect 114833 25959 114891 25965
rect 114833 25956 114845 25959
rect 114796 25928 114845 25956
rect 114796 25916 114802 25928
rect 114833 25925 114845 25928
rect 114879 25925 114891 25959
rect 114833 25919 114891 25925
rect 115109 25891 115167 25897
rect 115109 25857 115121 25891
rect 115155 25888 115167 25891
rect 115290 25888 115296 25900
rect 115155 25860 115296 25888
rect 115155 25857 115167 25860
rect 115109 25851 115167 25857
rect 115290 25848 115296 25860
rect 115348 25848 115354 25900
rect 114833 25755 114891 25761
rect 114833 25721 114845 25755
rect 114879 25752 114891 25755
rect 115014 25752 115020 25764
rect 114879 25724 115020 25752
rect 114879 25721 114891 25724
rect 114833 25715 114891 25721
rect 115014 25712 115020 25724
rect 115072 25712 115078 25764
rect 1104 25594 7912 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 7912 25594
rect 1104 25520 7912 25542
rect 108008 25594 118864 25616
rect 108008 25542 112914 25594
rect 112966 25542 112978 25594
rect 113030 25542 113042 25594
rect 113094 25542 113106 25594
rect 113158 25542 113170 25594
rect 113222 25542 118864 25594
rect 108008 25520 118864 25542
rect 1104 25050 7912 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 7912 25050
rect 1104 24976 7912 24998
rect 108008 25050 118864 25072
rect 108008 24998 113650 25050
rect 113702 24998 113714 25050
rect 113766 24998 113778 25050
rect 113830 24998 113842 25050
rect 113894 24998 113906 25050
rect 113958 24998 118864 25050
rect 108008 24976 118864 24998
rect 1104 24506 7912 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 7912 24506
rect 1104 24432 7912 24454
rect 108008 24506 118864 24528
rect 108008 24454 112914 24506
rect 112966 24454 112978 24506
rect 113030 24454 113042 24506
rect 113094 24454 113106 24506
rect 113158 24454 113170 24506
rect 113222 24454 118864 24506
rect 108008 24432 118864 24454
rect 1104 23962 7912 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 7912 23962
rect 1104 23888 7912 23910
rect 108008 23962 118864 23984
rect 108008 23910 113650 23962
rect 113702 23910 113714 23962
rect 113766 23910 113778 23962
rect 113830 23910 113842 23962
rect 113894 23910 113906 23962
rect 113958 23910 118864 23962
rect 108008 23888 118864 23910
rect 1104 23418 7912 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 7912 23418
rect 1104 23344 7912 23366
rect 108008 23418 118864 23440
rect 108008 23366 112914 23418
rect 112966 23366 112978 23418
rect 113030 23366 113042 23418
rect 113094 23366 113106 23418
rect 113158 23366 113170 23418
rect 113222 23366 118864 23418
rect 108008 23344 118864 23366
rect 1104 22874 7912 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 7912 22874
rect 1104 22800 7912 22822
rect 108008 22874 118864 22896
rect 108008 22822 113650 22874
rect 113702 22822 113714 22874
rect 113766 22822 113778 22874
rect 113830 22822 113842 22874
rect 113894 22822 113906 22874
rect 113958 22822 118864 22874
rect 108008 22800 118864 22822
rect 1104 22330 7912 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 7912 22330
rect 1104 22256 7912 22278
rect 108008 22330 118864 22352
rect 108008 22278 112914 22330
rect 112966 22278 112978 22330
rect 113030 22278 113042 22330
rect 113094 22278 113106 22330
rect 113158 22278 113170 22330
rect 113222 22278 118864 22330
rect 108008 22256 118864 22278
rect 1104 21786 7912 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 7912 21786
rect 1104 21712 7912 21734
rect 108008 21786 118864 21808
rect 108008 21734 113650 21786
rect 113702 21734 113714 21786
rect 113766 21734 113778 21786
rect 113830 21734 113842 21786
rect 113894 21734 113906 21786
rect 113958 21734 118864 21786
rect 108008 21712 118864 21734
rect 1104 21242 7912 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 7912 21242
rect 1104 21168 7912 21190
rect 108008 21242 118864 21264
rect 108008 21190 112914 21242
rect 112966 21190 112978 21242
rect 113030 21190 113042 21242
rect 113094 21190 113106 21242
rect 113158 21190 113170 21242
rect 113222 21190 118864 21242
rect 108008 21168 118864 21190
rect 1104 20698 7912 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 7912 20698
rect 1104 20624 7912 20646
rect 108008 20698 118864 20720
rect 108008 20646 113650 20698
rect 113702 20646 113714 20698
rect 113766 20646 113778 20698
rect 113830 20646 113842 20698
rect 113894 20646 113906 20698
rect 113958 20646 118864 20698
rect 108008 20624 118864 20646
rect 1104 20154 7912 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 7912 20154
rect 1104 20080 7912 20102
rect 108008 20154 118864 20176
rect 108008 20102 112914 20154
rect 112966 20102 112978 20154
rect 113030 20102 113042 20154
rect 113094 20102 113106 20154
rect 113158 20102 113170 20154
rect 113222 20102 118864 20154
rect 108008 20080 118864 20102
rect 1104 19610 7912 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 7912 19610
rect 1104 19536 7912 19558
rect 108008 19610 118864 19632
rect 108008 19558 113650 19610
rect 113702 19558 113714 19610
rect 113766 19558 113778 19610
rect 113830 19558 113842 19610
rect 113894 19558 113906 19610
rect 113958 19558 118864 19610
rect 108008 19536 118864 19558
rect 1104 19066 7912 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 7912 19066
rect 1104 18992 7912 19014
rect 108008 19066 118864 19088
rect 108008 19014 112914 19066
rect 112966 19014 112978 19066
rect 113030 19014 113042 19066
rect 113094 19014 113106 19066
rect 113158 19014 113170 19066
rect 113222 19014 118864 19066
rect 108008 18992 118864 19014
rect 1104 18522 7912 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 7912 18522
rect 1104 18448 7912 18470
rect 108008 18522 118864 18544
rect 108008 18470 113650 18522
rect 113702 18470 113714 18522
rect 113766 18470 113778 18522
rect 113830 18470 113842 18522
rect 113894 18470 113906 18522
rect 113958 18470 118864 18522
rect 108008 18448 118864 18470
rect 1104 17978 7912 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 7912 17978
rect 1104 17904 7912 17926
rect 108008 17978 118864 18000
rect 108008 17926 112914 17978
rect 112966 17926 112978 17978
rect 113030 17926 113042 17978
rect 113094 17926 113106 17978
rect 113158 17926 113170 17978
rect 113222 17926 118864 17978
rect 108008 17904 118864 17926
rect 7561 17663 7619 17669
rect 7561 17629 7573 17663
rect 7607 17660 7619 17663
rect 9674 17660 9680 17672
rect 7607 17632 9680 17660
rect 7607 17629 7619 17632
rect 7561 17623 7619 17629
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 1104 17434 7912 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 7912 17434
rect 1104 17360 7912 17382
rect 108008 17434 118864 17456
rect 108008 17382 113650 17434
rect 113702 17382 113714 17434
rect 113766 17382 113778 17434
rect 113830 17382 113842 17434
rect 113894 17382 113906 17434
rect 113958 17382 118864 17434
rect 108008 17360 118864 17382
rect 1104 16890 7912 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 7912 16890
rect 1104 16816 7912 16838
rect 108008 16890 118864 16912
rect 108008 16838 112914 16890
rect 112966 16838 112978 16890
rect 113030 16838 113042 16890
rect 113094 16838 113106 16890
rect 113158 16838 113170 16890
rect 113222 16838 118864 16890
rect 108008 16816 118864 16838
rect 1104 16346 7912 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 7912 16346
rect 1104 16272 7912 16294
rect 108008 16346 118864 16368
rect 108008 16294 113650 16346
rect 113702 16294 113714 16346
rect 113766 16294 113778 16346
rect 113830 16294 113842 16346
rect 113894 16294 113906 16346
rect 113958 16294 118864 16346
rect 108008 16272 118864 16294
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 1360 16068 1409 16096
rect 1360 16056 1366 16068
rect 1397 16065 1409 16068
rect 1443 16096 1455 16099
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1443 16068 1685 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 9674 15960 9680 15972
rect 1627 15932 9680 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 1104 15802 7912 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 7912 15802
rect 1104 15728 7912 15750
rect 108008 15802 118864 15824
rect 108008 15750 112914 15802
rect 112966 15750 112978 15802
rect 113030 15750 113042 15802
rect 113094 15750 113106 15802
rect 113158 15750 113170 15802
rect 113222 15750 118864 15802
rect 108008 15728 118864 15750
rect 1104 15258 7912 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 7912 15258
rect 1104 15184 7912 15206
rect 108008 15258 118864 15280
rect 108008 15206 113650 15258
rect 113702 15206 113714 15258
rect 113766 15206 113778 15258
rect 113830 15206 113842 15258
rect 113894 15206 113906 15258
rect 113958 15206 118864 15258
rect 108008 15184 118864 15206
rect 1104 14714 7912 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 7912 14714
rect 1104 14640 7912 14662
rect 108008 14714 118864 14736
rect 108008 14662 112914 14714
rect 112966 14662 112978 14714
rect 113030 14662 113042 14714
rect 113094 14662 113106 14714
rect 113158 14662 113170 14714
rect 113222 14662 118864 14714
rect 108008 14640 118864 14662
rect 1104 14170 7912 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 7912 14170
rect 1104 14096 7912 14118
rect 108008 14170 118864 14192
rect 108008 14118 113650 14170
rect 113702 14118 113714 14170
rect 113766 14118 113778 14170
rect 113830 14118 113842 14170
rect 113894 14118 113906 14170
rect 113958 14118 118864 14170
rect 108008 14096 118864 14118
rect 1104 13626 7912 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 7912 13626
rect 1104 13552 7912 13574
rect 108008 13626 118864 13648
rect 108008 13574 112914 13626
rect 112966 13574 112978 13626
rect 113030 13574 113042 13626
rect 113094 13574 113106 13626
rect 113158 13574 113170 13626
rect 113222 13574 118864 13626
rect 108008 13552 118864 13574
rect 1104 13082 7912 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 7912 13082
rect 1104 13008 7912 13030
rect 108008 13082 118864 13104
rect 108008 13030 113650 13082
rect 113702 13030 113714 13082
rect 113766 13030 113778 13082
rect 113830 13030 113842 13082
rect 113894 13030 113906 13082
rect 113958 13030 118864 13082
rect 108008 13008 118864 13030
rect 1104 12538 7912 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 7912 12538
rect 1104 12464 7912 12486
rect 108008 12538 118864 12560
rect 108008 12486 112914 12538
rect 112966 12486 112978 12538
rect 113030 12486 113042 12538
rect 113094 12486 113106 12538
rect 113158 12486 113170 12538
rect 113222 12486 118864 12538
rect 108008 12464 118864 12486
rect 1104 11994 7912 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 7912 11994
rect 1104 11920 7912 11942
rect 108008 11994 118864 12016
rect 108008 11942 113650 11994
rect 113702 11942 113714 11994
rect 113766 11942 113778 11994
rect 113830 11942 113842 11994
rect 113894 11942 113906 11994
rect 113958 11942 118864 11994
rect 108008 11920 118864 11942
rect 1104 11450 7912 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 7912 11450
rect 1104 11376 7912 11398
rect 108008 11450 118864 11472
rect 108008 11398 112914 11450
rect 112966 11398 112978 11450
rect 113030 11398 113042 11450
rect 113094 11398 113106 11450
rect 113158 11398 113170 11450
rect 113222 11398 118864 11450
rect 108008 11376 118864 11398
rect 1104 10906 7912 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 7912 10906
rect 1104 10832 7912 10854
rect 108008 10906 118864 10928
rect 108008 10854 113650 10906
rect 113702 10854 113714 10906
rect 113766 10854 113778 10906
rect 113830 10854 113842 10906
rect 113894 10854 113906 10906
rect 113958 10854 118864 10906
rect 108008 10832 118864 10854
rect 1104 10362 7912 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 7912 10362
rect 1104 10288 7912 10310
rect 108008 10362 118864 10384
rect 108008 10310 112914 10362
rect 112966 10310 112978 10362
rect 113030 10310 113042 10362
rect 113094 10310 113106 10362
rect 113158 10310 113170 10362
rect 113222 10310 118864 10362
rect 108008 10288 118864 10310
rect 93394 10004 93400 10056
rect 93452 10044 93458 10056
rect 109494 10044 109500 10056
rect 93452 10016 109500 10044
rect 93452 10004 93458 10016
rect 109494 10004 109500 10016
rect 109552 10004 109558 10056
rect 92842 9936 92848 9988
rect 92900 9976 92906 9988
rect 108298 9976 108304 9988
rect 92900 9948 108304 9976
rect 92900 9936 92906 9948
rect 108298 9936 108304 9948
rect 108356 9936 108362 9988
rect 93026 9868 93032 9920
rect 93084 9908 93090 9920
rect 106458 9908 106464 9920
rect 93084 9880 106464 9908
rect 93084 9868 93090 9880
rect 106458 9868 106464 9880
rect 106516 9868 106522 9920
rect 1104 9818 7912 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 7912 9818
rect 1104 9744 7912 9766
rect 108008 9818 118864 9840
rect 108008 9766 113650 9818
rect 113702 9766 113714 9818
rect 113766 9766 113778 9818
rect 113830 9766 113842 9818
rect 113894 9766 113906 9818
rect 113958 9766 118864 9818
rect 108008 9744 118864 9766
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 15838 9636 15844 9648
rect 8260 9608 15844 9636
rect 8260 9596 8266 9608
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 1104 9274 7912 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 7912 9274
rect 1104 9200 7912 9222
rect 108008 9274 118864 9296
rect 108008 9222 112914 9274
rect 112966 9222 112978 9274
rect 113030 9222 113042 9274
rect 113094 9222 113106 9274
rect 113158 9222 113170 9274
rect 113222 9222 118864 9274
rect 108008 9200 118864 9222
rect 1104 8730 7912 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 7912 8730
rect 1104 8656 7912 8678
rect 108008 8730 118864 8752
rect 108008 8678 113650 8730
rect 113702 8678 113714 8730
rect 113766 8678 113778 8730
rect 113830 8678 113842 8730
rect 113894 8678 113906 8730
rect 113958 8678 118864 8730
rect 108008 8656 118864 8678
rect 1104 8186 7912 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 7912 8186
rect 1104 8112 7912 8134
rect 108008 8186 118864 8208
rect 108008 8134 112914 8186
rect 112966 8134 112978 8186
rect 113030 8134 113042 8186
rect 113094 8134 113106 8186
rect 113158 8134 113170 8186
rect 113222 8134 118864 8186
rect 108008 8112 118864 8134
rect 1104 7642 118864 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 66314 7642
rect 66366 7590 66378 7642
rect 66430 7590 66442 7642
rect 66494 7590 66506 7642
rect 66558 7590 66570 7642
rect 66622 7590 97034 7642
rect 97086 7590 97098 7642
rect 97150 7590 97162 7642
rect 97214 7590 97226 7642
rect 97278 7590 97290 7642
rect 97342 7590 113650 7642
rect 113702 7590 113714 7642
rect 113766 7590 113778 7642
rect 113830 7590 113842 7642
rect 113894 7590 113906 7642
rect 113958 7590 118864 7642
rect 1104 7568 118864 7590
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 15933 7531 15991 7537
rect 15933 7528 15945 7531
rect 15896 7500 15945 7528
rect 15896 7488 15902 7500
rect 15933 7497 15945 7500
rect 15979 7497 15991 7531
rect 15933 7491 15991 7497
rect 26970 7488 26976 7540
rect 27028 7488 27034 7540
rect 27798 7488 27804 7540
rect 27856 7528 27862 7540
rect 27893 7531 27951 7537
rect 27893 7528 27905 7531
rect 27856 7500 27905 7528
rect 27856 7488 27862 7500
rect 27893 7497 27905 7500
rect 27939 7497 27951 7531
rect 27893 7491 27951 7497
rect 29546 7488 29552 7540
rect 29604 7488 29610 7540
rect 30190 7488 30196 7540
rect 30248 7488 30254 7540
rect 92842 7488 92848 7540
rect 92900 7488 92906 7540
rect 93026 7488 93032 7540
rect 93084 7488 93090 7540
rect 93210 7488 93216 7540
rect 93268 7488 93274 7540
rect 93394 7488 93400 7540
rect 93452 7488 93458 7540
rect 1104 7098 118864 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 112914 7098
rect 112966 7046 112978 7098
rect 113030 7046 113042 7098
rect 113094 7046 113106 7098
rect 113158 7046 113170 7098
rect 113222 7046 118864 7098
rect 1104 7024 118864 7046
rect 1104 6554 118864 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 66314 6554
rect 66366 6502 66378 6554
rect 66430 6502 66442 6554
rect 66494 6502 66506 6554
rect 66558 6502 66570 6554
rect 66622 6502 97034 6554
rect 97086 6502 97098 6554
rect 97150 6502 97162 6554
rect 97214 6502 97226 6554
rect 97278 6502 97290 6554
rect 97342 6502 118864 6554
rect 1104 6480 118864 6502
rect 1104 6010 118864 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 118864 6010
rect 1104 5936 118864 5958
rect 1104 5466 118864 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 66314 5466
rect 66366 5414 66378 5466
rect 66430 5414 66442 5466
rect 66494 5414 66506 5466
rect 66558 5414 66570 5466
rect 66622 5414 97034 5466
rect 97086 5414 97098 5466
rect 97150 5414 97162 5466
rect 97214 5414 97226 5466
rect 97278 5414 97290 5466
rect 97342 5414 118864 5466
rect 1104 5392 118864 5414
rect 1104 4922 118864 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 118864 4922
rect 1104 4848 118864 4870
rect 1104 4378 118864 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 66314 4378
rect 66366 4326 66378 4378
rect 66430 4326 66442 4378
rect 66494 4326 66506 4378
rect 66558 4326 66570 4378
rect 66622 4326 97034 4378
rect 97086 4326 97098 4378
rect 97150 4326 97162 4378
rect 97214 4326 97226 4378
rect 97278 4326 97290 4378
rect 97342 4326 118864 4378
rect 1104 4304 118864 4326
rect 1104 3834 118864 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 118864 3834
rect 1104 3760 118864 3782
rect 1104 3290 118864 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 66314 3290
rect 66366 3238 66378 3290
rect 66430 3238 66442 3290
rect 66494 3238 66506 3290
rect 66558 3238 66570 3290
rect 66622 3238 97034 3290
rect 97086 3238 97098 3290
rect 97150 3238 97162 3290
rect 97214 3238 97226 3290
rect 97278 3238 97290 3290
rect 97342 3238 118864 3290
rect 1104 3216 118864 3238
rect 1104 2746 118864 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 118864 2746
rect 1104 2672 118864 2694
rect 25866 2592 25872 2644
rect 25924 2592 25930 2644
rect 31662 2592 31668 2644
rect 31720 2592 31726 2644
rect 32950 2592 32956 2644
rect 33008 2592 33014 2644
rect 33778 2592 33784 2644
rect 33836 2592 33842 2644
rect 34790 2592 34796 2644
rect 34848 2632 34854 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 34848 2604 35081 2632
rect 34848 2592 34854 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 36170 2592 36176 2644
rect 36228 2592 36234 2644
rect 37458 2592 37464 2644
rect 37516 2592 37522 2644
rect 38286 2592 38292 2644
rect 38344 2592 38350 2644
rect 40034 2592 40040 2644
rect 40092 2592 40098 2644
rect 40862 2592 40868 2644
rect 40920 2592 40926 2644
rect 41966 2592 41972 2644
rect 42024 2592 42030 2644
rect 43254 2592 43260 2644
rect 43312 2592 43318 2644
rect 44542 2592 44548 2644
rect 44600 2592 44606 2644
rect 45830 2592 45836 2644
rect 45888 2592 45894 2644
rect 46658 2592 46664 2644
rect 46716 2592 46722 2644
rect 47762 2592 47768 2644
rect 47820 2592 47826 2644
rect 49050 2592 49056 2644
rect 49108 2592 49114 2644
rect 50338 2592 50344 2644
rect 50396 2592 50402 2644
rect 51626 2592 51632 2644
rect 51684 2592 51690 2644
rect 52454 2592 52460 2644
rect 52512 2592 52518 2644
rect 53558 2592 53564 2644
rect 53616 2592 53622 2644
rect 55030 2592 55036 2644
rect 55088 2592 55094 2644
rect 56134 2592 56140 2644
rect 56192 2592 56198 2644
rect 57422 2592 57428 2644
rect 57480 2592 57486 2644
rect 58250 2592 58256 2644
rect 58308 2592 58314 2644
rect 59538 2592 59544 2644
rect 59596 2592 59602 2644
rect 60826 2592 60832 2644
rect 60884 2592 60890 2644
rect 61930 2592 61936 2644
rect 61988 2592 61994 2644
rect 63218 2592 63224 2644
rect 63276 2592 63282 2644
rect 64046 2592 64052 2644
rect 64104 2592 64110 2644
rect 65334 2592 65340 2644
rect 65392 2592 65398 2644
rect 66625 2635 66683 2641
rect 66625 2601 66637 2635
rect 66671 2632 66683 2635
rect 66714 2632 66720 2644
rect 66671 2604 66720 2632
rect 66671 2601 66683 2604
rect 66625 2595 66683 2601
rect 66714 2592 66720 2604
rect 66772 2592 66778 2644
rect 67726 2592 67732 2644
rect 67784 2592 67790 2644
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25792 2400 26065 2428
rect 25792 2304 25820 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 31849 2431 31907 2437
rect 31849 2428 31861 2431
rect 26053 2391 26111 2397
rect 31588 2400 31861 2428
rect 31588 2304 31616 2400
rect 31849 2397 31861 2400
rect 31895 2397 31907 2431
rect 33137 2431 33195 2437
rect 33137 2428 33149 2431
rect 31849 2391 31907 2397
rect 32876 2400 33149 2428
rect 32876 2304 32904 2400
rect 33137 2397 33149 2400
rect 33183 2397 33195 2431
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33137 2391 33195 2397
rect 33520 2400 33609 2428
rect 33520 2304 33548 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 33597 2391 33655 2397
rect 34808 2400 34897 2428
rect 34808 2304 34836 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 34885 2391 34943 2397
rect 36096 2400 36369 2428
rect 36096 2304 36124 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 37645 2431 37703 2437
rect 37645 2428 37657 2431
rect 36357 2391 36415 2397
rect 37384 2400 37657 2428
rect 37384 2304 37412 2400
rect 37645 2397 37657 2400
rect 37691 2397 37703 2431
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 37645 2391 37703 2397
rect 38028 2400 38117 2428
rect 38028 2304 38056 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 38105 2391 38163 2397
rect 39960 2400 40233 2428
rect 39960 2304 39988 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 40221 2391 40279 2397
rect 40604 2400 40693 2428
rect 40604 2304 40632 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 42153 2431 42211 2437
rect 42153 2428 42165 2431
rect 40681 2391 40739 2397
rect 41892 2400 42165 2428
rect 41892 2304 41920 2400
rect 42153 2397 42165 2400
rect 42199 2397 42211 2431
rect 43441 2431 43499 2437
rect 43441 2428 43453 2431
rect 42153 2391 42211 2397
rect 43180 2400 43453 2428
rect 43180 2304 43208 2400
rect 43441 2397 43453 2400
rect 43487 2397 43499 2431
rect 44729 2431 44787 2437
rect 44729 2428 44741 2431
rect 43441 2391 43499 2397
rect 44468 2400 44741 2428
rect 44468 2304 44496 2400
rect 44729 2397 44741 2400
rect 44775 2397 44787 2431
rect 46017 2431 46075 2437
rect 46017 2428 46029 2431
rect 44729 2391 44787 2397
rect 45756 2400 46029 2428
rect 45756 2304 45784 2400
rect 46017 2397 46029 2400
rect 46063 2397 46075 2431
rect 46477 2431 46535 2437
rect 46477 2428 46489 2431
rect 46017 2391 46075 2397
rect 46400 2400 46489 2428
rect 46400 2304 46428 2400
rect 46477 2397 46489 2400
rect 46523 2397 46535 2431
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 46477 2391 46535 2397
rect 47688 2400 47961 2428
rect 47688 2304 47716 2400
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 49237 2431 49295 2437
rect 49237 2428 49249 2431
rect 47949 2391 48007 2397
rect 48976 2400 49249 2428
rect 48976 2304 49004 2400
rect 49237 2397 49249 2400
rect 49283 2397 49295 2431
rect 50525 2431 50583 2437
rect 50525 2428 50537 2431
rect 49237 2391 49295 2397
rect 50264 2400 50537 2428
rect 50264 2304 50292 2400
rect 50525 2397 50537 2400
rect 50571 2397 50583 2431
rect 51813 2431 51871 2437
rect 51813 2428 51825 2431
rect 50525 2391 50583 2397
rect 51552 2400 51825 2428
rect 51552 2304 51580 2400
rect 51813 2397 51825 2400
rect 51859 2397 51871 2431
rect 52273 2431 52331 2437
rect 52273 2428 52285 2431
rect 51813 2391 51871 2397
rect 52196 2400 52285 2428
rect 52196 2304 52224 2400
rect 52273 2397 52285 2400
rect 52319 2397 52331 2431
rect 53745 2431 53803 2437
rect 53745 2428 53757 2431
rect 52273 2391 52331 2397
rect 53484 2400 53757 2428
rect 53484 2304 53512 2400
rect 53745 2397 53757 2400
rect 53791 2397 53803 2431
rect 54849 2431 54907 2437
rect 54849 2428 54861 2431
rect 53745 2391 53803 2397
rect 54772 2400 54861 2428
rect 54772 2304 54800 2400
rect 54849 2397 54861 2400
rect 54895 2397 54907 2431
rect 56321 2431 56379 2437
rect 56321 2428 56333 2431
rect 54849 2391 54907 2397
rect 56060 2400 56333 2428
rect 56060 2304 56088 2400
rect 56321 2397 56333 2400
rect 56367 2397 56379 2431
rect 57609 2431 57667 2437
rect 57609 2428 57621 2431
rect 56321 2391 56379 2397
rect 57348 2400 57621 2428
rect 57348 2304 57376 2400
rect 57609 2397 57621 2400
rect 57655 2397 57667 2431
rect 58069 2431 58127 2437
rect 58069 2428 58081 2431
rect 57609 2391 57667 2397
rect 57992 2400 58081 2428
rect 57992 2304 58020 2400
rect 58069 2397 58081 2400
rect 58115 2397 58127 2431
rect 59357 2431 59415 2437
rect 59357 2428 59369 2431
rect 58069 2391 58127 2397
rect 59280 2400 59369 2428
rect 59280 2304 59308 2400
rect 59357 2397 59369 2400
rect 59403 2397 59415 2431
rect 60645 2431 60703 2437
rect 60645 2428 60657 2431
rect 59357 2391 59415 2397
rect 60568 2400 60657 2428
rect 60568 2304 60596 2400
rect 60645 2397 60657 2400
rect 60691 2397 60703 2431
rect 62117 2431 62175 2437
rect 62117 2428 62129 2431
rect 60645 2391 60703 2397
rect 61856 2400 62129 2428
rect 61856 2304 61884 2400
rect 62117 2397 62129 2400
rect 62163 2397 62175 2431
rect 63405 2431 63463 2437
rect 63405 2428 63417 2431
rect 62117 2391 62175 2397
rect 63144 2400 63417 2428
rect 63144 2304 63172 2400
rect 63405 2397 63417 2400
rect 63451 2397 63463 2431
rect 63865 2431 63923 2437
rect 63865 2428 63877 2431
rect 63405 2391 63463 2397
rect 63788 2400 63877 2428
rect 63788 2304 63816 2400
rect 63865 2397 63877 2400
rect 63911 2397 63923 2431
rect 65153 2431 65211 2437
rect 65153 2428 65165 2431
rect 63865 2391 63923 2397
rect 65076 2400 65165 2428
rect 65076 2304 65104 2400
rect 65153 2397 65165 2400
rect 65199 2397 65211 2431
rect 65153 2391 65211 2397
rect 66441 2431 66499 2437
rect 66441 2397 66453 2431
rect 66487 2397 66499 2431
rect 67913 2431 67971 2437
rect 67913 2428 67925 2431
rect 66441 2391 66499 2397
rect 67652 2400 67925 2428
rect 25774 2252 25780 2304
rect 25832 2252 25838 2304
rect 31570 2252 31576 2304
rect 31628 2252 31634 2304
rect 32858 2252 32864 2304
rect 32916 2252 32922 2304
rect 33502 2252 33508 2304
rect 33560 2252 33566 2304
rect 34790 2252 34796 2304
rect 34848 2252 34854 2304
rect 36078 2252 36084 2304
rect 36136 2252 36142 2304
rect 37366 2252 37372 2304
rect 37424 2252 37430 2304
rect 38010 2252 38016 2304
rect 38068 2252 38074 2304
rect 39942 2252 39948 2304
rect 40000 2252 40006 2304
rect 40586 2252 40592 2304
rect 40644 2252 40650 2304
rect 41874 2252 41880 2304
rect 41932 2252 41938 2304
rect 43162 2252 43168 2304
rect 43220 2252 43226 2304
rect 44450 2252 44456 2304
rect 44508 2252 44514 2304
rect 45738 2252 45744 2304
rect 45796 2252 45802 2304
rect 46382 2252 46388 2304
rect 46440 2252 46446 2304
rect 47670 2252 47676 2304
rect 47728 2252 47734 2304
rect 48958 2252 48964 2304
rect 49016 2252 49022 2304
rect 50246 2252 50252 2304
rect 50304 2252 50310 2304
rect 51534 2252 51540 2304
rect 51592 2252 51598 2304
rect 52178 2252 52184 2304
rect 52236 2252 52242 2304
rect 53466 2252 53472 2304
rect 53524 2252 53530 2304
rect 54754 2252 54760 2304
rect 54812 2252 54818 2304
rect 56042 2252 56048 2304
rect 56100 2252 56106 2304
rect 57330 2252 57336 2304
rect 57388 2252 57394 2304
rect 57974 2252 57980 2304
rect 58032 2252 58038 2304
rect 59262 2252 59268 2304
rect 59320 2252 59326 2304
rect 60550 2252 60556 2304
rect 60608 2252 60614 2304
rect 61838 2252 61844 2304
rect 61896 2252 61902 2304
rect 63126 2252 63132 2304
rect 63184 2252 63190 2304
rect 63770 2252 63776 2304
rect 63828 2252 63834 2304
rect 65058 2252 65064 2304
rect 65116 2252 65122 2304
rect 66349 2295 66407 2301
rect 66349 2261 66361 2295
rect 66395 2292 66407 2295
rect 66456 2292 66484 2391
rect 67652 2304 67680 2400
rect 67913 2397 67925 2400
rect 67959 2397 67971 2431
rect 67913 2391 67971 2397
rect 66714 2292 66720 2304
rect 66395 2264 66720 2292
rect 66395 2261 66407 2264
rect 66349 2255 66407 2261
rect 66714 2252 66720 2264
rect 66772 2252 66778 2304
rect 67634 2252 67640 2304
rect 67692 2252 67698 2304
rect 1104 2202 118864 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 66314 2202
rect 66366 2150 66378 2202
rect 66430 2150 66442 2202
rect 66494 2150 66506 2202
rect 66558 2150 66570 2202
rect 66622 2150 97034 2202
rect 97086 2150 97098 2202
rect 97150 2150 97162 2202
rect 97214 2150 97226 2202
rect 97278 2150 97290 2202
rect 97342 2150 118864 2202
rect 1104 2128 118864 2150
<< via1 >>
rect 4214 97350 4266 97402
rect 4278 97350 4330 97402
rect 4342 97350 4394 97402
rect 4406 97350 4458 97402
rect 4470 97350 4522 97402
rect 34934 97350 34986 97402
rect 34998 97350 35050 97402
rect 35062 97350 35114 97402
rect 35126 97350 35178 97402
rect 35190 97350 35242 97402
rect 65654 97350 65706 97402
rect 65718 97350 65770 97402
rect 65782 97350 65834 97402
rect 65846 97350 65898 97402
rect 65910 97350 65962 97402
rect 96374 97350 96426 97402
rect 96438 97350 96490 97402
rect 96502 97350 96554 97402
rect 96566 97350 96618 97402
rect 96630 97350 96682 97402
rect 55772 97248 55824 97300
rect 57704 97248 57756 97300
rect 58808 97291 58860 97300
rect 58808 97257 58817 97291
rect 58817 97257 58851 97291
rect 58851 97257 58860 97291
rect 58808 97248 58860 97257
rect 60096 97291 60148 97300
rect 60096 97257 60105 97291
rect 60105 97257 60139 97291
rect 60139 97257 60148 97291
rect 60096 97248 60148 97257
rect 60648 97248 60700 97300
rect 62672 97291 62724 97300
rect 62672 97257 62681 97291
rect 62681 97257 62715 97291
rect 62715 97257 62724 97291
rect 62672 97248 62724 97257
rect 63316 97291 63368 97300
rect 63316 97257 63325 97291
rect 63325 97257 63359 97291
rect 63359 97257 63368 97291
rect 63316 97248 63368 97257
rect 64604 97291 64656 97300
rect 64604 97257 64613 97291
rect 64613 97257 64647 97291
rect 64647 97257 64656 97291
rect 64604 97248 64656 97257
rect 65248 97291 65300 97300
rect 65248 97257 65257 97291
rect 65257 97257 65291 97291
rect 65291 97257 65300 97291
rect 65248 97248 65300 97257
rect 65340 97248 65392 97300
rect 107844 97248 107896 97300
rect 67180 97223 67232 97232
rect 67180 97189 67189 97223
rect 67189 97189 67223 97223
rect 67223 97189 67232 97223
rect 67180 97180 67232 97189
rect 67824 97223 67876 97232
rect 67824 97189 67833 97223
rect 67833 97189 67867 97223
rect 67867 97189 67876 97223
rect 67824 97180 67876 97189
rect 70308 97180 70360 97232
rect 71688 97223 71740 97232
rect 71688 97189 71697 97223
rect 71697 97189 71731 97223
rect 71731 97189 71740 97223
rect 71688 97180 71740 97189
rect 72332 97223 72384 97232
rect 72332 97189 72341 97223
rect 72341 97189 72375 97223
rect 72375 97189 72384 97223
rect 72332 97180 72384 97189
rect 74356 97223 74408 97232
rect 74356 97189 74365 97223
rect 74365 97189 74399 97223
rect 74399 97189 74408 97223
rect 74356 97180 74408 97189
rect 107476 97223 107528 97232
rect 107476 97189 107485 97223
rect 107485 97189 107519 97223
rect 107519 97189 107528 97223
rect 107476 97180 107528 97189
rect 67640 97112 67692 97164
rect 57428 97044 57480 97096
rect 58164 97087 58216 97096
rect 58164 97053 58173 97087
rect 58173 97053 58207 97087
rect 58207 97053 58216 97087
rect 58164 97044 58216 97053
rect 59268 97044 59320 97096
rect 60556 97044 60608 97096
rect 60924 97087 60976 97096
rect 60924 97053 60933 97087
rect 60933 97053 60967 97087
rect 60967 97053 60976 97087
rect 60924 97044 60976 97053
rect 62856 97087 62908 97096
rect 62856 97053 62865 97087
rect 62865 97053 62899 97087
rect 62899 97053 62908 97087
rect 62856 97044 62908 97053
rect 63500 97087 63552 97096
rect 63500 97053 63509 97087
rect 63509 97053 63543 97087
rect 63543 97053 63552 97087
rect 63500 97044 63552 97053
rect 64972 97044 65024 97096
rect 66720 97044 66772 97096
rect 67364 97087 67416 97096
rect 67364 97053 67373 97087
rect 67373 97053 67407 97087
rect 67407 97053 67416 97087
rect 67364 97044 67416 97053
rect 68008 97087 68060 97096
rect 68008 97053 68017 97087
rect 68017 97053 68051 97087
rect 68051 97053 68060 97087
rect 68008 97044 68060 97053
rect 70032 97044 70084 97096
rect 71872 97087 71924 97096
rect 71872 97053 71881 97087
rect 71881 97053 71915 97087
rect 71915 97053 71924 97087
rect 71872 97044 71924 97053
rect 72516 97087 72568 97096
rect 72516 97053 72525 97087
rect 72525 97053 72559 97087
rect 72559 97053 72568 97087
rect 72516 97044 72568 97053
rect 74172 97087 74224 97096
rect 74172 97053 74181 97087
rect 74181 97053 74215 97087
rect 74215 97053 74224 97087
rect 74172 97044 74224 97053
rect 56600 96976 56652 97028
rect 67456 96976 67508 97028
rect 56232 96908 56284 96960
rect 67640 96951 67692 96960
rect 67640 96917 67649 96951
rect 67649 96917 67683 96951
rect 67683 96917 67692 96951
rect 67640 96908 67692 96917
rect 107844 96951 107896 96960
rect 107844 96917 107853 96951
rect 107853 96917 107887 96951
rect 107887 96917 107896 96951
rect 107844 96908 107896 96917
rect 4874 96806 4926 96858
rect 4938 96806 4990 96858
rect 5002 96806 5054 96858
rect 5066 96806 5118 96858
rect 5130 96806 5182 96858
rect 35594 96806 35646 96858
rect 35658 96806 35710 96858
rect 35722 96806 35774 96858
rect 35786 96806 35838 96858
rect 35850 96806 35902 96858
rect 66314 96806 66366 96858
rect 66378 96806 66430 96858
rect 66442 96806 66494 96858
rect 66506 96806 66558 96858
rect 66570 96806 66622 96858
rect 97034 96806 97086 96858
rect 97098 96806 97150 96858
rect 97162 96806 97214 96858
rect 97226 96806 97278 96858
rect 97290 96806 97342 96858
rect 56232 96679 56284 96688
rect 56232 96645 56241 96679
rect 56241 96645 56275 96679
rect 56275 96645 56284 96679
rect 56232 96636 56284 96645
rect 56784 96636 56836 96688
rect 69296 96611 69348 96620
rect 69296 96577 69305 96611
rect 69305 96577 69339 96611
rect 69339 96577 69348 96611
rect 69296 96568 69348 96577
rect 68836 96432 68888 96484
rect 4214 96262 4266 96314
rect 4278 96262 4330 96314
rect 4342 96262 4394 96314
rect 4406 96262 4458 96314
rect 4470 96262 4522 96314
rect 34934 96262 34986 96314
rect 34998 96262 35050 96314
rect 35062 96262 35114 96314
rect 35126 96262 35178 96314
rect 35190 96262 35242 96314
rect 65654 96262 65706 96314
rect 65718 96262 65770 96314
rect 65782 96262 65834 96314
rect 65846 96262 65898 96314
rect 65910 96262 65962 96314
rect 96374 96262 96426 96314
rect 96438 96262 96490 96314
rect 96502 96262 96554 96314
rect 96566 96262 96618 96314
rect 96630 96262 96682 96314
rect 58164 96160 58216 96212
rect 68008 96160 68060 96212
rect 74172 96160 74224 96212
rect 67456 96092 67508 96144
rect 56784 96067 56836 96076
rect 56784 96033 56793 96067
rect 56793 96033 56827 96067
rect 56827 96033 56836 96067
rect 56784 96024 56836 96033
rect 70768 95956 70820 96008
rect 57060 95931 57112 95940
rect 57060 95897 57069 95931
rect 57069 95897 57103 95931
rect 57103 95897 57112 95931
rect 57060 95888 57112 95897
rect 59176 95888 59228 95940
rect 69112 95888 69164 95940
rect 71964 95931 72016 95940
rect 71964 95897 71973 95931
rect 71973 95897 72007 95931
rect 72007 95897 72016 95931
rect 71964 95888 72016 95897
rect 74724 95888 74776 95940
rect 66996 95820 67048 95872
rect 4874 95718 4926 95770
rect 4938 95718 4990 95770
rect 5002 95718 5054 95770
rect 5066 95718 5118 95770
rect 5130 95718 5182 95770
rect 35594 95718 35646 95770
rect 35658 95718 35710 95770
rect 35722 95718 35774 95770
rect 35786 95718 35838 95770
rect 35850 95718 35902 95770
rect 66314 95718 66366 95770
rect 66378 95718 66430 95770
rect 66442 95718 66494 95770
rect 66506 95718 66558 95770
rect 66570 95718 66622 95770
rect 97034 95718 97086 95770
rect 97098 95718 97150 95770
rect 97162 95718 97214 95770
rect 97226 95718 97278 95770
rect 97290 95718 97342 95770
rect 57428 95659 57480 95668
rect 57428 95625 57437 95659
rect 57437 95625 57471 95659
rect 57471 95625 57480 95659
rect 57428 95616 57480 95625
rect 60924 95616 60976 95668
rect 54484 95548 54536 95600
rect 57704 95548 57756 95600
rect 57612 95480 57664 95532
rect 62764 95616 62816 95668
rect 62856 95659 62908 95668
rect 62856 95625 62865 95659
rect 62865 95625 62899 95659
rect 62899 95625 62908 95659
rect 62856 95616 62908 95625
rect 64880 95616 64932 95668
rect 64972 95659 65024 95668
rect 64972 95625 64981 95659
rect 64981 95625 65015 95659
rect 65015 95625 65024 95659
rect 64972 95616 65024 95625
rect 66628 95616 66680 95668
rect 66720 95616 66772 95668
rect 67088 95548 67140 95600
rect 69940 95548 69992 95600
rect 71872 95616 71924 95668
rect 70584 95548 70636 95600
rect 71688 95548 71740 95600
rect 55680 95455 55732 95464
rect 55680 95421 55689 95455
rect 55689 95421 55723 95455
rect 55723 95421 55732 95455
rect 55680 95412 55732 95421
rect 57888 95412 57940 95464
rect 59544 95276 59596 95328
rect 60740 95344 60792 95396
rect 63592 95412 63644 95464
rect 65064 95455 65116 95464
rect 62028 95276 62080 95328
rect 65064 95421 65073 95455
rect 65073 95421 65107 95455
rect 65107 95421 65116 95455
rect 65064 95412 65116 95421
rect 64788 95344 64840 95396
rect 67732 95412 67784 95464
rect 69020 95412 69072 95464
rect 70032 95344 70084 95396
rect 4214 95174 4266 95226
rect 4278 95174 4330 95226
rect 4342 95174 4394 95226
rect 4406 95174 4458 95226
rect 4470 95174 4522 95226
rect 34934 95174 34986 95226
rect 34998 95174 35050 95226
rect 35062 95174 35114 95226
rect 35126 95174 35178 95226
rect 35190 95174 35242 95226
rect 65654 95174 65706 95226
rect 65718 95174 65770 95226
rect 65782 95174 65834 95226
rect 65846 95174 65898 95226
rect 65910 95174 65962 95226
rect 96374 95174 96426 95226
rect 96438 95174 96490 95226
rect 96502 95174 96554 95226
rect 96566 95174 96618 95226
rect 96630 95174 96682 95226
rect 59268 95072 59320 95124
rect 63500 95072 63552 95124
rect 67364 95115 67416 95124
rect 67364 95081 67373 95115
rect 67373 95081 67407 95115
rect 67407 95081 67416 95115
rect 67364 95072 67416 95081
rect 69296 95072 69348 95124
rect 72516 95115 72568 95124
rect 72516 95081 72525 95115
rect 72525 95081 72559 95115
rect 72559 95081 72568 95115
rect 72516 95072 72568 95081
rect 54668 94936 54720 94988
rect 56784 94936 56836 94988
rect 57888 94979 57940 94988
rect 57888 94945 57897 94979
rect 57897 94945 57931 94979
rect 57931 94945 57940 94979
rect 57888 94936 57940 94945
rect 62028 94979 62080 94988
rect 62028 94945 62037 94979
rect 62037 94945 62071 94979
rect 62071 94945 62080 94979
rect 62028 94936 62080 94945
rect 65064 94936 65116 94988
rect 66904 94936 66956 94988
rect 67456 94979 67508 94988
rect 67456 94945 67465 94979
rect 67465 94945 67499 94979
rect 67499 94945 67508 94979
rect 67456 94936 67508 94945
rect 56876 94868 56928 94920
rect 66996 94868 67048 94920
rect 68836 94868 68888 94920
rect 70768 94911 70820 94920
rect 70768 94877 70777 94911
rect 70777 94877 70811 94911
rect 70811 94877 70820 94911
rect 70768 94868 70820 94877
rect 57796 94800 57848 94852
rect 55220 94732 55272 94784
rect 61752 94800 61804 94852
rect 62304 94843 62356 94852
rect 62304 94809 62313 94843
rect 62313 94809 62347 94843
rect 62347 94809 62356 94843
rect 62304 94800 62356 94809
rect 65248 94800 65300 94852
rect 64144 94732 64196 94784
rect 67180 94800 67232 94852
rect 69756 94800 69808 94852
rect 72976 94800 73028 94852
rect 4874 94630 4926 94682
rect 4938 94630 4990 94682
rect 5002 94630 5054 94682
rect 5066 94630 5118 94682
rect 5130 94630 5182 94682
rect 35594 94630 35646 94682
rect 35658 94630 35710 94682
rect 35722 94630 35774 94682
rect 35786 94630 35838 94682
rect 35850 94630 35902 94682
rect 66314 94630 66366 94682
rect 66378 94630 66430 94682
rect 66442 94630 66494 94682
rect 66506 94630 66558 94682
rect 66570 94630 66622 94682
rect 97034 94630 97086 94682
rect 97098 94630 97150 94682
rect 97162 94630 97214 94682
rect 97226 94630 97278 94682
rect 97290 94630 97342 94682
rect 57060 94528 57112 94580
rect 60004 94528 60056 94580
rect 60556 94528 60608 94580
rect 61752 94571 61804 94580
rect 61752 94537 61761 94571
rect 61761 94537 61795 94571
rect 61795 94537 61804 94571
rect 61752 94528 61804 94537
rect 65248 94528 65300 94580
rect 57704 94460 57756 94512
rect 52460 94392 52512 94444
rect 55496 94392 55548 94444
rect 55680 94392 55732 94444
rect 55864 94435 55916 94444
rect 55864 94401 55898 94435
rect 55898 94401 55916 94435
rect 55864 94392 55916 94401
rect 58440 94435 58492 94444
rect 58440 94401 58449 94435
rect 58449 94401 58483 94435
rect 58483 94401 58492 94435
rect 58440 94392 58492 94401
rect 60096 94460 60148 94512
rect 63224 94460 63276 94512
rect 59544 94435 59596 94444
rect 59544 94401 59553 94435
rect 59553 94401 59587 94435
rect 59587 94401 59596 94435
rect 59544 94392 59596 94401
rect 53840 94324 53892 94376
rect 54668 94367 54720 94376
rect 54668 94333 54677 94367
rect 54677 94333 54711 94367
rect 54711 94333 54720 94367
rect 54668 94324 54720 94333
rect 55404 94324 55456 94376
rect 56876 94324 56928 94376
rect 57888 94324 57940 94376
rect 60188 94324 60240 94376
rect 63316 94324 63368 94376
rect 55588 94188 55640 94240
rect 55864 94188 55916 94240
rect 63776 94256 63828 94308
rect 65432 94435 65484 94444
rect 65432 94401 65441 94435
rect 65441 94401 65475 94435
rect 65475 94401 65484 94435
rect 65432 94392 65484 94401
rect 70492 94256 70544 94308
rect 63592 94188 63644 94240
rect 4214 94086 4266 94138
rect 4278 94086 4330 94138
rect 4342 94086 4394 94138
rect 4406 94086 4458 94138
rect 4470 94086 4522 94138
rect 34934 94086 34986 94138
rect 34998 94086 35050 94138
rect 35062 94086 35114 94138
rect 35126 94086 35178 94138
rect 35190 94086 35242 94138
rect 65654 94086 65706 94138
rect 65718 94086 65770 94138
rect 65782 94086 65834 94138
rect 65846 94086 65898 94138
rect 65910 94086 65962 94138
rect 96374 94086 96426 94138
rect 96438 94086 96490 94138
rect 96502 94086 96554 94138
rect 96566 94086 96618 94138
rect 96630 94086 96682 94138
rect 57796 94027 57848 94036
rect 57796 93993 57805 94027
rect 57805 93993 57839 94027
rect 57839 93993 57848 94027
rect 57796 93984 57848 93993
rect 57888 93984 57940 94036
rect 55588 93959 55640 93968
rect 55588 93925 55597 93959
rect 55597 93925 55631 93959
rect 55631 93925 55640 93959
rect 55588 93916 55640 93925
rect 60740 93984 60792 94036
rect 64144 94027 64196 94036
rect 64144 93993 64153 94027
rect 64153 93993 64187 94027
rect 64187 93993 64196 94027
rect 64144 93984 64196 93993
rect 67180 93984 67232 94036
rect 68836 93984 68888 94036
rect 65432 93916 65484 93968
rect 63592 93891 63644 93900
rect 63592 93857 63601 93891
rect 63601 93857 63635 93891
rect 63635 93857 63644 93891
rect 63592 93848 63644 93857
rect 66168 93848 66220 93900
rect 55496 93780 55548 93832
rect 56508 93780 56560 93832
rect 59544 93780 59596 93832
rect 59636 93823 59688 93832
rect 59636 93789 59645 93823
rect 59645 93789 59679 93823
rect 59679 93789 59688 93823
rect 59636 93780 59688 93789
rect 60096 93780 60148 93832
rect 61476 93780 61528 93832
rect 61660 93780 61712 93832
rect 62764 93780 62816 93832
rect 63316 93780 63368 93832
rect 63776 93823 63828 93832
rect 63776 93789 63785 93823
rect 63785 93789 63819 93823
rect 63819 93789 63828 93823
rect 63776 93780 63828 93789
rect 64696 93780 64748 93832
rect 64880 93780 64932 93832
rect 65432 93780 65484 93832
rect 65892 93823 65944 93832
rect 65892 93789 65901 93823
rect 65901 93789 65935 93823
rect 65935 93789 65944 93823
rect 65892 93780 65944 93789
rect 67088 93823 67140 93832
rect 67088 93789 67097 93823
rect 67097 93789 67131 93823
rect 67131 93789 67140 93823
rect 67088 93780 67140 93789
rect 53380 93644 53432 93696
rect 58164 93712 58216 93764
rect 55772 93687 55824 93696
rect 55772 93653 55781 93687
rect 55781 93653 55815 93687
rect 55815 93653 55824 93687
rect 55772 93644 55824 93653
rect 59268 93712 59320 93764
rect 60372 93712 60424 93764
rect 59360 93644 59412 93696
rect 60648 93644 60700 93696
rect 62304 93712 62356 93764
rect 61384 93644 61436 93696
rect 61752 93687 61804 93696
rect 61752 93653 61761 93687
rect 61761 93653 61795 93687
rect 61795 93653 61804 93687
rect 61752 93644 61804 93653
rect 63500 93712 63552 93764
rect 62856 93644 62908 93696
rect 64788 93712 64840 93764
rect 64512 93644 64564 93696
rect 64604 93644 64656 93696
rect 66812 93712 66864 93764
rect 67272 93712 67324 93764
rect 68284 93712 68336 93764
rect 69112 93823 69164 93832
rect 69112 93789 69121 93823
rect 69121 93789 69155 93823
rect 69155 93789 69164 93823
rect 69112 93780 69164 93789
rect 72240 93780 72292 93832
rect 70124 93712 70176 93764
rect 70492 93755 70544 93764
rect 70492 93721 70501 93755
rect 70501 93721 70535 93755
rect 70535 93721 70544 93755
rect 70492 93712 70544 93721
rect 65984 93687 66036 93696
rect 65984 93653 65993 93687
rect 65993 93653 66027 93687
rect 66027 93653 66036 93687
rect 65984 93644 66036 93653
rect 66720 93644 66772 93696
rect 66996 93644 67048 93696
rect 70860 93687 70912 93696
rect 70860 93653 70869 93687
rect 70869 93653 70903 93687
rect 70903 93653 70912 93687
rect 70860 93644 70912 93653
rect 71136 93687 71188 93696
rect 71136 93653 71145 93687
rect 71145 93653 71179 93687
rect 71179 93653 71188 93687
rect 71136 93644 71188 93653
rect 72148 93644 72200 93696
rect 4874 93542 4926 93594
rect 4938 93542 4990 93594
rect 5002 93542 5054 93594
rect 5066 93542 5118 93594
rect 5130 93542 5182 93594
rect 35594 93542 35646 93594
rect 35658 93542 35710 93594
rect 35722 93542 35774 93594
rect 35786 93542 35838 93594
rect 35850 93542 35902 93594
rect 66314 93542 66366 93594
rect 66378 93542 66430 93594
rect 66442 93542 66494 93594
rect 66506 93542 66558 93594
rect 66570 93542 66622 93594
rect 97034 93542 97086 93594
rect 97098 93542 97150 93594
rect 97162 93542 97214 93594
rect 97226 93542 97278 93594
rect 97290 93542 97342 93594
rect 54484 93483 54536 93492
rect 54484 93449 54493 93483
rect 54493 93449 54527 93483
rect 54527 93449 54536 93483
rect 54484 93440 54536 93449
rect 57612 93440 57664 93492
rect 55772 93372 55824 93424
rect 56232 93372 56284 93424
rect 59636 93440 59688 93492
rect 60004 93483 60056 93492
rect 60004 93449 60013 93483
rect 60013 93449 60047 93483
rect 60047 93449 60056 93483
rect 60004 93440 60056 93449
rect 60648 93440 60700 93492
rect 61568 93440 61620 93492
rect 63500 93440 63552 93492
rect 65984 93440 66036 93492
rect 69848 93440 69900 93492
rect 69940 93440 69992 93492
rect 70860 93440 70912 93492
rect 71688 93440 71740 93492
rect 72976 93483 73028 93492
rect 72976 93449 72985 93483
rect 72985 93449 73019 93483
rect 73019 93449 73028 93483
rect 72976 93440 73028 93449
rect 74724 93483 74776 93492
rect 74724 93449 74733 93483
rect 74733 93449 74767 93483
rect 74767 93449 74776 93483
rect 74724 93440 74776 93449
rect 58900 93372 58952 93424
rect 59544 93372 59596 93424
rect 49332 93304 49384 93356
rect 46848 93236 46900 93288
rect 49516 93279 49568 93288
rect 49516 93245 49525 93279
rect 49525 93245 49559 93279
rect 49559 93245 49568 93279
rect 49516 93236 49568 93245
rect 49332 93211 49384 93220
rect 49332 93177 49341 93211
rect 49341 93177 49375 93211
rect 49375 93177 49384 93211
rect 49332 93168 49384 93177
rect 46940 93100 46992 93152
rect 54668 93347 54720 93356
rect 54668 93313 54677 93347
rect 54677 93313 54711 93347
rect 54711 93313 54720 93347
rect 56600 93347 56652 93356
rect 54668 93304 54720 93313
rect 56600 93313 56609 93347
rect 56609 93313 56643 93347
rect 56643 93313 56652 93347
rect 56600 93304 56652 93313
rect 53840 93279 53892 93288
rect 53840 93245 53849 93279
rect 53849 93245 53883 93279
rect 53883 93245 53892 93279
rect 53840 93236 53892 93245
rect 53932 93236 53984 93288
rect 56324 93236 56376 93288
rect 56508 93236 56560 93288
rect 59820 93304 59872 93356
rect 60740 93372 60792 93424
rect 63592 93372 63644 93424
rect 56876 93236 56928 93288
rect 63224 93347 63276 93356
rect 63224 93313 63233 93347
rect 63233 93313 63267 93347
rect 63267 93313 63276 93347
rect 63224 93304 63276 93313
rect 63316 93347 63368 93356
rect 63316 93313 63325 93347
rect 63325 93313 63359 93347
rect 63359 93313 63368 93347
rect 63316 93304 63368 93313
rect 66904 93372 66956 93424
rect 68376 93372 68428 93424
rect 52184 93100 52236 93152
rect 56232 93100 56284 93152
rect 56324 93100 56376 93152
rect 60372 93100 60424 93152
rect 60464 93100 60516 93152
rect 61660 93100 61712 93152
rect 63776 93236 63828 93288
rect 65248 93236 65300 93288
rect 66352 93304 66404 93356
rect 66720 93347 66772 93356
rect 66720 93313 66729 93347
rect 66729 93313 66763 93347
rect 66763 93313 66772 93347
rect 66720 93304 66772 93313
rect 67824 93304 67876 93356
rect 64788 93168 64840 93220
rect 68376 93279 68428 93288
rect 68376 93245 68385 93279
rect 68385 93245 68419 93279
rect 68419 93245 68428 93279
rect 68376 93236 68428 93245
rect 70124 93372 70176 93424
rect 72056 93372 72108 93424
rect 72240 93415 72292 93424
rect 72240 93381 72249 93415
rect 72249 93381 72283 93415
rect 72283 93381 72292 93415
rect 72240 93372 72292 93381
rect 69204 93304 69256 93356
rect 70308 93347 70360 93356
rect 70308 93313 70317 93347
rect 70317 93313 70351 93347
rect 70351 93313 70360 93347
rect 70308 93304 70360 93313
rect 62856 93100 62908 93152
rect 63408 93100 63460 93152
rect 66812 93168 66864 93220
rect 67732 93168 67784 93220
rect 69940 93236 69992 93288
rect 70124 93279 70176 93288
rect 70124 93245 70133 93279
rect 70133 93245 70167 93279
rect 70167 93245 70176 93279
rect 70124 93236 70176 93245
rect 72148 93279 72200 93288
rect 72148 93245 72157 93279
rect 72157 93245 72191 93279
rect 72191 93245 72200 93279
rect 72148 93236 72200 93245
rect 74172 93236 74224 93288
rect 68560 93100 68612 93152
rect 69020 93100 69072 93152
rect 69756 93143 69808 93152
rect 69756 93109 69765 93143
rect 69765 93109 69799 93143
rect 69799 93109 69808 93143
rect 69756 93100 69808 93109
rect 69848 93100 69900 93152
rect 70584 93100 70636 93152
rect 71964 93100 72016 93152
rect 107844 93168 107896 93220
rect 108580 93100 108632 93152
rect 4214 92998 4266 93050
rect 4278 92998 4330 93050
rect 4342 92998 4394 93050
rect 4406 92998 4458 93050
rect 4470 92998 4522 93050
rect 34934 92998 34986 93050
rect 34998 92998 35050 93050
rect 35062 92998 35114 93050
rect 35126 92998 35178 93050
rect 35190 92998 35242 93050
rect 65654 92998 65706 93050
rect 65718 92998 65770 93050
rect 65782 92998 65834 93050
rect 65846 92998 65898 93050
rect 65910 92998 65962 93050
rect 96374 92998 96426 93050
rect 96438 92998 96490 93050
rect 96502 92998 96554 93050
rect 96566 92998 96618 93050
rect 96630 92998 96682 93050
rect 46940 92939 46992 92948
rect 46940 92905 46949 92939
rect 46949 92905 46983 92939
rect 46983 92905 46992 92939
rect 46940 92896 46992 92905
rect 52184 92939 52236 92948
rect 52184 92905 52193 92939
rect 52193 92905 52227 92939
rect 52227 92905 52236 92939
rect 52184 92896 52236 92905
rect 52460 92896 52512 92948
rect 53932 92896 53984 92948
rect 55404 92896 55456 92948
rect 61292 92896 61344 92948
rect 61384 92896 61436 92948
rect 63408 92896 63460 92948
rect 63500 92939 63552 92948
rect 63500 92905 63509 92939
rect 63509 92905 63543 92939
rect 63543 92905 63552 92939
rect 63500 92896 63552 92905
rect 60464 92828 60516 92880
rect 62948 92828 63000 92880
rect 64604 92828 64656 92880
rect 70308 92896 70360 92948
rect 70584 92896 70636 92948
rect 46848 92760 46900 92812
rect 50620 92803 50672 92812
rect 50620 92769 50629 92803
rect 50629 92769 50663 92803
rect 50663 92769 50672 92803
rect 50620 92760 50672 92769
rect 57980 92803 58032 92812
rect 57980 92769 57989 92803
rect 57989 92769 58023 92803
rect 58023 92769 58032 92803
rect 57980 92760 58032 92769
rect 63592 92803 63644 92812
rect 63592 92769 63601 92803
rect 63601 92769 63635 92803
rect 63635 92769 63644 92803
rect 63592 92760 63644 92769
rect 68560 92871 68612 92880
rect 68560 92837 68569 92871
rect 68569 92837 68603 92871
rect 68603 92837 68612 92871
rect 68560 92828 68612 92837
rect 69940 92828 69992 92880
rect 45652 92692 45704 92744
rect 44180 92624 44232 92676
rect 47124 92624 47176 92676
rect 53380 92692 53432 92744
rect 52552 92667 52604 92676
rect 52552 92633 52586 92667
rect 52586 92633 52604 92667
rect 52552 92624 52604 92633
rect 54024 92667 54076 92676
rect 54024 92633 54058 92667
rect 54058 92633 54076 92667
rect 56508 92692 56560 92744
rect 58900 92692 58952 92744
rect 54024 92624 54076 92633
rect 58440 92667 58492 92676
rect 58440 92633 58474 92667
rect 58474 92633 58492 92667
rect 58440 92624 58492 92633
rect 59268 92624 59320 92676
rect 63224 92624 63276 92676
rect 63500 92624 63552 92676
rect 59452 92556 59504 92608
rect 61292 92556 61344 92608
rect 64880 92556 64932 92608
rect 72148 92735 72200 92744
rect 72148 92701 72157 92735
rect 72157 92701 72191 92735
rect 72191 92701 72200 92735
rect 72148 92692 72200 92701
rect 72976 92692 73028 92744
rect 67548 92624 67600 92676
rect 69204 92624 69256 92676
rect 69572 92624 69624 92676
rect 70492 92624 70544 92676
rect 73252 92624 73304 92676
rect 73712 92624 73764 92676
rect 77484 92667 77536 92676
rect 77484 92633 77493 92667
rect 77493 92633 77527 92667
rect 77527 92633 77536 92667
rect 77484 92624 77536 92633
rect 74724 92556 74776 92608
rect 79416 92599 79468 92608
rect 79416 92565 79425 92599
rect 79425 92565 79459 92599
rect 79459 92565 79468 92599
rect 79416 92556 79468 92565
rect 4874 92454 4926 92506
rect 4938 92454 4990 92506
rect 5002 92454 5054 92506
rect 5066 92454 5118 92506
rect 5130 92454 5182 92506
rect 35594 92454 35646 92506
rect 35658 92454 35710 92506
rect 35722 92454 35774 92506
rect 35786 92454 35838 92506
rect 35850 92454 35902 92506
rect 66314 92454 66366 92506
rect 66378 92454 66430 92506
rect 66442 92454 66494 92506
rect 66506 92454 66558 92506
rect 66570 92454 66622 92506
rect 97034 92454 97086 92506
rect 97098 92454 97150 92506
rect 97162 92454 97214 92506
rect 97226 92454 97278 92506
rect 97290 92454 97342 92506
rect 113650 92454 113702 92506
rect 113714 92454 113766 92506
rect 113778 92454 113830 92506
rect 113842 92454 113894 92506
rect 113906 92454 113958 92506
rect 45652 92395 45704 92404
rect 45652 92361 45661 92395
rect 45661 92361 45695 92395
rect 45695 92361 45704 92395
rect 45652 92352 45704 92361
rect 54668 92352 54720 92404
rect 52920 92284 52972 92336
rect 54852 92352 54904 92404
rect 58348 92352 58400 92404
rect 49516 92216 49568 92268
rect 53380 92259 53432 92268
rect 53380 92225 53389 92259
rect 53389 92225 53423 92259
rect 53423 92225 53432 92259
rect 53380 92216 53432 92225
rect 8208 92012 8260 92064
rect 45652 92012 45704 92064
rect 46848 92012 46900 92064
rect 53196 92148 53248 92200
rect 56048 92284 56100 92336
rect 63500 92395 63552 92404
rect 63500 92361 63509 92395
rect 63509 92361 63543 92395
rect 63543 92361 63552 92395
rect 63500 92352 63552 92361
rect 56416 92216 56468 92268
rect 58900 92259 58952 92268
rect 58900 92225 58909 92259
rect 58909 92225 58943 92259
rect 58943 92225 58952 92259
rect 58900 92216 58952 92225
rect 60740 92259 60792 92268
rect 60740 92225 60749 92259
rect 60749 92225 60783 92259
rect 60783 92225 60792 92259
rect 60740 92216 60792 92225
rect 65340 92395 65392 92404
rect 65340 92361 65349 92395
rect 65349 92361 65383 92395
rect 65383 92361 65392 92395
rect 65340 92352 65392 92361
rect 67640 92352 67692 92404
rect 72976 92395 73028 92404
rect 72976 92361 72985 92395
rect 72985 92361 73019 92395
rect 73019 92361 73028 92395
rect 72976 92352 73028 92361
rect 77484 92352 77536 92404
rect 69572 92216 69624 92268
rect 66720 92148 66772 92200
rect 50252 92123 50304 92132
rect 50252 92089 50261 92123
rect 50261 92089 50295 92123
rect 50295 92089 50304 92123
rect 50252 92080 50304 92089
rect 49608 92055 49660 92064
rect 49608 92021 49617 92055
rect 49617 92021 49651 92055
rect 49651 92021 49660 92055
rect 49608 92012 49660 92021
rect 53196 92055 53248 92064
rect 53196 92021 53205 92055
rect 53205 92021 53239 92055
rect 53239 92021 53248 92055
rect 53196 92012 53248 92021
rect 58716 92123 58768 92132
rect 58716 92089 58725 92123
rect 58725 92089 58759 92123
rect 58759 92089 58768 92123
rect 58716 92080 58768 92089
rect 60556 92123 60608 92132
rect 60556 92089 60565 92123
rect 60565 92089 60599 92123
rect 60599 92089 60608 92123
rect 60556 92080 60608 92089
rect 67824 92080 67876 92132
rect 68284 92123 68336 92132
rect 68284 92089 68293 92123
rect 68293 92089 68327 92123
rect 68327 92089 68336 92123
rect 68284 92080 68336 92089
rect 71872 92148 71924 92200
rect 74724 92259 74776 92268
rect 74724 92225 74733 92259
rect 74733 92225 74767 92259
rect 74767 92225 74776 92259
rect 74724 92216 74776 92225
rect 75920 92148 75972 92200
rect 70768 92080 70820 92132
rect 72056 92080 72108 92132
rect 54852 92012 54904 92064
rect 64696 92012 64748 92064
rect 79416 92012 79468 92064
rect 100024 92080 100076 92132
rect 89444 92055 89496 92064
rect 89444 92021 89453 92055
rect 89453 92021 89487 92055
rect 89487 92021 89496 92055
rect 89444 92012 89496 92021
rect 4214 91910 4266 91962
rect 4278 91910 4330 91962
rect 4342 91910 4394 91962
rect 4406 91910 4458 91962
rect 4470 91910 4522 91962
rect 34934 91910 34986 91962
rect 34998 91910 35050 91962
rect 35062 91910 35114 91962
rect 35126 91910 35178 91962
rect 35190 91910 35242 91962
rect 65654 91910 65706 91962
rect 65718 91910 65770 91962
rect 65782 91910 65834 91962
rect 65846 91910 65898 91962
rect 65910 91910 65962 91962
rect 96374 91910 96426 91962
rect 96438 91910 96490 91962
rect 96502 91910 96554 91962
rect 96566 91910 96618 91962
rect 96630 91910 96682 91962
rect 112914 91910 112966 91962
rect 112978 91910 113030 91962
rect 113042 91910 113094 91962
rect 113106 91910 113158 91962
rect 113170 91910 113222 91962
rect 49608 91808 49660 91860
rect 55220 91808 55272 91860
rect 56048 91808 56100 91860
rect 61752 91808 61804 91860
rect 77484 91740 77536 91792
rect 108304 91740 108356 91792
rect 4874 91366 4926 91418
rect 4938 91366 4990 91418
rect 5002 91366 5054 91418
rect 5066 91366 5118 91418
rect 5130 91366 5182 91418
rect 113650 91366 113702 91418
rect 113714 91366 113766 91418
rect 113778 91366 113830 91418
rect 113842 91366 113894 91418
rect 113906 91366 113958 91418
rect 4214 90822 4266 90874
rect 4278 90822 4330 90874
rect 4342 90822 4394 90874
rect 4406 90822 4458 90874
rect 4470 90822 4522 90874
rect 112914 90822 112966 90874
rect 112978 90822 113030 90874
rect 113042 90822 113094 90874
rect 113106 90822 113158 90874
rect 113170 90822 113222 90874
rect 71136 90380 71188 90432
rect 108396 90380 108448 90432
rect 4874 90278 4926 90330
rect 4938 90278 4990 90330
rect 5002 90278 5054 90330
rect 5066 90278 5118 90330
rect 5130 90278 5182 90330
rect 113650 90278 113702 90330
rect 113714 90278 113766 90330
rect 113778 90278 113830 90330
rect 113842 90278 113894 90330
rect 113906 90278 113958 90330
rect 4214 89734 4266 89786
rect 4278 89734 4330 89786
rect 4342 89734 4394 89786
rect 4406 89734 4458 89786
rect 4470 89734 4522 89786
rect 112914 89734 112966 89786
rect 112978 89734 113030 89786
rect 113042 89734 113094 89786
rect 113106 89734 113158 89786
rect 113170 89734 113222 89786
rect 4874 89190 4926 89242
rect 4938 89190 4990 89242
rect 5002 89190 5054 89242
rect 5066 89190 5118 89242
rect 5130 89190 5182 89242
rect 113650 89190 113702 89242
rect 113714 89190 113766 89242
rect 113778 89190 113830 89242
rect 113842 89190 113894 89242
rect 113906 89190 113958 89242
rect 4214 88646 4266 88698
rect 4278 88646 4330 88698
rect 4342 88646 4394 88698
rect 4406 88646 4458 88698
rect 4470 88646 4522 88698
rect 112914 88646 112966 88698
rect 112978 88646 113030 88698
rect 113042 88646 113094 88698
rect 113106 88646 113158 88698
rect 113170 88646 113222 88698
rect 4874 88102 4926 88154
rect 4938 88102 4990 88154
rect 5002 88102 5054 88154
rect 5066 88102 5118 88154
rect 5130 88102 5182 88154
rect 113650 88102 113702 88154
rect 113714 88102 113766 88154
rect 113778 88102 113830 88154
rect 113842 88102 113894 88154
rect 113906 88102 113958 88154
rect 4214 87558 4266 87610
rect 4278 87558 4330 87610
rect 4342 87558 4394 87610
rect 4406 87558 4458 87610
rect 4470 87558 4522 87610
rect 112914 87558 112966 87610
rect 112978 87558 113030 87610
rect 113042 87558 113094 87610
rect 113106 87558 113158 87610
rect 113170 87558 113222 87610
rect 4874 87014 4926 87066
rect 4938 87014 4990 87066
rect 5002 87014 5054 87066
rect 5066 87014 5118 87066
rect 5130 87014 5182 87066
rect 113650 87014 113702 87066
rect 113714 87014 113766 87066
rect 113778 87014 113830 87066
rect 113842 87014 113894 87066
rect 113906 87014 113958 87066
rect 106188 86572 106240 86624
rect 4214 86470 4266 86522
rect 4278 86470 4330 86522
rect 4342 86470 4394 86522
rect 4406 86470 4458 86522
rect 4470 86470 4522 86522
rect 112914 86470 112966 86522
rect 112978 86470 113030 86522
rect 113042 86470 113094 86522
rect 113106 86470 113158 86522
rect 113170 86470 113222 86522
rect 4874 85926 4926 85978
rect 4938 85926 4990 85978
rect 5002 85926 5054 85978
rect 5066 85926 5118 85978
rect 5130 85926 5182 85978
rect 113650 85926 113702 85978
rect 113714 85926 113766 85978
rect 113778 85926 113830 85978
rect 113842 85926 113894 85978
rect 113906 85926 113958 85978
rect 4214 85382 4266 85434
rect 4278 85382 4330 85434
rect 4342 85382 4394 85434
rect 4406 85382 4458 85434
rect 4470 85382 4522 85434
rect 112914 85382 112966 85434
rect 112978 85382 113030 85434
rect 113042 85382 113094 85434
rect 113106 85382 113158 85434
rect 113170 85382 113222 85434
rect 4874 84838 4926 84890
rect 4938 84838 4990 84890
rect 5002 84838 5054 84890
rect 5066 84838 5118 84890
rect 5130 84838 5182 84890
rect 113650 84838 113702 84890
rect 113714 84838 113766 84890
rect 113778 84838 113830 84890
rect 113842 84838 113894 84890
rect 113906 84838 113958 84890
rect 4214 84294 4266 84346
rect 4278 84294 4330 84346
rect 4342 84294 4394 84346
rect 4406 84294 4458 84346
rect 4470 84294 4522 84346
rect 112914 84294 112966 84346
rect 112978 84294 113030 84346
rect 113042 84294 113094 84346
rect 113106 84294 113158 84346
rect 113170 84294 113222 84346
rect 4874 83750 4926 83802
rect 4938 83750 4990 83802
rect 5002 83750 5054 83802
rect 5066 83750 5118 83802
rect 5130 83750 5182 83802
rect 113650 83750 113702 83802
rect 113714 83750 113766 83802
rect 113778 83750 113830 83802
rect 113842 83750 113894 83802
rect 113906 83750 113958 83802
rect 4214 83206 4266 83258
rect 4278 83206 4330 83258
rect 4342 83206 4394 83258
rect 4406 83206 4458 83258
rect 4470 83206 4522 83258
rect 112914 83206 112966 83258
rect 112978 83206 113030 83258
rect 113042 83206 113094 83258
rect 113106 83206 113158 83258
rect 113170 83206 113222 83258
rect 4874 82662 4926 82714
rect 4938 82662 4990 82714
rect 5002 82662 5054 82714
rect 5066 82662 5118 82714
rect 5130 82662 5182 82714
rect 113650 82662 113702 82714
rect 113714 82662 113766 82714
rect 113778 82662 113830 82714
rect 113842 82662 113894 82714
rect 113906 82662 113958 82714
rect 4214 82118 4266 82170
rect 4278 82118 4330 82170
rect 4342 82118 4394 82170
rect 4406 82118 4458 82170
rect 4470 82118 4522 82170
rect 112914 82118 112966 82170
rect 112978 82118 113030 82170
rect 113042 82118 113094 82170
rect 113106 82118 113158 82170
rect 113170 82118 113222 82170
rect 4874 81574 4926 81626
rect 4938 81574 4990 81626
rect 5002 81574 5054 81626
rect 5066 81574 5118 81626
rect 5130 81574 5182 81626
rect 113650 81574 113702 81626
rect 113714 81574 113766 81626
rect 113778 81574 113830 81626
rect 113842 81574 113894 81626
rect 113906 81574 113958 81626
rect 4214 81030 4266 81082
rect 4278 81030 4330 81082
rect 4342 81030 4394 81082
rect 4406 81030 4458 81082
rect 4470 81030 4522 81082
rect 112914 81030 112966 81082
rect 112978 81030 113030 81082
rect 113042 81030 113094 81082
rect 113106 81030 113158 81082
rect 113170 81030 113222 81082
rect 4874 80486 4926 80538
rect 4938 80486 4990 80538
rect 5002 80486 5054 80538
rect 5066 80486 5118 80538
rect 5130 80486 5182 80538
rect 113650 80486 113702 80538
rect 113714 80486 113766 80538
rect 113778 80486 113830 80538
rect 113842 80486 113894 80538
rect 113906 80486 113958 80538
rect 4214 79942 4266 79994
rect 4278 79942 4330 79994
rect 4342 79942 4394 79994
rect 4406 79942 4458 79994
rect 4470 79942 4522 79994
rect 112914 79942 112966 79994
rect 112978 79942 113030 79994
rect 113042 79942 113094 79994
rect 113106 79942 113158 79994
rect 113170 79942 113222 79994
rect 4874 79398 4926 79450
rect 4938 79398 4990 79450
rect 5002 79398 5054 79450
rect 5066 79398 5118 79450
rect 5130 79398 5182 79450
rect 113650 79398 113702 79450
rect 113714 79398 113766 79450
rect 113778 79398 113830 79450
rect 113842 79398 113894 79450
rect 113906 79398 113958 79450
rect 4214 78854 4266 78906
rect 4278 78854 4330 78906
rect 4342 78854 4394 78906
rect 4406 78854 4458 78906
rect 4470 78854 4522 78906
rect 112914 78854 112966 78906
rect 112978 78854 113030 78906
rect 113042 78854 113094 78906
rect 113106 78854 113158 78906
rect 113170 78854 113222 78906
rect 4874 78310 4926 78362
rect 4938 78310 4990 78362
rect 5002 78310 5054 78362
rect 5066 78310 5118 78362
rect 5130 78310 5182 78362
rect 113650 78310 113702 78362
rect 113714 78310 113766 78362
rect 113778 78310 113830 78362
rect 113842 78310 113894 78362
rect 113906 78310 113958 78362
rect 4214 77766 4266 77818
rect 4278 77766 4330 77818
rect 4342 77766 4394 77818
rect 4406 77766 4458 77818
rect 4470 77766 4522 77818
rect 112914 77766 112966 77818
rect 112978 77766 113030 77818
rect 113042 77766 113094 77818
rect 113106 77766 113158 77818
rect 113170 77766 113222 77818
rect 4874 77222 4926 77274
rect 4938 77222 4990 77274
rect 5002 77222 5054 77274
rect 5066 77222 5118 77274
rect 5130 77222 5182 77274
rect 113650 77222 113702 77274
rect 113714 77222 113766 77274
rect 113778 77222 113830 77274
rect 113842 77222 113894 77274
rect 113906 77222 113958 77274
rect 4214 76678 4266 76730
rect 4278 76678 4330 76730
rect 4342 76678 4394 76730
rect 4406 76678 4458 76730
rect 4470 76678 4522 76730
rect 112914 76678 112966 76730
rect 112978 76678 113030 76730
rect 113042 76678 113094 76730
rect 113106 76678 113158 76730
rect 113170 76678 113222 76730
rect 4874 76134 4926 76186
rect 4938 76134 4990 76186
rect 5002 76134 5054 76186
rect 5066 76134 5118 76186
rect 5130 76134 5182 76186
rect 113650 76134 113702 76186
rect 113714 76134 113766 76186
rect 113778 76134 113830 76186
rect 113842 76134 113894 76186
rect 113906 76134 113958 76186
rect 4214 75590 4266 75642
rect 4278 75590 4330 75642
rect 4342 75590 4394 75642
rect 4406 75590 4458 75642
rect 4470 75590 4522 75642
rect 112914 75590 112966 75642
rect 112978 75590 113030 75642
rect 113042 75590 113094 75642
rect 113106 75590 113158 75642
rect 113170 75590 113222 75642
rect 4874 75046 4926 75098
rect 4938 75046 4990 75098
rect 5002 75046 5054 75098
rect 5066 75046 5118 75098
rect 5130 75046 5182 75098
rect 113650 75046 113702 75098
rect 113714 75046 113766 75098
rect 113778 75046 113830 75098
rect 113842 75046 113894 75098
rect 113906 75046 113958 75098
rect 4214 74502 4266 74554
rect 4278 74502 4330 74554
rect 4342 74502 4394 74554
rect 4406 74502 4458 74554
rect 4470 74502 4522 74554
rect 112914 74502 112966 74554
rect 112978 74502 113030 74554
rect 113042 74502 113094 74554
rect 113106 74502 113158 74554
rect 113170 74502 113222 74554
rect 4874 73958 4926 74010
rect 4938 73958 4990 74010
rect 5002 73958 5054 74010
rect 5066 73958 5118 74010
rect 5130 73958 5182 74010
rect 113650 73958 113702 74010
rect 113714 73958 113766 74010
rect 113778 73958 113830 74010
rect 113842 73958 113894 74010
rect 113906 73958 113958 74010
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 112914 73414 112966 73466
rect 112978 73414 113030 73466
rect 113042 73414 113094 73466
rect 113106 73414 113158 73466
rect 113170 73414 113222 73466
rect 4874 72870 4926 72922
rect 4938 72870 4990 72922
rect 5002 72870 5054 72922
rect 5066 72870 5118 72922
rect 5130 72870 5182 72922
rect 113650 72870 113702 72922
rect 113714 72870 113766 72922
rect 113778 72870 113830 72922
rect 113842 72870 113894 72922
rect 113906 72870 113958 72922
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 112914 72326 112966 72378
rect 112978 72326 113030 72378
rect 113042 72326 113094 72378
rect 113106 72326 113158 72378
rect 113170 72326 113222 72378
rect 4874 71782 4926 71834
rect 4938 71782 4990 71834
rect 5002 71782 5054 71834
rect 5066 71782 5118 71834
rect 5130 71782 5182 71834
rect 113650 71782 113702 71834
rect 113714 71782 113766 71834
rect 113778 71782 113830 71834
rect 113842 71782 113894 71834
rect 113906 71782 113958 71834
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 112914 71238 112966 71290
rect 112978 71238 113030 71290
rect 113042 71238 113094 71290
rect 113106 71238 113158 71290
rect 113170 71238 113222 71290
rect 4874 70694 4926 70746
rect 4938 70694 4990 70746
rect 5002 70694 5054 70746
rect 5066 70694 5118 70746
rect 5130 70694 5182 70746
rect 113650 70694 113702 70746
rect 113714 70694 113766 70746
rect 113778 70694 113830 70746
rect 113842 70694 113894 70746
rect 113906 70694 113958 70746
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 112914 70150 112966 70202
rect 112978 70150 113030 70202
rect 113042 70150 113094 70202
rect 113106 70150 113158 70202
rect 113170 70150 113222 70202
rect 4874 69606 4926 69658
rect 4938 69606 4990 69658
rect 5002 69606 5054 69658
rect 5066 69606 5118 69658
rect 5130 69606 5182 69658
rect 113650 69606 113702 69658
rect 113714 69606 113766 69658
rect 113778 69606 113830 69658
rect 113842 69606 113894 69658
rect 113906 69606 113958 69658
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 112914 69062 112966 69114
rect 112978 69062 113030 69114
rect 113042 69062 113094 69114
rect 113106 69062 113158 69114
rect 113170 69062 113222 69114
rect 4874 68518 4926 68570
rect 4938 68518 4990 68570
rect 5002 68518 5054 68570
rect 5066 68518 5118 68570
rect 5130 68518 5182 68570
rect 113650 68518 113702 68570
rect 113714 68518 113766 68570
rect 113778 68518 113830 68570
rect 113842 68518 113894 68570
rect 113906 68518 113958 68570
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 112914 67974 112966 68026
rect 112978 67974 113030 68026
rect 113042 67974 113094 68026
rect 113106 67974 113158 68026
rect 113170 67974 113222 68026
rect 4874 67430 4926 67482
rect 4938 67430 4990 67482
rect 5002 67430 5054 67482
rect 5066 67430 5118 67482
rect 5130 67430 5182 67482
rect 113650 67430 113702 67482
rect 113714 67430 113766 67482
rect 113778 67430 113830 67482
rect 113842 67430 113894 67482
rect 113906 67430 113958 67482
rect 108396 67371 108448 67380
rect 108396 67337 108405 67371
rect 108405 67337 108439 67371
rect 108439 67337 108448 67371
rect 108396 67328 108448 67337
rect 109684 67192 109736 67244
rect 109960 66988 110012 67040
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 112914 66886 112966 66938
rect 112978 66886 113030 66938
rect 113042 66886 113094 66938
rect 113106 66886 113158 66938
rect 113170 66886 113222 66938
rect 4874 66342 4926 66394
rect 4938 66342 4990 66394
rect 5002 66342 5054 66394
rect 5066 66342 5118 66394
rect 5130 66342 5182 66394
rect 113650 66342 113702 66394
rect 113714 66342 113766 66394
rect 113778 66342 113830 66394
rect 113842 66342 113894 66394
rect 113906 66342 113958 66394
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 112914 65798 112966 65850
rect 112978 65798 113030 65850
rect 113042 65798 113094 65850
rect 113106 65798 113158 65850
rect 113170 65798 113222 65850
rect 4874 65254 4926 65306
rect 4938 65254 4990 65306
rect 5002 65254 5054 65306
rect 5066 65254 5118 65306
rect 5130 65254 5182 65306
rect 113650 65254 113702 65306
rect 113714 65254 113766 65306
rect 113778 65254 113830 65306
rect 113842 65254 113894 65306
rect 113906 65254 113958 65306
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 112914 64710 112966 64762
rect 112978 64710 113030 64762
rect 113042 64710 113094 64762
rect 113106 64710 113158 64762
rect 113170 64710 113222 64762
rect 4874 64166 4926 64218
rect 4938 64166 4990 64218
rect 5002 64166 5054 64218
rect 5066 64166 5118 64218
rect 5130 64166 5182 64218
rect 113650 64166 113702 64218
rect 113714 64166 113766 64218
rect 113778 64166 113830 64218
rect 113842 64166 113894 64218
rect 113906 64166 113958 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 112914 63622 112966 63674
rect 112978 63622 113030 63674
rect 113042 63622 113094 63674
rect 113106 63622 113158 63674
rect 113170 63622 113222 63674
rect 4874 63078 4926 63130
rect 4938 63078 4990 63130
rect 5002 63078 5054 63130
rect 5066 63078 5118 63130
rect 5130 63078 5182 63130
rect 113650 63078 113702 63130
rect 113714 63078 113766 63130
rect 113778 63078 113830 63130
rect 113842 63078 113894 63130
rect 113906 63078 113958 63130
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 112914 62534 112966 62586
rect 112978 62534 113030 62586
rect 113042 62534 113094 62586
rect 113106 62534 113158 62586
rect 113170 62534 113222 62586
rect 4874 61990 4926 62042
rect 4938 61990 4990 62042
rect 5002 61990 5054 62042
rect 5066 61990 5118 62042
rect 5130 61990 5182 62042
rect 113650 61990 113702 62042
rect 113714 61990 113766 62042
rect 113778 61990 113830 62042
rect 113842 61990 113894 62042
rect 113906 61990 113958 62042
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 112914 61446 112966 61498
rect 112978 61446 113030 61498
rect 113042 61446 113094 61498
rect 113106 61446 113158 61498
rect 113170 61446 113222 61498
rect 4874 60902 4926 60954
rect 4938 60902 4990 60954
rect 5002 60902 5054 60954
rect 5066 60902 5118 60954
rect 5130 60902 5182 60954
rect 113650 60902 113702 60954
rect 113714 60902 113766 60954
rect 113778 60902 113830 60954
rect 113842 60902 113894 60954
rect 113906 60902 113958 60954
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 112914 60358 112966 60410
rect 112978 60358 113030 60410
rect 113042 60358 113094 60410
rect 113106 60358 113158 60410
rect 113170 60358 113222 60410
rect 4874 59814 4926 59866
rect 4938 59814 4990 59866
rect 5002 59814 5054 59866
rect 5066 59814 5118 59866
rect 5130 59814 5182 59866
rect 113650 59814 113702 59866
rect 113714 59814 113766 59866
rect 113778 59814 113830 59866
rect 113842 59814 113894 59866
rect 113906 59814 113958 59866
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 112914 59270 112966 59322
rect 112978 59270 113030 59322
rect 113042 59270 113094 59322
rect 113106 59270 113158 59322
rect 113170 59270 113222 59322
rect 4874 58726 4926 58778
rect 4938 58726 4990 58778
rect 5002 58726 5054 58778
rect 5066 58726 5118 58778
rect 5130 58726 5182 58778
rect 113650 58726 113702 58778
rect 113714 58726 113766 58778
rect 113778 58726 113830 58778
rect 113842 58726 113894 58778
rect 113906 58726 113958 58778
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 112914 58182 112966 58234
rect 112978 58182 113030 58234
rect 113042 58182 113094 58234
rect 113106 58182 113158 58234
rect 113170 58182 113222 58234
rect 109960 57919 110012 57928
rect 109960 57885 109969 57919
rect 109969 57885 110003 57919
rect 110003 57885 110012 57919
rect 109960 57876 110012 57885
rect 108672 57808 108724 57860
rect 109684 57783 109736 57792
rect 109684 57749 109693 57783
rect 109693 57749 109727 57783
rect 109727 57749 109736 57783
rect 109684 57740 109736 57749
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 113650 57638 113702 57690
rect 113714 57638 113766 57690
rect 113778 57638 113830 57690
rect 113842 57638 113894 57690
rect 113906 57638 113958 57690
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 112914 57094 112966 57146
rect 112978 57094 113030 57146
rect 113042 57094 113094 57146
rect 113106 57094 113158 57146
rect 113170 57094 113222 57146
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 113650 56550 113702 56602
rect 113714 56550 113766 56602
rect 113778 56550 113830 56602
rect 113842 56550 113894 56602
rect 113906 56550 113958 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 112914 56006 112966 56058
rect 112978 56006 113030 56058
rect 113042 56006 113094 56058
rect 113106 56006 113158 56058
rect 113170 56006 113222 56058
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 113650 55462 113702 55514
rect 113714 55462 113766 55514
rect 113778 55462 113830 55514
rect 113842 55462 113894 55514
rect 113906 55462 113958 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 112914 54918 112966 54970
rect 112978 54918 113030 54970
rect 113042 54918 113094 54970
rect 113106 54918 113158 54970
rect 113170 54918 113222 54970
rect 108580 54859 108632 54868
rect 108580 54825 108589 54859
rect 108589 54825 108623 54859
rect 108623 54825 108632 54859
rect 108580 54816 108632 54825
rect 108580 54612 108632 54664
rect 109132 54544 109184 54596
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 113650 54374 113702 54426
rect 113714 54374 113766 54426
rect 113778 54374 113830 54426
rect 113842 54374 113894 54426
rect 113906 54374 113958 54426
rect 108304 54315 108356 54324
rect 108304 54281 108313 54315
rect 108313 54281 108347 54315
rect 108347 54281 108356 54315
rect 108304 54272 108356 54281
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 112914 53830 112966 53882
rect 112978 53830 113030 53882
rect 113042 53830 113094 53882
rect 113106 53830 113158 53882
rect 113170 53830 113222 53882
rect 108304 53567 108356 53576
rect 108304 53533 108313 53567
rect 108313 53533 108347 53567
rect 108347 53533 108356 53567
rect 108304 53524 108356 53533
rect 109040 53388 109092 53440
rect 109960 53388 110012 53440
rect 110696 53388 110748 53440
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 113650 53286 113702 53338
rect 113714 53286 113766 53338
rect 113778 53286 113830 53338
rect 113842 53286 113894 53338
rect 113906 53286 113958 53338
rect 109040 53227 109092 53236
rect 109040 53193 109049 53227
rect 109049 53193 109083 53227
rect 109083 53193 109092 53227
rect 109040 53184 109092 53193
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 112914 52742 112966 52794
rect 112978 52742 113030 52794
rect 113042 52742 113094 52794
rect 113106 52742 113158 52794
rect 113170 52742 113222 52794
rect 109040 52504 109092 52556
rect 110696 52436 110748 52488
rect 108580 52411 108632 52420
rect 108580 52377 108589 52411
rect 108589 52377 108623 52411
rect 108623 52377 108632 52411
rect 108580 52368 108632 52377
rect 109132 52368 109184 52420
rect 109408 52300 109460 52352
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 113650 52198 113702 52250
rect 113714 52198 113766 52250
rect 113778 52198 113830 52250
rect 113842 52198 113894 52250
rect 113906 52198 113958 52250
rect 108304 52139 108356 52148
rect 108304 52105 108313 52139
rect 108313 52105 108347 52139
rect 108347 52105 108356 52139
rect 108304 52096 108356 52105
rect 106924 52028 106976 52080
rect 109408 51960 109460 52012
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 112914 51654 112966 51706
rect 112978 51654 113030 51706
rect 113042 51654 113094 51706
rect 113106 51654 113158 51706
rect 113170 51654 113222 51706
rect 108304 51391 108356 51400
rect 108304 51357 108313 51391
rect 108313 51357 108347 51391
rect 108347 51357 108356 51391
rect 108304 51348 108356 51357
rect 109592 51255 109644 51264
rect 109592 51221 109601 51255
rect 109601 51221 109635 51255
rect 109635 51221 109644 51255
rect 109592 51212 109644 51221
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 113650 51110 113702 51162
rect 113714 51110 113766 51162
rect 113778 51110 113830 51162
rect 113842 51110 113894 51162
rect 113906 51110 113958 51162
rect 109592 50940 109644 50992
rect 108672 50872 108724 50924
rect 108948 50711 109000 50720
rect 108948 50677 108957 50711
rect 108957 50677 108991 50711
rect 108991 50677 109000 50711
rect 108948 50668 109000 50677
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 112914 50566 112966 50618
rect 112978 50566 113030 50618
rect 113042 50566 113094 50618
rect 113106 50566 113158 50618
rect 113170 50566 113222 50618
rect 108672 50507 108724 50516
rect 108672 50473 108681 50507
rect 108681 50473 108715 50507
rect 108715 50473 108724 50507
rect 108672 50464 108724 50473
rect 108672 50260 108724 50312
rect 109132 50192 109184 50244
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 113650 50022 113702 50074
rect 113714 50022 113766 50074
rect 113778 50022 113830 50074
rect 113842 50022 113894 50074
rect 113906 50022 113958 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 112914 49478 112966 49530
rect 112978 49478 113030 49530
rect 113042 49478 113094 49530
rect 113106 49478 113158 49530
rect 113170 49478 113222 49530
rect 108580 49376 108632 49428
rect 108672 49351 108724 49360
rect 108672 49317 108681 49351
rect 108681 49317 108715 49351
rect 108715 49317 108724 49351
rect 108672 49308 108724 49317
rect 109500 49308 109552 49360
rect 108304 49215 108356 49224
rect 108304 49181 108313 49215
rect 108313 49181 108347 49215
rect 108347 49181 108356 49215
rect 108304 49172 108356 49181
rect 109040 49104 109092 49156
rect 109408 49147 109460 49156
rect 109408 49113 109417 49147
rect 109417 49113 109451 49147
rect 109451 49113 109460 49147
rect 109408 49104 109460 49113
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 113650 48934 113702 48986
rect 113714 48934 113766 48986
rect 113778 48934 113830 48986
rect 113842 48934 113894 48986
rect 113906 48934 113958 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 112914 48390 112966 48442
rect 112978 48390 113030 48442
rect 113042 48390 113094 48442
rect 113106 48390 113158 48442
rect 113170 48390 113222 48442
rect 109592 48152 109644 48204
rect 110328 48195 110380 48204
rect 110328 48161 110337 48195
rect 110337 48161 110371 48195
rect 110371 48161 110380 48195
rect 110328 48152 110380 48161
rect 108948 48084 109000 48136
rect 110052 48059 110104 48068
rect 110052 48025 110061 48059
rect 110061 48025 110095 48059
rect 110095 48025 110104 48059
rect 110052 48016 110104 48025
rect 108580 47991 108632 48000
rect 108580 47957 108589 47991
rect 108589 47957 108623 47991
rect 108623 47957 108632 47991
rect 108580 47948 108632 47957
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 113650 47846 113702 47898
rect 113714 47846 113766 47898
rect 113778 47846 113830 47898
rect 113842 47846 113894 47898
rect 113906 47846 113958 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 112914 47302 112966 47354
rect 112978 47302 113030 47354
rect 113042 47302 113094 47354
rect 113106 47302 113158 47354
rect 113170 47302 113222 47354
rect 108764 47200 108816 47252
rect 110512 47200 110564 47252
rect 110420 47107 110472 47116
rect 110420 47073 110429 47107
rect 110429 47073 110463 47107
rect 110463 47073 110472 47107
rect 110420 47064 110472 47073
rect 109132 46928 109184 46980
rect 110144 46971 110196 46980
rect 110144 46937 110153 46971
rect 110153 46937 110187 46971
rect 110187 46937 110196 46971
rect 110144 46928 110196 46937
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 113650 46758 113702 46810
rect 113714 46758 113766 46810
rect 113778 46758 113830 46810
rect 113842 46758 113894 46810
rect 113906 46758 113958 46810
rect 108580 46520 108632 46572
rect 109684 46359 109736 46368
rect 109684 46325 109693 46359
rect 109693 46325 109727 46359
rect 109727 46325 109736 46359
rect 109684 46316 109736 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 112914 46214 112966 46266
rect 112978 46214 113030 46266
rect 113042 46214 113094 46266
rect 113106 46214 113158 46266
rect 113170 46214 113222 46266
rect 110328 46112 110380 46164
rect 108304 45951 108356 45960
rect 108304 45917 108313 45951
rect 108313 45917 108347 45951
rect 108347 45917 108356 45951
rect 108304 45908 108356 45917
rect 109040 45908 109092 45960
rect 110420 45840 110472 45892
rect 108488 45772 108540 45824
rect 109224 45772 109276 45824
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 113650 45670 113702 45722
rect 113714 45670 113766 45722
rect 113778 45670 113830 45722
rect 113842 45670 113894 45722
rect 113906 45670 113958 45722
rect 108304 45611 108356 45620
rect 108304 45577 108313 45611
rect 108313 45577 108347 45611
rect 108347 45577 108356 45611
rect 108304 45568 108356 45577
rect 109316 45500 109368 45552
rect 109408 45543 109460 45552
rect 109408 45509 109417 45543
rect 109417 45509 109451 45543
rect 109451 45509 109460 45543
rect 109408 45500 109460 45509
rect 109500 45500 109552 45552
rect 108580 45432 108632 45484
rect 109592 45432 109644 45484
rect 109684 45432 109736 45484
rect 110052 45364 110104 45416
rect 109132 45228 109184 45280
rect 109592 45228 109644 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 112914 45126 112966 45178
rect 112978 45126 113030 45178
rect 113042 45126 113094 45178
rect 113106 45126 113158 45178
rect 113170 45126 113222 45178
rect 109316 45024 109368 45076
rect 109500 44820 109552 44872
rect 109592 44863 109644 44872
rect 109592 44829 109601 44863
rect 109601 44829 109635 44863
rect 109635 44829 109644 44863
rect 109592 44820 109644 44829
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 113650 44582 113702 44634
rect 113714 44582 113766 44634
rect 113778 44582 113830 44634
rect 113842 44582 113894 44634
rect 113906 44582 113958 44634
rect 1308 44344 1360 44396
rect 108304 44387 108356 44396
rect 108304 44353 108313 44387
rect 108313 44353 108347 44387
rect 108347 44353 108356 44387
rect 108304 44344 108356 44353
rect 108856 44208 108908 44260
rect 9680 44140 9732 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 112914 44038 112966 44090
rect 112978 44038 113030 44090
rect 113042 44038 113094 44090
rect 113106 44038 113158 44090
rect 113170 44038 113222 44090
rect 108304 43936 108356 43988
rect 110144 43936 110196 43988
rect 110236 43979 110288 43988
rect 110236 43945 110245 43979
rect 110245 43945 110279 43979
rect 110279 43945 110288 43979
rect 110236 43936 110288 43945
rect 110420 43979 110472 43988
rect 110420 43945 110429 43979
rect 110429 43945 110463 43979
rect 110463 43945 110472 43979
rect 110420 43936 110472 43945
rect 109684 43800 109736 43852
rect 108304 43775 108356 43784
rect 108304 43741 108313 43775
rect 108313 43741 108347 43775
rect 108347 43741 108356 43775
rect 108304 43732 108356 43741
rect 109776 43775 109828 43784
rect 109776 43741 109785 43775
rect 109785 43741 109819 43775
rect 109819 43741 109828 43775
rect 109776 43732 109828 43741
rect 108672 43664 108724 43716
rect 109408 43664 109460 43716
rect 109868 43596 109920 43648
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 113650 43494 113702 43546
rect 113714 43494 113766 43546
rect 113778 43494 113830 43546
rect 113842 43494 113894 43546
rect 113906 43494 113958 43546
rect 110236 43392 110288 43444
rect 109132 43324 109184 43376
rect 1308 43256 1360 43308
rect 109224 43256 109276 43308
rect 109592 43299 109644 43308
rect 109592 43265 109601 43299
rect 109601 43265 109635 43299
rect 109635 43265 109644 43299
rect 109592 43256 109644 43265
rect 110144 43256 110196 43308
rect 9680 43120 9732 43172
rect 109960 43120 110012 43172
rect 109592 43052 109644 43104
rect 110144 43095 110196 43104
rect 110144 43061 110153 43095
rect 110153 43061 110187 43095
rect 110187 43061 110196 43095
rect 110144 43052 110196 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 112914 42950 112966 43002
rect 112978 42950 113030 43002
rect 113042 42950 113094 43002
rect 113106 42950 113158 43002
rect 113170 42950 113222 43002
rect 108304 42848 108356 42900
rect 109868 42891 109920 42900
rect 109868 42857 109877 42891
rect 109877 42857 109911 42891
rect 109911 42857 109920 42891
rect 109868 42848 109920 42857
rect 109500 42687 109552 42696
rect 109500 42653 109509 42687
rect 109509 42653 109543 42687
rect 109543 42653 109552 42687
rect 109500 42644 109552 42653
rect 110144 42644 110196 42696
rect 109592 42576 109644 42628
rect 109868 42576 109920 42628
rect 108488 42551 108540 42560
rect 108488 42517 108497 42551
rect 108497 42517 108531 42551
rect 108531 42517 108540 42551
rect 108488 42508 108540 42517
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 113650 42406 113702 42458
rect 113714 42406 113766 42458
rect 113778 42406 113830 42458
rect 113842 42406 113894 42458
rect 113906 42406 113958 42458
rect 108580 42236 108632 42288
rect 110328 42211 110380 42220
rect 110328 42177 110337 42211
rect 110337 42177 110371 42211
rect 110371 42177 110380 42211
rect 110328 42168 110380 42177
rect 110052 42143 110104 42152
rect 110052 42109 110061 42143
rect 110061 42109 110095 42143
rect 110095 42109 110104 42143
rect 110052 42100 110104 42109
rect 109500 41964 109552 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 112914 41862 112966 41914
rect 112978 41862 113030 41914
rect 113042 41862 113094 41914
rect 113106 41862 113158 41914
rect 113170 41862 113222 41914
rect 108304 41760 108356 41812
rect 109776 41760 109828 41812
rect 108948 41624 109000 41676
rect 108304 41599 108356 41608
rect 108304 41565 108313 41599
rect 108313 41565 108347 41599
rect 108347 41565 108356 41599
rect 108304 41556 108356 41565
rect 110512 41624 110564 41676
rect 109592 41488 109644 41540
rect 110236 41556 110288 41608
rect 110604 41488 110656 41540
rect 108396 41463 108448 41472
rect 108396 41429 108405 41463
rect 108405 41429 108439 41463
rect 108439 41429 108448 41463
rect 108396 41420 108448 41429
rect 110788 41463 110840 41472
rect 110788 41429 110797 41463
rect 110797 41429 110831 41463
rect 110831 41429 110840 41463
rect 110788 41420 110840 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 113650 41318 113702 41370
rect 113714 41318 113766 41370
rect 113778 41318 113830 41370
rect 113842 41318 113894 41370
rect 113906 41318 113958 41370
rect 1308 41080 1360 41132
rect 108764 41080 108816 41132
rect 108948 41080 109000 41132
rect 109684 41080 109736 41132
rect 109868 41080 109920 41132
rect 110236 41080 110288 41132
rect 110604 41123 110656 41132
rect 110604 41089 110613 41123
rect 110613 41089 110647 41123
rect 110647 41089 110656 41123
rect 110604 41080 110656 41089
rect 110880 41123 110932 41132
rect 110880 41089 110889 41123
rect 110889 41089 110923 41123
rect 110923 41089 110932 41123
rect 110880 41080 110932 41089
rect 9680 40944 9732 40996
rect 108948 40944 109000 40996
rect 110328 40944 110380 40996
rect 110236 40876 110288 40928
rect 110512 40876 110564 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 112914 40774 112966 40826
rect 112978 40774 113030 40826
rect 113042 40774 113094 40826
rect 113106 40774 113158 40826
rect 113170 40774 113222 40826
rect 110052 40672 110104 40724
rect 110328 40715 110380 40724
rect 110328 40681 110337 40715
rect 110337 40681 110371 40715
rect 110371 40681 110380 40715
rect 110328 40672 110380 40681
rect 109684 40604 109736 40656
rect 110604 40604 110656 40656
rect 108948 40536 109000 40588
rect 1308 40468 1360 40520
rect 109868 40468 109920 40520
rect 9680 40400 9732 40452
rect 108580 40443 108632 40452
rect 108580 40409 108589 40443
rect 108589 40409 108623 40443
rect 108623 40409 108632 40443
rect 108580 40400 108632 40409
rect 108856 40400 108908 40452
rect 113456 40468 113508 40520
rect 110144 40332 110196 40384
rect 110604 40332 110656 40384
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 113650 40230 113702 40282
rect 113714 40230 113766 40282
rect 113778 40230 113830 40282
rect 113842 40230 113894 40282
rect 113906 40230 113958 40282
rect 110144 40128 110196 40180
rect 110420 40171 110472 40180
rect 110420 40137 110429 40171
rect 110429 40137 110463 40171
rect 110463 40137 110472 40171
rect 110420 40128 110472 40137
rect 110788 40128 110840 40180
rect 109500 40035 109552 40044
rect 109500 40001 109509 40035
rect 109509 40001 109543 40035
rect 109543 40001 109552 40035
rect 109500 39992 109552 40001
rect 109592 40035 109644 40044
rect 109592 40001 109601 40035
rect 109601 40001 109635 40035
rect 109635 40001 109644 40035
rect 109592 39992 109644 40001
rect 109684 40035 109736 40044
rect 109684 40001 109693 40035
rect 109693 40001 109727 40035
rect 109727 40001 109736 40035
rect 109684 39992 109736 40001
rect 109960 39992 110012 40044
rect 110512 40060 110564 40112
rect 110880 40103 110932 40112
rect 110880 40069 110889 40103
rect 110889 40069 110923 40103
rect 110923 40069 110932 40103
rect 110880 40060 110932 40069
rect 110420 39924 110472 39976
rect 111340 39992 111392 40044
rect 110144 39788 110196 39840
rect 111156 39788 111208 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 112914 39686 112966 39738
rect 112978 39686 113030 39738
rect 113042 39686 113094 39738
rect 113106 39686 113158 39738
rect 113170 39686 113222 39738
rect 109776 39584 109828 39636
rect 110236 39584 110288 39636
rect 110696 39627 110748 39636
rect 110696 39593 110705 39627
rect 110705 39593 110739 39627
rect 110739 39593 110748 39627
rect 110696 39584 110748 39593
rect 110420 39448 110472 39500
rect 106924 39312 106976 39364
rect 108212 39244 108264 39296
rect 108672 39312 108724 39364
rect 109684 39312 109736 39364
rect 110236 39312 110288 39364
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 113650 39142 113702 39194
rect 113714 39142 113766 39194
rect 113778 39142 113830 39194
rect 113842 39142 113894 39194
rect 113906 39142 113958 39194
rect 109500 39083 109552 39092
rect 109500 39049 109509 39083
rect 109509 39049 109543 39083
rect 109543 39049 109552 39083
rect 109500 39040 109552 39049
rect 109592 39040 109644 39092
rect 109776 38972 109828 39024
rect 110328 39083 110380 39092
rect 110328 39049 110337 39083
rect 110337 39049 110371 39083
rect 110371 39049 110380 39083
rect 110328 39040 110380 39049
rect 110512 39040 110564 39092
rect 109960 38947 110012 38956
rect 109960 38913 109969 38947
rect 109969 38913 110003 38947
rect 110003 38913 110012 38947
rect 109960 38904 110012 38913
rect 109592 38768 109644 38820
rect 111340 38904 111392 38956
rect 110144 38743 110196 38752
rect 110144 38709 110153 38743
rect 110153 38709 110187 38743
rect 110187 38709 110196 38743
rect 110144 38700 110196 38709
rect 110972 38700 111024 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 112914 38598 112966 38650
rect 112978 38598 113030 38650
rect 113042 38598 113094 38650
rect 113106 38598 113158 38650
rect 113170 38598 113222 38650
rect 110880 38496 110932 38548
rect 108948 38428 109000 38480
rect 1216 38292 1268 38344
rect 111892 38335 111944 38344
rect 111892 38301 111901 38335
rect 111901 38301 111935 38335
rect 111935 38301 111944 38335
rect 111892 38292 111944 38301
rect 112352 38292 112404 38344
rect 9680 38224 9732 38276
rect 108488 38224 108540 38276
rect 110052 38267 110104 38276
rect 110052 38233 110061 38267
rect 110061 38233 110095 38267
rect 110095 38233 110104 38267
rect 110052 38224 110104 38233
rect 108672 38156 108724 38208
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 113650 38054 113702 38106
rect 113714 38054 113766 38106
rect 113778 38054 113830 38106
rect 113842 38054 113894 38106
rect 113906 38054 113958 38106
rect 108580 37952 108632 38004
rect 109868 37952 109920 38004
rect 109316 37927 109368 37936
rect 109316 37893 109343 37927
rect 109343 37893 109368 37927
rect 109316 37884 109368 37893
rect 109408 37884 109460 37936
rect 110144 37884 110196 37936
rect 1308 37816 1360 37868
rect 110604 37816 110656 37868
rect 112812 37816 112864 37868
rect 113456 37859 113508 37868
rect 113456 37825 113465 37859
rect 113465 37825 113499 37859
rect 113499 37825 113508 37859
rect 113456 37816 113508 37825
rect 114560 37859 114612 37868
rect 114560 37825 114569 37859
rect 114569 37825 114603 37859
rect 114603 37825 114612 37859
rect 114560 37816 114612 37825
rect 110328 37748 110380 37800
rect 110788 37791 110840 37800
rect 110788 37757 110797 37791
rect 110797 37757 110831 37791
rect 110831 37757 110840 37791
rect 110788 37748 110840 37757
rect 111892 37748 111944 37800
rect 9496 37680 9548 37732
rect 108764 37680 108816 37732
rect 111064 37723 111116 37732
rect 111064 37689 111073 37723
rect 111073 37689 111107 37723
rect 111107 37689 111116 37723
rect 111064 37680 111116 37689
rect 112352 37791 112404 37800
rect 112352 37757 112361 37791
rect 112361 37757 112395 37791
rect 112395 37757 112404 37791
rect 112352 37748 112404 37757
rect 113824 37791 113876 37800
rect 113824 37757 113833 37791
rect 113833 37757 113867 37791
rect 113867 37757 113876 37791
rect 113824 37748 113876 37757
rect 109960 37612 110012 37664
rect 110512 37612 110564 37664
rect 111248 37612 111300 37664
rect 112444 37612 112496 37664
rect 114100 37655 114152 37664
rect 114100 37621 114109 37655
rect 114109 37621 114143 37655
rect 114143 37621 114152 37655
rect 114100 37612 114152 37621
rect 114468 37655 114520 37664
rect 114468 37621 114477 37655
rect 114477 37621 114511 37655
rect 114511 37621 114520 37655
rect 114468 37612 114520 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 112914 37510 112966 37562
rect 112978 37510 113030 37562
rect 113042 37510 113094 37562
rect 113106 37510 113158 37562
rect 113170 37510 113222 37562
rect 108488 37408 108540 37460
rect 108856 37408 108908 37460
rect 110052 37408 110104 37460
rect 110788 37408 110840 37460
rect 113548 37408 113600 37460
rect 111248 37383 111300 37392
rect 111248 37349 111257 37383
rect 111257 37349 111291 37383
rect 111291 37349 111300 37383
rect 111248 37340 111300 37349
rect 112812 37383 112864 37392
rect 112812 37349 112821 37383
rect 112821 37349 112855 37383
rect 112855 37349 112864 37383
rect 112812 37340 112864 37349
rect 107016 37272 107068 37324
rect 109408 37204 109460 37256
rect 110144 37204 110196 37256
rect 113180 37204 113232 37256
rect 113456 37340 113508 37392
rect 113824 37272 113876 37324
rect 116400 37315 116452 37324
rect 116400 37281 116409 37315
rect 116409 37281 116443 37315
rect 116443 37281 116452 37315
rect 116400 37272 116452 37281
rect 109960 37136 110012 37188
rect 111708 37136 111760 37188
rect 114008 37204 114060 37256
rect 114284 37247 114336 37256
rect 114284 37213 114293 37247
rect 114293 37213 114327 37247
rect 114327 37213 114336 37247
rect 114284 37204 114336 37213
rect 114376 37247 114428 37256
rect 114376 37213 114385 37247
rect 114385 37213 114419 37247
rect 114419 37213 114428 37247
rect 114376 37204 114428 37213
rect 114192 37136 114244 37188
rect 115020 37204 115072 37256
rect 116308 37204 116360 37256
rect 114560 37136 114612 37188
rect 108856 37068 108908 37120
rect 112444 37111 112496 37120
rect 112444 37077 112453 37111
rect 112453 37077 112487 37111
rect 112487 37077 112496 37111
rect 112444 37068 112496 37077
rect 112536 37111 112588 37120
rect 112536 37077 112545 37111
rect 112545 37077 112579 37111
rect 112579 37077 112588 37111
rect 112536 37068 112588 37077
rect 114836 37179 114888 37188
rect 114836 37145 114845 37179
rect 114845 37145 114879 37179
rect 114879 37145 114888 37179
rect 114836 37136 114888 37145
rect 116216 37111 116268 37120
rect 116216 37077 116225 37111
rect 116225 37077 116259 37111
rect 116259 37077 116268 37111
rect 116216 37068 116268 37077
rect 116492 37068 116544 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 113650 36966 113702 37018
rect 113714 36966 113766 37018
rect 113778 36966 113830 37018
rect 113842 36966 113894 37018
rect 113906 36966 113958 37018
rect 108396 36796 108448 36848
rect 110420 36864 110472 36916
rect 112444 36864 112496 36916
rect 114652 36864 114704 36916
rect 114836 36864 114888 36916
rect 111064 36796 111116 36848
rect 112812 36796 112864 36848
rect 111892 36728 111944 36780
rect 109776 36703 109828 36712
rect 109776 36669 109785 36703
rect 109785 36669 109819 36703
rect 109819 36669 109828 36703
rect 109776 36660 109828 36669
rect 110788 36703 110840 36712
rect 110788 36669 110797 36703
rect 110797 36669 110831 36703
rect 110831 36669 110840 36703
rect 110788 36660 110840 36669
rect 111156 36660 111208 36712
rect 113180 36728 113232 36780
rect 113364 36728 113416 36780
rect 114100 36796 114152 36848
rect 114468 36796 114520 36848
rect 115112 36839 115164 36848
rect 115112 36805 115121 36839
rect 115121 36805 115155 36839
rect 115155 36805 115164 36839
rect 115112 36796 115164 36805
rect 113916 36771 113968 36780
rect 113916 36737 113925 36771
rect 113925 36737 113959 36771
rect 113959 36737 113968 36771
rect 113916 36728 113968 36737
rect 114008 36771 114060 36780
rect 114008 36737 114017 36771
rect 114017 36737 114051 36771
rect 114051 36737 114060 36771
rect 114008 36728 114060 36737
rect 114284 36771 114336 36780
rect 114284 36737 114293 36771
rect 114293 36737 114327 36771
rect 114327 36737 114336 36771
rect 114284 36728 114336 36737
rect 114376 36771 114428 36780
rect 114376 36737 114385 36771
rect 114385 36737 114419 36771
rect 114419 36737 114428 36771
rect 114376 36728 114428 36737
rect 114652 36771 114704 36780
rect 114652 36737 114661 36771
rect 114661 36737 114695 36771
rect 114695 36737 114704 36771
rect 114652 36728 114704 36737
rect 114928 36771 114980 36780
rect 114928 36737 114937 36771
rect 114937 36737 114971 36771
rect 114971 36737 114980 36771
rect 114928 36728 114980 36737
rect 115020 36771 115072 36780
rect 115020 36737 115029 36771
rect 115029 36737 115063 36771
rect 115063 36737 115072 36771
rect 115020 36728 115072 36737
rect 116124 36864 116176 36916
rect 116216 36907 116268 36916
rect 116216 36873 116225 36907
rect 116225 36873 116259 36907
rect 116259 36873 116268 36907
rect 116216 36864 116268 36873
rect 115572 36796 115624 36848
rect 116400 36796 116452 36848
rect 115848 36771 115900 36780
rect 115848 36737 115882 36771
rect 115882 36737 115900 36771
rect 115848 36728 115900 36737
rect 116124 36728 116176 36780
rect 108304 36567 108356 36576
rect 108304 36533 108313 36567
rect 108313 36533 108347 36567
rect 108347 36533 108356 36567
rect 108304 36524 108356 36533
rect 110696 36567 110748 36576
rect 110696 36533 110705 36567
rect 110705 36533 110739 36567
rect 110739 36533 110748 36567
rect 110696 36524 110748 36533
rect 110880 36567 110932 36576
rect 110880 36533 110889 36567
rect 110889 36533 110923 36567
rect 110923 36533 110932 36567
rect 110880 36524 110932 36533
rect 112168 36524 112220 36576
rect 113364 36592 113416 36644
rect 116492 36771 116544 36780
rect 116492 36737 116501 36771
rect 116501 36737 116535 36771
rect 116535 36737 116544 36771
rect 116492 36728 116544 36737
rect 116952 36771 117004 36780
rect 116952 36737 116961 36771
rect 116961 36737 116995 36771
rect 116995 36737 117004 36771
rect 116952 36728 117004 36737
rect 117136 36660 117188 36712
rect 113916 36524 113968 36576
rect 115204 36524 115256 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 112914 36422 112966 36474
rect 112978 36422 113030 36474
rect 113042 36422 113094 36474
rect 113106 36422 113158 36474
rect 113170 36422 113222 36474
rect 109408 36320 109460 36372
rect 109684 36320 109736 36372
rect 110788 36363 110840 36372
rect 110788 36329 110797 36363
rect 110797 36329 110831 36363
rect 110831 36329 110840 36363
rect 110788 36320 110840 36329
rect 112536 36320 112588 36372
rect 112352 36252 112404 36304
rect 113364 36320 113416 36372
rect 115020 36320 115072 36372
rect 115572 36363 115624 36372
rect 115572 36329 115581 36363
rect 115581 36329 115615 36363
rect 115615 36329 115624 36363
rect 115572 36320 115624 36329
rect 116952 36363 117004 36372
rect 116952 36329 116961 36363
rect 116961 36329 116995 36363
rect 116995 36329 117004 36363
rect 116952 36320 117004 36329
rect 113548 36252 113600 36304
rect 114376 36252 114428 36304
rect 114928 36252 114980 36304
rect 115388 36252 115440 36304
rect 110972 36227 111024 36236
rect 110972 36193 110981 36227
rect 110981 36193 111015 36227
rect 111015 36193 111024 36227
rect 110972 36184 111024 36193
rect 107108 36116 107160 36168
rect 110236 36116 110288 36168
rect 112352 36159 112404 36168
rect 112352 36125 112360 36159
rect 112360 36125 112394 36159
rect 112394 36125 112404 36159
rect 112352 36116 112404 36125
rect 112444 36159 112496 36168
rect 112444 36125 112453 36159
rect 112453 36125 112487 36159
rect 112487 36125 112496 36159
rect 112444 36116 112496 36125
rect 112536 36159 112588 36168
rect 112536 36125 112545 36159
rect 112545 36125 112579 36159
rect 112579 36125 112588 36159
rect 112536 36116 112588 36125
rect 109040 36048 109092 36100
rect 109868 36048 109920 36100
rect 112076 36091 112128 36100
rect 112076 36057 112085 36091
rect 112085 36057 112119 36091
rect 112119 36057 112128 36091
rect 112076 36048 112128 36057
rect 112168 36091 112220 36100
rect 112168 36057 112177 36091
rect 112177 36057 112211 36091
rect 112211 36057 112220 36091
rect 112168 36048 112220 36057
rect 112812 36116 112864 36168
rect 113088 36116 113140 36168
rect 113272 36116 113324 36168
rect 114100 36184 114152 36236
rect 113824 36159 113876 36168
rect 113824 36125 113833 36159
rect 113833 36125 113867 36159
rect 113867 36125 113876 36159
rect 113824 36116 113876 36125
rect 114008 36159 114060 36168
rect 114008 36125 114017 36159
rect 114017 36125 114051 36159
rect 114051 36125 114060 36159
rect 114008 36116 114060 36125
rect 114468 36048 114520 36100
rect 109224 35980 109276 36032
rect 113272 35980 113324 36032
rect 113824 35980 113876 36032
rect 115204 36184 115256 36236
rect 115204 36048 115256 36100
rect 115756 36116 115808 36168
rect 116124 36184 116176 36236
rect 117412 36184 117464 36236
rect 115480 36048 115532 36100
rect 116860 36159 116912 36168
rect 116860 36125 116869 36159
rect 116869 36125 116903 36159
rect 116903 36125 116912 36159
rect 116860 36116 116912 36125
rect 116952 36159 117004 36168
rect 116952 36125 116961 36159
rect 116961 36125 116995 36159
rect 116995 36125 117004 36159
rect 116952 36116 117004 36125
rect 117136 36159 117188 36168
rect 117136 36125 117145 36159
rect 117145 36125 117179 36159
rect 117179 36125 117188 36159
rect 117136 36116 117188 36125
rect 116492 36048 116544 36100
rect 114836 36023 114888 36032
rect 114836 35989 114845 36023
rect 114845 35989 114879 36023
rect 114879 35989 114888 36023
rect 114836 35980 114888 35989
rect 114928 36023 114980 36032
rect 114928 35989 114937 36023
rect 114937 35989 114971 36023
rect 114971 35989 114980 36023
rect 114928 35980 114980 35989
rect 115296 35980 115348 36032
rect 117320 35980 117372 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 113650 35878 113702 35930
rect 113714 35878 113766 35930
rect 113778 35878 113830 35930
rect 113842 35878 113894 35930
rect 113906 35878 113958 35930
rect 108764 35819 108816 35828
rect 108764 35785 108773 35819
rect 108773 35785 108807 35819
rect 108807 35785 108816 35819
rect 108764 35776 108816 35785
rect 9496 35708 9548 35760
rect 108948 35776 109000 35828
rect 109040 35751 109092 35760
rect 109040 35717 109065 35751
rect 109065 35717 109092 35751
rect 109316 35819 109368 35828
rect 109316 35785 109325 35819
rect 109325 35785 109359 35819
rect 109359 35785 109368 35819
rect 109316 35776 109368 35785
rect 111892 35819 111944 35828
rect 111892 35785 111901 35819
rect 111901 35785 111935 35819
rect 111935 35785 111944 35819
rect 111892 35776 111944 35785
rect 113364 35819 113416 35828
rect 113364 35785 113373 35819
rect 113373 35785 113407 35819
rect 113407 35785 113416 35819
rect 113364 35776 113416 35785
rect 114008 35776 114060 35828
rect 114836 35776 114888 35828
rect 116952 35819 117004 35828
rect 116952 35785 116961 35819
rect 116961 35785 116995 35819
rect 116995 35785 117004 35819
rect 116952 35776 117004 35785
rect 109040 35708 109092 35717
rect 109776 35708 109828 35760
rect 1308 35640 1360 35692
rect 108396 35504 108448 35556
rect 109592 35640 109644 35692
rect 110420 35683 110472 35692
rect 110420 35649 110429 35683
rect 110429 35649 110463 35683
rect 110463 35649 110472 35683
rect 110420 35640 110472 35649
rect 111708 35708 111760 35760
rect 114284 35708 114336 35760
rect 117412 35819 117464 35828
rect 117412 35785 117421 35819
rect 117421 35785 117455 35819
rect 117455 35785 117464 35819
rect 117412 35776 117464 35785
rect 110604 35640 110656 35692
rect 112536 35640 112588 35692
rect 112812 35640 112864 35692
rect 113088 35683 113140 35692
rect 113088 35649 113097 35683
rect 113097 35649 113131 35683
rect 113131 35649 113140 35683
rect 113088 35640 113140 35649
rect 113548 35683 113600 35692
rect 113548 35649 113557 35683
rect 113557 35649 113591 35683
rect 113591 35649 113600 35683
rect 113548 35640 113600 35649
rect 109592 35504 109644 35556
rect 110972 35572 111024 35624
rect 111616 35615 111668 35624
rect 111616 35581 111625 35615
rect 111625 35581 111659 35615
rect 111659 35581 111668 35615
rect 111616 35572 111668 35581
rect 113456 35572 113508 35624
rect 114192 35572 114244 35624
rect 112536 35504 112588 35556
rect 114376 35683 114428 35692
rect 114376 35649 114385 35683
rect 114385 35649 114419 35683
rect 114419 35649 114428 35683
rect 114376 35640 114428 35649
rect 115204 35683 115256 35692
rect 115204 35649 115213 35683
rect 115213 35649 115247 35683
rect 115247 35649 115256 35683
rect 115204 35640 115256 35649
rect 115296 35683 115348 35692
rect 115296 35649 115305 35683
rect 115305 35649 115339 35683
rect 115339 35649 115348 35683
rect 115296 35640 115348 35649
rect 115480 35683 115532 35692
rect 115480 35649 115489 35683
rect 115489 35649 115523 35683
rect 115523 35649 115532 35683
rect 115480 35640 115532 35649
rect 114468 35615 114520 35624
rect 114468 35581 114477 35615
rect 114477 35581 114511 35615
rect 114511 35581 114520 35615
rect 114468 35572 114520 35581
rect 115940 35572 115992 35624
rect 116032 35572 116084 35624
rect 116584 35683 116636 35692
rect 116584 35649 116593 35683
rect 116593 35649 116627 35683
rect 116627 35649 116636 35683
rect 116584 35640 116636 35649
rect 117044 35640 117096 35692
rect 115572 35504 115624 35556
rect 117872 35615 117924 35624
rect 117872 35581 117881 35615
rect 117881 35581 117915 35615
rect 117915 35581 117924 35615
rect 118240 35683 118292 35692
rect 118240 35649 118249 35683
rect 118249 35649 118283 35683
rect 118283 35649 118292 35683
rect 118240 35640 118292 35649
rect 117872 35572 117924 35581
rect 109040 35479 109092 35488
rect 109040 35445 109049 35479
rect 109049 35445 109083 35479
rect 109083 35445 109092 35479
rect 109040 35436 109092 35445
rect 109500 35436 109552 35488
rect 115204 35436 115256 35488
rect 118240 35436 118292 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 112914 35334 112966 35386
rect 112978 35334 113030 35386
rect 113042 35334 113094 35386
rect 113106 35334 113158 35386
rect 113170 35334 113222 35386
rect 109040 35232 109092 35284
rect 111616 35275 111668 35284
rect 111616 35241 111625 35275
rect 111625 35241 111659 35275
rect 111659 35241 111668 35275
rect 111616 35232 111668 35241
rect 112444 35232 112496 35284
rect 112536 35232 112588 35284
rect 112996 35232 113048 35284
rect 110880 35164 110932 35216
rect 112076 35164 112128 35216
rect 113272 35164 113324 35216
rect 113640 35164 113692 35216
rect 114100 35275 114152 35284
rect 114100 35241 114109 35275
rect 114109 35241 114143 35275
rect 114143 35241 114152 35275
rect 114100 35232 114152 35241
rect 115112 35232 115164 35284
rect 116584 35232 116636 35284
rect 117320 35275 117372 35284
rect 117320 35241 117329 35275
rect 117329 35241 117363 35275
rect 117363 35241 117372 35275
rect 117320 35232 117372 35241
rect 118240 35232 118292 35284
rect 111248 35096 111300 35148
rect 108764 35028 108816 35080
rect 110604 35028 110656 35080
rect 111984 34960 112036 35012
rect 112904 35071 112956 35080
rect 112904 35037 112913 35071
rect 112913 35037 112947 35071
rect 112947 35037 112956 35071
rect 112904 35028 112956 35037
rect 113456 35096 113508 35148
rect 114192 35096 114244 35148
rect 114560 35164 114612 35216
rect 113364 35028 113416 35080
rect 112812 34960 112864 35012
rect 113640 35071 113692 35080
rect 113640 35037 113649 35071
rect 113649 35037 113683 35071
rect 113683 35037 113692 35071
rect 113640 35028 113692 35037
rect 114652 35096 114704 35148
rect 114468 35071 114520 35080
rect 114468 35037 114477 35071
rect 114477 35037 114511 35071
rect 114511 35037 114520 35071
rect 114468 35028 114520 35037
rect 116124 35139 116176 35148
rect 116124 35105 116133 35139
rect 116133 35105 116167 35139
rect 116167 35105 116176 35139
rect 116124 35096 116176 35105
rect 117596 35139 117648 35148
rect 117596 35105 117605 35139
rect 117605 35105 117639 35139
rect 117639 35105 117648 35139
rect 117596 35096 117648 35105
rect 115204 35071 115256 35080
rect 115204 35037 115213 35071
rect 115213 35037 115247 35071
rect 115247 35037 115256 35071
rect 115204 35028 115256 35037
rect 115296 35071 115348 35080
rect 115296 35037 115305 35071
rect 115305 35037 115339 35071
rect 115339 35037 115348 35071
rect 115296 35028 115348 35037
rect 115480 35071 115532 35080
rect 115480 35037 115489 35071
rect 115489 35037 115523 35071
rect 115523 35037 115532 35071
rect 115480 35028 115532 35037
rect 116308 35028 116360 35080
rect 110604 34892 110656 34944
rect 111064 34892 111116 34944
rect 112996 34892 113048 34944
rect 116492 34960 116544 35012
rect 117136 34960 117188 35012
rect 117964 34960 118016 35012
rect 118148 35003 118200 35012
rect 118148 34969 118157 35003
rect 118157 34969 118191 35003
rect 118191 34969 118200 35003
rect 118148 34960 118200 34969
rect 118332 35003 118384 35012
rect 118332 34969 118341 35003
rect 118341 34969 118375 35003
rect 118375 34969 118384 35003
rect 118332 34960 118384 34969
rect 114008 34892 114060 34944
rect 114100 34892 114152 34944
rect 114376 34892 114428 34944
rect 114652 34892 114704 34944
rect 115296 34892 115348 34944
rect 117228 34892 117280 34944
rect 117872 34892 117924 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 113650 34790 113702 34842
rect 113714 34790 113766 34842
rect 113778 34790 113830 34842
rect 113842 34790 113894 34842
rect 113906 34790 113958 34842
rect 108488 34688 108540 34740
rect 109224 34731 109276 34740
rect 109224 34697 109233 34731
rect 109233 34697 109267 34731
rect 109267 34697 109276 34731
rect 109224 34688 109276 34697
rect 109408 34731 109460 34740
rect 109408 34697 109417 34731
rect 109417 34697 109451 34731
rect 109451 34697 109460 34731
rect 109408 34688 109460 34697
rect 108212 34620 108264 34672
rect 109960 34663 110012 34672
rect 109960 34629 109969 34663
rect 109969 34629 110003 34663
rect 110003 34629 110012 34663
rect 109960 34620 110012 34629
rect 110696 34663 110748 34672
rect 110696 34629 110705 34663
rect 110705 34629 110739 34663
rect 110739 34629 110748 34663
rect 110696 34620 110748 34629
rect 111064 34620 111116 34672
rect 111248 34688 111300 34740
rect 112076 34688 112128 34740
rect 108488 34595 108540 34604
rect 108488 34561 108497 34595
rect 108497 34561 108531 34595
rect 108531 34561 108540 34595
rect 108488 34552 108540 34561
rect 108580 34552 108632 34604
rect 108764 34552 108816 34604
rect 109040 34595 109092 34604
rect 109040 34561 109049 34595
rect 109049 34561 109083 34595
rect 109083 34561 109092 34595
rect 109040 34552 109092 34561
rect 110604 34552 110656 34604
rect 109960 34484 110012 34536
rect 110328 34527 110380 34536
rect 110328 34493 110337 34527
rect 110337 34493 110371 34527
rect 110371 34493 110380 34527
rect 110328 34484 110380 34493
rect 111340 34620 111392 34672
rect 111708 34552 111760 34604
rect 110512 34459 110564 34468
rect 110512 34425 110540 34459
rect 110540 34425 110564 34459
rect 110512 34416 110564 34425
rect 111892 34416 111944 34468
rect 114100 34731 114152 34740
rect 114100 34697 114109 34731
rect 114109 34697 114143 34731
rect 114143 34697 114152 34731
rect 114100 34688 114152 34697
rect 114468 34688 114520 34740
rect 116124 34688 116176 34740
rect 114100 34552 114152 34604
rect 114284 34552 114336 34604
rect 113548 34484 113600 34536
rect 114928 34620 114980 34672
rect 115480 34620 115532 34672
rect 115020 34595 115072 34604
rect 115020 34561 115029 34595
rect 115029 34561 115063 34595
rect 115063 34561 115072 34595
rect 115020 34552 115072 34561
rect 115664 34595 115716 34604
rect 115664 34561 115673 34595
rect 115673 34561 115707 34595
rect 115707 34561 115716 34595
rect 115664 34552 115716 34561
rect 117228 34595 117280 34604
rect 117228 34561 117237 34595
rect 117237 34561 117271 34595
rect 117271 34561 117280 34595
rect 117228 34552 117280 34561
rect 117504 34595 117556 34604
rect 117504 34561 117513 34595
rect 117513 34561 117547 34595
rect 117547 34561 117556 34595
rect 117504 34552 117556 34561
rect 117688 34595 117740 34604
rect 117688 34561 117697 34595
rect 117697 34561 117731 34595
rect 117731 34561 117740 34595
rect 117688 34552 117740 34561
rect 109868 34391 109920 34400
rect 109868 34357 109877 34391
rect 109877 34357 109911 34391
rect 109911 34357 109920 34391
rect 109868 34348 109920 34357
rect 110144 34348 110196 34400
rect 110788 34391 110840 34400
rect 110788 34357 110797 34391
rect 110797 34357 110831 34391
rect 110831 34357 110840 34391
rect 110788 34348 110840 34357
rect 110972 34391 111024 34400
rect 110972 34357 110981 34391
rect 110981 34357 111015 34391
rect 111015 34357 111024 34391
rect 110972 34348 111024 34357
rect 111616 34348 111668 34400
rect 114560 34416 114612 34468
rect 115112 34527 115164 34536
rect 115112 34493 115121 34527
rect 115121 34493 115155 34527
rect 115155 34493 115164 34527
rect 115112 34484 115164 34493
rect 115572 34527 115624 34536
rect 115572 34493 115581 34527
rect 115581 34493 115615 34527
rect 115615 34493 115624 34527
rect 115572 34484 115624 34493
rect 116032 34484 116084 34536
rect 117780 34484 117832 34536
rect 118332 34484 118384 34536
rect 113732 34348 113784 34400
rect 114192 34348 114244 34400
rect 117412 34459 117464 34468
rect 117412 34425 117421 34459
rect 117421 34425 117455 34459
rect 117455 34425 117464 34459
rect 117412 34416 117464 34425
rect 118148 34416 118200 34468
rect 117044 34391 117096 34400
rect 117044 34357 117053 34391
rect 117053 34357 117087 34391
rect 117087 34357 117096 34391
rect 117044 34348 117096 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 112914 34246 112966 34298
rect 112978 34246 113030 34298
rect 113042 34246 113094 34298
rect 113106 34246 113158 34298
rect 113170 34246 113222 34298
rect 108856 34187 108908 34196
rect 108856 34153 108865 34187
rect 108865 34153 108899 34187
rect 108899 34153 108908 34187
rect 108856 34144 108908 34153
rect 109592 34144 109644 34196
rect 110512 34144 110564 34196
rect 113456 34144 113508 34196
rect 110052 34076 110104 34128
rect 110972 34076 111024 34128
rect 112812 34076 112864 34128
rect 114008 34187 114060 34196
rect 114008 34153 114017 34187
rect 114017 34153 114051 34187
rect 114051 34153 114060 34187
rect 114008 34144 114060 34153
rect 114284 34144 114336 34196
rect 115020 34144 115072 34196
rect 116492 34144 116544 34196
rect 108488 33983 108540 33992
rect 108488 33949 108497 33983
rect 108497 33949 108531 33983
rect 108531 33949 108540 33983
rect 108488 33940 108540 33949
rect 108580 33940 108632 33992
rect 109040 33983 109092 33992
rect 109040 33949 109049 33983
rect 109049 33949 109083 33983
rect 109083 33949 109092 33983
rect 109040 33940 109092 33949
rect 110788 34008 110840 34060
rect 109868 33940 109920 33992
rect 110236 33983 110288 33992
rect 110236 33949 110245 33983
rect 110245 33949 110279 33983
rect 110279 33949 110288 33983
rect 110236 33940 110288 33949
rect 110420 33940 110472 33992
rect 108764 33872 108816 33924
rect 111340 33940 111392 33992
rect 111708 34008 111760 34060
rect 114192 33940 114244 33992
rect 117044 34076 117096 34128
rect 114928 33983 114980 33992
rect 114928 33949 114937 33983
rect 114937 33949 114971 33983
rect 114971 33949 114980 33983
rect 114928 33940 114980 33949
rect 116308 34008 116360 34060
rect 117412 34144 117464 34196
rect 117688 34144 117740 34196
rect 109224 33847 109276 33856
rect 109224 33813 109233 33847
rect 109233 33813 109267 33847
rect 109267 33813 109276 33847
rect 109224 33804 109276 33813
rect 111432 33872 111484 33924
rect 113732 33915 113784 33924
rect 113732 33881 113759 33915
rect 113759 33881 113784 33915
rect 113732 33872 113784 33881
rect 116032 33983 116084 33992
rect 116032 33949 116041 33983
rect 116041 33949 116075 33983
rect 116075 33949 116084 33983
rect 116032 33940 116084 33949
rect 116124 33983 116176 33992
rect 116124 33949 116133 33983
rect 116133 33949 116167 33983
rect 116167 33949 116176 33983
rect 116124 33940 116176 33949
rect 116492 33940 116544 33992
rect 117780 34008 117832 34060
rect 117964 33983 118016 33992
rect 117964 33949 117973 33983
rect 117973 33949 118007 33983
rect 118007 33949 118016 33983
rect 117964 33940 118016 33949
rect 110972 33847 111024 33856
rect 110972 33813 110981 33847
rect 110981 33813 111015 33847
rect 111015 33813 111024 33847
rect 110972 33804 111024 33813
rect 111616 33804 111668 33856
rect 111708 33847 111760 33856
rect 111708 33813 111717 33847
rect 111717 33813 111751 33847
rect 111751 33813 111760 33847
rect 111708 33804 111760 33813
rect 111800 33847 111852 33856
rect 111800 33813 111809 33847
rect 111809 33813 111843 33847
rect 111843 33813 111852 33847
rect 111800 33804 111852 33813
rect 114376 33804 114428 33856
rect 115572 33804 115624 33856
rect 117596 33872 117648 33924
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 113650 33702 113702 33754
rect 113714 33702 113766 33754
rect 113778 33702 113830 33754
rect 113842 33702 113894 33754
rect 113906 33702 113958 33754
rect 108488 33600 108540 33652
rect 109684 33600 109736 33652
rect 109224 33532 109276 33584
rect 108304 33507 108356 33516
rect 108304 33473 108313 33507
rect 108313 33473 108347 33507
rect 108347 33473 108356 33507
rect 108304 33464 108356 33473
rect 108672 33464 108724 33516
rect 109132 33507 109184 33516
rect 109132 33473 109141 33507
rect 109141 33473 109175 33507
rect 109175 33473 109184 33507
rect 109132 33464 109184 33473
rect 109776 33464 109828 33516
rect 110604 33396 110656 33448
rect 111340 33507 111392 33516
rect 111340 33473 111349 33507
rect 111349 33473 111383 33507
rect 111383 33473 111392 33507
rect 111340 33464 111392 33473
rect 111432 33507 111484 33516
rect 111432 33473 111441 33507
rect 111441 33473 111475 33507
rect 111475 33473 111484 33507
rect 111432 33464 111484 33473
rect 115112 33600 115164 33652
rect 115204 33600 115256 33652
rect 115572 33643 115624 33652
rect 115572 33609 115581 33643
rect 115581 33609 115615 33643
rect 115615 33609 115624 33643
rect 115572 33600 115624 33609
rect 116308 33600 116360 33652
rect 109592 33371 109644 33380
rect 109592 33337 109601 33371
rect 109601 33337 109635 33371
rect 109635 33337 109644 33371
rect 109592 33328 109644 33337
rect 111616 33439 111668 33448
rect 111616 33405 111625 33439
rect 111625 33405 111659 33439
rect 111659 33405 111668 33439
rect 111616 33396 111668 33405
rect 108948 33260 109000 33312
rect 109408 33303 109460 33312
rect 109408 33269 109417 33303
rect 109417 33269 109451 33303
rect 109451 33269 109460 33303
rect 109408 33260 109460 33269
rect 111800 33464 111852 33516
rect 111984 33507 112036 33516
rect 111984 33473 111993 33507
rect 111993 33473 112027 33507
rect 112027 33473 112036 33507
rect 111984 33464 112036 33473
rect 115756 33532 115808 33584
rect 116216 33532 116268 33584
rect 112628 33507 112680 33516
rect 112628 33473 112637 33507
rect 112637 33473 112671 33507
rect 112671 33473 112680 33507
rect 112628 33464 112680 33473
rect 112720 33464 112772 33516
rect 114560 33464 114612 33516
rect 114836 33507 114888 33516
rect 114836 33473 114845 33507
rect 114845 33473 114879 33507
rect 114879 33473 114888 33507
rect 114836 33464 114888 33473
rect 115664 33464 115716 33516
rect 117504 33600 117556 33652
rect 114008 33396 114060 33448
rect 116032 33396 116084 33448
rect 116124 33396 116176 33448
rect 115480 33328 115532 33380
rect 117136 33439 117188 33448
rect 117136 33405 117145 33439
rect 117145 33405 117179 33439
rect 117179 33405 117188 33439
rect 117136 33396 117188 33405
rect 117688 33396 117740 33448
rect 115388 33260 115440 33312
rect 116676 33328 116728 33380
rect 117964 33328 118016 33380
rect 116952 33260 117004 33312
rect 117780 33260 117832 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 112914 33158 112966 33210
rect 112978 33158 113030 33210
rect 113042 33158 113094 33210
rect 113106 33158 113158 33210
rect 113170 33158 113222 33210
rect 108856 33056 108908 33108
rect 109132 33056 109184 33108
rect 109684 33099 109736 33108
rect 109684 33065 109693 33099
rect 109693 33065 109727 33099
rect 109727 33065 109736 33099
rect 109684 33056 109736 33065
rect 110236 33056 110288 33108
rect 114560 33056 114612 33108
rect 115204 33099 115256 33108
rect 115204 33065 115213 33099
rect 115213 33065 115247 33099
rect 115247 33065 115256 33099
rect 115204 33056 115256 33065
rect 116032 33056 116084 33108
rect 116676 33099 116728 33108
rect 116676 33065 116685 33099
rect 116685 33065 116719 33099
rect 116719 33065 116728 33099
rect 116676 33056 116728 33065
rect 117596 33099 117648 33108
rect 117596 33065 117605 33099
rect 117605 33065 117639 33099
rect 117639 33065 117648 33099
rect 117596 33056 117648 33065
rect 117688 33099 117740 33108
rect 117688 33065 117697 33099
rect 117697 33065 117731 33099
rect 117731 33065 117740 33099
rect 117688 33056 117740 33065
rect 108304 32988 108356 33040
rect 110052 32988 110104 33040
rect 111984 32988 112036 33040
rect 108304 32895 108356 32904
rect 108304 32861 108313 32895
rect 108313 32861 108347 32895
rect 108347 32861 108356 32895
rect 108304 32852 108356 32861
rect 110972 32920 111024 32972
rect 111616 32920 111668 32972
rect 109224 32895 109276 32904
rect 109224 32861 109233 32895
rect 109233 32861 109267 32895
rect 109267 32861 109276 32895
rect 109224 32852 109276 32861
rect 111800 32852 111852 32904
rect 112720 32895 112772 32904
rect 112720 32861 112729 32895
rect 112729 32861 112763 32895
rect 112763 32861 112772 32895
rect 112720 32852 112772 32861
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 109776 32784 109828 32836
rect 112536 32784 112588 32836
rect 115020 32852 115072 32904
rect 115756 32920 115808 32972
rect 117136 32988 117188 33040
rect 118148 32963 118200 32972
rect 118148 32929 118157 32963
rect 118157 32929 118191 32963
rect 118191 32929 118200 32963
rect 118148 32920 118200 32929
rect 112996 32784 113048 32836
rect 115296 32784 115348 32836
rect 115848 32895 115900 32904
rect 115848 32861 115857 32895
rect 115857 32861 115891 32895
rect 115891 32861 115900 32895
rect 115848 32852 115900 32861
rect 115940 32895 115992 32904
rect 115940 32861 115949 32895
rect 115949 32861 115983 32895
rect 115983 32861 115992 32895
rect 115940 32852 115992 32861
rect 109408 32716 109460 32768
rect 109868 32716 109920 32768
rect 113180 32716 113232 32768
rect 114284 32716 114336 32768
rect 115480 32716 115532 32768
rect 115848 32716 115900 32768
rect 116216 32895 116268 32904
rect 116216 32861 116225 32895
rect 116225 32861 116259 32895
rect 116259 32861 116268 32895
rect 116216 32852 116268 32861
rect 116400 32852 116452 32904
rect 117688 32852 117740 32904
rect 117136 32759 117188 32768
rect 117136 32725 117145 32759
rect 117145 32725 117179 32759
rect 117179 32725 117188 32759
rect 117136 32716 117188 32725
rect 117228 32759 117280 32768
rect 117228 32725 117237 32759
rect 117237 32725 117271 32759
rect 117271 32725 117280 32759
rect 117228 32716 117280 32725
rect 113650 32614 113702 32666
rect 113714 32614 113766 32666
rect 113778 32614 113830 32666
rect 113842 32614 113894 32666
rect 113906 32614 113958 32666
rect 108396 32512 108448 32564
rect 108672 32555 108724 32564
rect 108672 32521 108681 32555
rect 108681 32521 108715 32555
rect 108715 32521 108724 32555
rect 108672 32512 108724 32521
rect 110144 32512 110196 32564
rect 112628 32512 112680 32564
rect 114468 32512 114520 32564
rect 115664 32555 115716 32564
rect 115664 32521 115673 32555
rect 115673 32521 115707 32555
rect 115707 32521 115716 32555
rect 115664 32512 115716 32521
rect 116124 32512 116176 32564
rect 116216 32512 116268 32564
rect 117596 32512 117648 32564
rect 117688 32555 117740 32564
rect 117688 32521 117697 32555
rect 117697 32521 117731 32555
rect 117731 32521 117740 32555
rect 117688 32512 117740 32521
rect 118148 32555 118200 32564
rect 118148 32521 118157 32555
rect 118157 32521 118191 32555
rect 118191 32521 118200 32555
rect 118148 32512 118200 32521
rect 108948 32419 109000 32428
rect 108948 32385 108957 32419
rect 108957 32385 108991 32419
rect 108991 32385 109000 32419
rect 108948 32376 109000 32385
rect 109500 32376 109552 32428
rect 110972 32419 111024 32428
rect 110972 32385 110981 32419
rect 110981 32385 111015 32419
rect 111015 32385 111024 32419
rect 110972 32376 111024 32385
rect 111432 32376 111484 32428
rect 109868 32308 109920 32360
rect 111340 32308 111392 32360
rect 108488 32215 108540 32224
rect 108488 32181 108497 32215
rect 108497 32181 108531 32215
rect 108531 32181 108540 32215
rect 108488 32172 108540 32181
rect 109408 32172 109460 32224
rect 110880 32172 110932 32224
rect 112168 32419 112220 32428
rect 112168 32385 112177 32419
rect 112177 32385 112211 32419
rect 112211 32385 112220 32419
rect 112168 32376 112220 32385
rect 112720 32419 112772 32428
rect 112076 32308 112128 32360
rect 112720 32385 112729 32419
rect 112729 32385 112763 32419
rect 112763 32385 112772 32419
rect 112720 32376 112772 32385
rect 112996 32376 113048 32428
rect 112444 32308 112496 32360
rect 114284 32419 114336 32428
rect 114284 32385 114296 32419
rect 114296 32385 114330 32419
rect 114330 32385 114336 32419
rect 114284 32376 114336 32385
rect 113456 32240 113508 32292
rect 111984 32172 112036 32224
rect 112260 32172 112312 32224
rect 112352 32172 112404 32224
rect 114192 32240 114244 32292
rect 115204 32308 115256 32360
rect 115388 32376 115440 32428
rect 115480 32308 115532 32360
rect 116308 32376 116360 32428
rect 115848 32308 115900 32360
rect 115940 32240 115992 32292
rect 116216 32308 116268 32360
rect 116768 32419 116820 32428
rect 116768 32385 116777 32419
rect 116777 32385 116811 32419
rect 116811 32385 116820 32419
rect 116768 32376 116820 32385
rect 116860 32419 116912 32428
rect 116860 32385 116869 32419
rect 116869 32385 116903 32419
rect 116903 32385 116912 32419
rect 116860 32376 116912 32385
rect 116952 32376 117004 32428
rect 116584 32308 116636 32360
rect 117320 32376 117372 32428
rect 117504 32419 117556 32428
rect 117504 32385 117513 32419
rect 117513 32385 117547 32419
rect 117547 32385 117556 32419
rect 117504 32376 117556 32385
rect 117780 32419 117832 32428
rect 117780 32385 117789 32419
rect 117789 32385 117823 32419
rect 117823 32385 117832 32419
rect 117780 32376 117832 32385
rect 113916 32215 113968 32224
rect 113916 32181 113925 32215
rect 113925 32181 113959 32215
rect 113959 32181 113968 32215
rect 113916 32172 113968 32181
rect 114928 32215 114980 32224
rect 114928 32181 114937 32215
rect 114937 32181 114971 32215
rect 114971 32181 114980 32215
rect 114928 32172 114980 32181
rect 115112 32172 115164 32224
rect 116216 32172 116268 32224
rect 116308 32215 116360 32224
rect 116308 32181 116317 32215
rect 116317 32181 116351 32215
rect 116351 32181 116360 32215
rect 116308 32172 116360 32181
rect 117412 32240 117464 32292
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 112914 32070 112966 32122
rect 112978 32070 113030 32122
rect 113042 32070 113094 32122
rect 113106 32070 113158 32122
rect 113170 32070 113222 32122
rect 112076 31968 112128 32020
rect 115388 32011 115440 32020
rect 115388 31977 115397 32011
rect 115397 31977 115431 32011
rect 115431 31977 115440 32011
rect 115388 31968 115440 31977
rect 115480 32011 115532 32020
rect 115480 31977 115489 32011
rect 115489 31977 115523 32011
rect 115523 31977 115532 32011
rect 115480 31968 115532 31977
rect 108764 31832 108816 31884
rect 110328 31900 110380 31952
rect 110604 31900 110656 31952
rect 111708 31900 111760 31952
rect 113180 31900 113232 31952
rect 114100 31900 114152 31952
rect 109960 31832 110012 31884
rect 110880 31875 110932 31884
rect 110880 31841 110889 31875
rect 110889 31841 110923 31875
rect 110923 31841 110932 31875
rect 110880 31832 110932 31841
rect 111892 31832 111944 31884
rect 115204 31900 115256 31952
rect 116032 31968 116084 32020
rect 114468 31832 114520 31884
rect 108304 31807 108356 31816
rect 108304 31773 108313 31807
rect 108313 31773 108347 31807
rect 108347 31773 108356 31807
rect 108304 31764 108356 31773
rect 108488 31807 108540 31816
rect 108488 31773 108497 31807
rect 108497 31773 108531 31807
rect 108531 31773 108540 31807
rect 108488 31764 108540 31773
rect 108856 31807 108908 31816
rect 108856 31773 108865 31807
rect 108865 31773 108899 31807
rect 108899 31773 108908 31807
rect 108856 31764 108908 31773
rect 110420 31764 110472 31816
rect 111800 31807 111852 31816
rect 111800 31773 111809 31807
rect 111809 31773 111843 31807
rect 111843 31773 111852 31807
rect 111800 31764 111852 31773
rect 111432 31628 111484 31680
rect 111524 31628 111576 31680
rect 112352 31696 112404 31748
rect 113272 31807 113324 31816
rect 113272 31773 113281 31807
rect 113281 31773 113315 31807
rect 113315 31773 113324 31807
rect 113272 31764 113324 31773
rect 114008 31764 114060 31816
rect 114100 31807 114152 31816
rect 114100 31773 114109 31807
rect 114109 31773 114143 31807
rect 114143 31773 114152 31807
rect 114100 31764 114152 31773
rect 114928 31764 114980 31816
rect 117136 31968 117188 32020
rect 116860 31900 116912 31952
rect 117596 31900 117648 31952
rect 115940 31875 115992 31884
rect 115940 31841 115949 31875
rect 115949 31841 115983 31875
rect 115983 31841 115992 31875
rect 115940 31832 115992 31841
rect 116400 31832 116452 31884
rect 113456 31696 113508 31748
rect 113916 31696 113968 31748
rect 114284 31696 114336 31748
rect 115756 31764 115808 31816
rect 117320 31832 117372 31884
rect 116952 31764 117004 31816
rect 116216 31696 116268 31748
rect 117596 31807 117648 31816
rect 117596 31773 117605 31807
rect 117605 31773 117639 31807
rect 117639 31773 117648 31807
rect 117596 31764 117648 31773
rect 118516 31807 118568 31816
rect 118516 31773 118525 31807
rect 118525 31773 118559 31807
rect 118559 31773 118568 31807
rect 118516 31764 118568 31773
rect 117964 31696 118016 31748
rect 114376 31628 114428 31680
rect 115848 31628 115900 31680
rect 115940 31628 115992 31680
rect 116676 31628 116728 31680
rect 117228 31628 117280 31680
rect 118332 31671 118384 31680
rect 118332 31637 118341 31671
rect 118341 31637 118375 31671
rect 118375 31637 118384 31671
rect 118332 31628 118384 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 113650 31526 113702 31578
rect 113714 31526 113766 31578
rect 113778 31526 113830 31578
rect 113842 31526 113894 31578
rect 113906 31526 113958 31578
rect 110972 31424 111024 31476
rect 108856 31399 108908 31408
rect 108856 31365 108865 31399
rect 108865 31365 108899 31399
rect 108899 31365 108908 31399
rect 108856 31356 108908 31365
rect 110052 31356 110104 31408
rect 111892 31424 111944 31476
rect 112168 31424 112220 31476
rect 112444 31467 112496 31476
rect 112444 31433 112453 31467
rect 112453 31433 112487 31467
rect 112487 31433 112496 31467
rect 112444 31424 112496 31433
rect 114468 31467 114520 31476
rect 114468 31433 114477 31467
rect 114477 31433 114511 31467
rect 114511 31433 114520 31467
rect 114468 31424 114520 31433
rect 111800 31356 111852 31408
rect 113272 31356 113324 31408
rect 109592 31288 109644 31340
rect 108304 31152 108356 31204
rect 110512 31263 110564 31272
rect 110512 31229 110521 31263
rect 110521 31229 110555 31263
rect 110555 31229 110564 31263
rect 110512 31220 110564 31229
rect 110604 31152 110656 31204
rect 111892 31331 111944 31340
rect 111892 31297 111901 31331
rect 111901 31297 111935 31331
rect 111935 31297 111944 31331
rect 111892 31288 111944 31297
rect 111984 31288 112036 31340
rect 112260 31331 112312 31340
rect 112260 31297 112269 31331
rect 112269 31297 112303 31331
rect 112303 31297 112312 31331
rect 112260 31288 112312 31297
rect 112352 31220 112404 31272
rect 112536 31263 112588 31272
rect 112536 31229 112545 31263
rect 112545 31229 112579 31263
rect 112579 31229 112588 31263
rect 112536 31220 112588 31229
rect 112812 31288 112864 31340
rect 113456 31331 113508 31340
rect 113456 31297 113465 31331
rect 113465 31297 113499 31331
rect 113499 31297 113508 31331
rect 113456 31288 113508 31297
rect 113824 31331 113876 31340
rect 113824 31297 113833 31331
rect 113833 31297 113867 31331
rect 113867 31297 113876 31331
rect 113824 31288 113876 31297
rect 114100 31331 114152 31340
rect 114100 31297 114109 31331
rect 114109 31297 114143 31331
rect 114143 31297 114152 31331
rect 114100 31288 114152 31297
rect 114284 31288 114336 31340
rect 116124 31424 116176 31476
rect 116584 31467 116636 31476
rect 116584 31433 116593 31467
rect 116593 31433 116627 31467
rect 116627 31433 116636 31467
rect 116584 31424 116636 31433
rect 115112 31356 115164 31408
rect 117780 31424 117832 31476
rect 117964 31424 118016 31476
rect 116768 31356 116820 31408
rect 116952 31399 117004 31408
rect 116952 31365 116961 31399
rect 116961 31365 116995 31399
rect 116995 31365 117004 31399
rect 116952 31356 117004 31365
rect 114652 31288 114704 31340
rect 115940 31288 115992 31340
rect 116400 31331 116452 31340
rect 116400 31297 116409 31331
rect 116409 31297 116443 31331
rect 116443 31297 116452 31331
rect 116400 31288 116452 31297
rect 116492 31331 116544 31340
rect 116492 31297 116501 31331
rect 116501 31297 116535 31331
rect 116535 31297 116544 31331
rect 116492 31288 116544 31297
rect 116676 31331 116728 31340
rect 116676 31297 116685 31331
rect 116685 31297 116719 31331
rect 116719 31297 116728 31331
rect 116676 31288 116728 31297
rect 113364 31152 113416 31204
rect 114376 31152 114428 31204
rect 116584 31220 116636 31272
rect 117412 31331 117464 31340
rect 117412 31297 117421 31331
rect 117421 31297 117455 31331
rect 117455 31297 117464 31331
rect 117412 31288 117464 31297
rect 118516 31331 118568 31340
rect 118516 31297 118525 31331
rect 118525 31297 118559 31331
rect 118559 31297 118568 31331
rect 118516 31288 118568 31297
rect 108764 31127 108816 31136
rect 108764 31093 108773 31127
rect 108773 31093 108807 31127
rect 108807 31093 108816 31127
rect 108764 31084 108816 31093
rect 111340 31127 111392 31136
rect 111340 31093 111349 31127
rect 111349 31093 111383 31127
rect 111383 31093 111392 31127
rect 111340 31084 111392 31093
rect 111616 31084 111668 31136
rect 114192 31084 114244 31136
rect 114560 31127 114612 31136
rect 114560 31093 114569 31127
rect 114569 31093 114603 31127
rect 114603 31093 114612 31127
rect 114560 31084 114612 31093
rect 114836 31084 114888 31136
rect 117964 31152 118016 31204
rect 116308 31127 116360 31136
rect 116308 31093 116317 31127
rect 116317 31093 116351 31127
rect 116351 31093 116360 31127
rect 116308 31084 116360 31093
rect 117136 31084 117188 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 112914 30982 112966 31034
rect 112978 30982 113030 31034
rect 113042 30982 113094 31034
rect 113106 30982 113158 31034
rect 113170 30982 113222 31034
rect 109592 30880 109644 30932
rect 110512 30880 110564 30932
rect 111432 30923 111484 30932
rect 111432 30889 111441 30923
rect 111441 30889 111475 30923
rect 111475 30889 111484 30923
rect 111432 30880 111484 30889
rect 111708 30880 111760 30932
rect 114652 30880 114704 30932
rect 116032 30923 116084 30932
rect 116032 30889 116041 30923
rect 116041 30889 116075 30923
rect 116075 30889 116084 30923
rect 116032 30880 116084 30889
rect 110052 30855 110104 30864
rect 110052 30821 110061 30855
rect 110061 30821 110095 30855
rect 110095 30821 110104 30855
rect 110052 30812 110104 30821
rect 110880 30744 110932 30796
rect 111892 30744 111944 30796
rect 109224 30719 109276 30728
rect 109224 30685 109233 30719
rect 109233 30685 109267 30719
rect 109267 30685 109276 30719
rect 109224 30676 109276 30685
rect 109684 30719 109736 30728
rect 109684 30685 109693 30719
rect 109693 30685 109727 30719
rect 109727 30685 109736 30719
rect 109684 30676 109736 30685
rect 110328 30676 110380 30728
rect 110512 30676 110564 30728
rect 111340 30676 111392 30728
rect 111616 30719 111668 30728
rect 111616 30685 111625 30719
rect 111625 30685 111659 30719
rect 111659 30685 111668 30719
rect 111616 30676 111668 30685
rect 111892 30651 111944 30660
rect 111892 30617 111901 30651
rect 111901 30617 111935 30651
rect 111935 30617 111944 30651
rect 111892 30608 111944 30617
rect 115112 30812 115164 30864
rect 116584 30880 116636 30932
rect 117136 30923 117188 30932
rect 117136 30889 117145 30923
rect 117145 30889 117179 30923
rect 117179 30889 117188 30923
rect 117136 30880 117188 30889
rect 117320 30923 117372 30932
rect 117320 30889 117329 30923
rect 117329 30889 117363 30923
rect 117363 30889 117372 30923
rect 117320 30880 117372 30889
rect 113272 30744 113324 30796
rect 113088 30719 113140 30728
rect 113088 30685 113097 30719
rect 113097 30685 113131 30719
rect 113131 30685 113140 30719
rect 113088 30676 113140 30685
rect 113824 30676 113876 30728
rect 114284 30744 114336 30796
rect 114468 30744 114520 30796
rect 114928 30744 114980 30796
rect 115480 30744 115532 30796
rect 114652 30719 114704 30728
rect 114652 30685 114661 30719
rect 114661 30685 114695 30719
rect 114695 30685 114704 30719
rect 114652 30676 114704 30685
rect 113364 30608 113416 30660
rect 112076 30583 112128 30592
rect 112076 30549 112085 30583
rect 112085 30549 112119 30583
rect 112119 30549 112128 30583
rect 112076 30540 112128 30549
rect 113088 30540 113140 30592
rect 113548 30608 113600 30660
rect 114008 30540 114060 30592
rect 116032 30676 116084 30728
rect 116400 30812 116452 30864
rect 116860 30812 116912 30864
rect 116400 30676 116452 30728
rect 116952 30676 117004 30728
rect 117964 30719 118016 30728
rect 117964 30685 117973 30719
rect 117973 30685 118007 30719
rect 118007 30685 118016 30719
rect 117964 30676 118016 30685
rect 118332 30676 118384 30728
rect 115940 30608 115992 30660
rect 116492 30583 116544 30592
rect 116492 30549 116501 30583
rect 116501 30549 116535 30583
rect 116535 30549 116544 30583
rect 116492 30540 116544 30549
rect 116584 30540 116636 30592
rect 117136 30540 117188 30592
rect 117596 30583 117648 30592
rect 117596 30549 117605 30583
rect 117605 30549 117639 30583
rect 117639 30549 117648 30583
rect 117596 30540 117648 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 113650 30438 113702 30490
rect 113714 30438 113766 30490
rect 113778 30438 113830 30490
rect 113842 30438 113894 30490
rect 113906 30438 113958 30490
rect 109224 30379 109276 30388
rect 109224 30345 109233 30379
rect 109233 30345 109267 30379
rect 109267 30345 109276 30379
rect 109224 30336 109276 30345
rect 110880 30336 110932 30388
rect 109592 30268 109644 30320
rect 109776 30243 109828 30252
rect 109776 30209 109785 30243
rect 109785 30209 109819 30243
rect 109819 30209 109828 30243
rect 109776 30200 109828 30209
rect 109868 30200 109920 30252
rect 110420 30268 110472 30320
rect 110144 30243 110196 30252
rect 110144 30209 110153 30243
rect 110153 30209 110187 30243
rect 110187 30209 110196 30243
rect 110144 30200 110196 30209
rect 110604 30243 110656 30252
rect 110604 30209 110613 30243
rect 110613 30209 110647 30243
rect 110647 30209 110656 30243
rect 110604 30200 110656 30209
rect 110880 30243 110932 30252
rect 110880 30209 110889 30243
rect 110889 30209 110923 30243
rect 110923 30209 110932 30243
rect 110880 30200 110932 30209
rect 111248 30200 111300 30252
rect 111524 30336 111576 30388
rect 112076 30379 112128 30388
rect 112076 30345 112085 30379
rect 112085 30345 112119 30379
rect 112119 30345 112128 30379
rect 112076 30336 112128 30345
rect 113548 30336 113600 30388
rect 114928 30336 114980 30388
rect 111984 30243 112036 30252
rect 111984 30209 111993 30243
rect 111993 30209 112027 30243
rect 112027 30209 112036 30243
rect 111984 30200 112036 30209
rect 112076 30243 112128 30252
rect 112076 30209 112085 30243
rect 112085 30209 112119 30243
rect 112119 30209 112128 30243
rect 112536 30268 112588 30320
rect 114560 30268 114612 30320
rect 112076 30200 112128 30209
rect 112260 30243 112312 30252
rect 112260 30209 112269 30243
rect 112269 30209 112303 30243
rect 112303 30209 112312 30243
rect 112260 30200 112312 30209
rect 112812 30200 112864 30252
rect 113732 30243 113784 30252
rect 113732 30209 113741 30243
rect 113741 30209 113775 30243
rect 113775 30209 113784 30243
rect 113732 30200 113784 30209
rect 111892 30132 111944 30184
rect 114192 30175 114244 30184
rect 114192 30141 114201 30175
rect 114201 30141 114235 30175
rect 114235 30141 114244 30175
rect 114192 30132 114244 30141
rect 115020 30064 115072 30116
rect 116308 30268 116360 30320
rect 117136 30336 117188 30388
rect 117872 30336 117924 30388
rect 116860 30311 116912 30320
rect 116860 30277 116869 30311
rect 116869 30277 116903 30311
rect 116903 30277 116912 30311
rect 116860 30268 116912 30277
rect 116400 30200 116452 30252
rect 116492 30243 116544 30252
rect 116492 30209 116501 30243
rect 116501 30209 116535 30243
rect 116535 30209 116544 30243
rect 116492 30200 116544 30209
rect 116584 30200 116636 30252
rect 116952 30243 117004 30252
rect 116952 30209 116961 30243
rect 116961 30209 116995 30243
rect 116995 30209 117004 30243
rect 116952 30200 117004 30209
rect 117596 30268 117648 30320
rect 117228 30243 117280 30252
rect 117228 30209 117237 30243
rect 117237 30209 117271 30243
rect 117271 30209 117280 30243
rect 117228 30200 117280 30209
rect 117780 30200 117832 30252
rect 118516 30311 118568 30320
rect 118516 30277 118525 30311
rect 118525 30277 118559 30311
rect 118559 30277 118568 30311
rect 118516 30268 118568 30277
rect 116032 30132 116084 30184
rect 118056 30200 118108 30252
rect 111156 30039 111208 30048
rect 111156 30005 111165 30039
rect 111165 30005 111199 30039
rect 111199 30005 111208 30039
rect 111156 29996 111208 30005
rect 115388 30039 115440 30048
rect 115388 30005 115397 30039
rect 115397 30005 115431 30039
rect 115431 30005 115440 30039
rect 115388 29996 115440 30005
rect 116860 30064 116912 30116
rect 115756 29996 115808 30048
rect 115848 30039 115900 30048
rect 115848 30005 115857 30039
rect 115857 30005 115891 30039
rect 115891 30005 115900 30039
rect 115848 29996 115900 30005
rect 116124 30039 116176 30048
rect 116124 30005 116133 30039
rect 116133 30005 116167 30039
rect 116167 30005 116176 30039
rect 116124 29996 116176 30005
rect 116584 30039 116636 30048
rect 116584 30005 116593 30039
rect 116593 30005 116627 30039
rect 116627 30005 116636 30039
rect 116584 29996 116636 30005
rect 117412 29996 117464 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 112914 29894 112966 29946
rect 112978 29894 113030 29946
rect 113042 29894 113094 29946
rect 113106 29894 113158 29946
rect 113170 29894 113222 29946
rect 109684 29792 109736 29844
rect 109776 29792 109828 29844
rect 110144 29792 110196 29844
rect 110604 29792 110656 29844
rect 111156 29792 111208 29844
rect 110420 29724 110472 29776
rect 110972 29724 111024 29776
rect 111248 29767 111300 29776
rect 111248 29733 111257 29767
rect 111257 29733 111291 29767
rect 111291 29733 111300 29767
rect 111248 29724 111300 29733
rect 109868 29656 109920 29708
rect 110052 29656 110104 29708
rect 109592 29588 109644 29640
rect 109776 29631 109828 29640
rect 109776 29597 109785 29631
rect 109785 29597 109819 29631
rect 109819 29597 109828 29631
rect 109776 29588 109828 29597
rect 110144 29588 110196 29640
rect 110788 29631 110840 29640
rect 110788 29597 110797 29631
rect 110797 29597 110831 29631
rect 110831 29597 110840 29631
rect 110788 29588 110840 29597
rect 110972 29631 111024 29640
rect 110972 29597 110981 29631
rect 110981 29597 111015 29631
rect 111015 29597 111024 29631
rect 110972 29588 111024 29597
rect 111064 29631 111116 29640
rect 111064 29597 111073 29631
rect 111073 29597 111107 29631
rect 111107 29597 111116 29631
rect 111064 29588 111116 29597
rect 112076 29656 112128 29708
rect 114192 29792 114244 29844
rect 114100 29656 114152 29708
rect 111708 29631 111760 29640
rect 111708 29597 111717 29631
rect 111717 29597 111751 29631
rect 111751 29597 111760 29631
rect 111708 29588 111760 29597
rect 111892 29631 111944 29640
rect 111892 29597 111901 29631
rect 111901 29597 111935 29631
rect 111935 29597 111944 29631
rect 111892 29588 111944 29597
rect 112260 29520 112312 29572
rect 114928 29631 114980 29640
rect 114928 29597 114937 29631
rect 114937 29597 114971 29631
rect 114971 29597 114980 29631
rect 114928 29588 114980 29597
rect 115296 29588 115348 29640
rect 115388 29588 115440 29640
rect 115848 29631 115900 29640
rect 115848 29597 115857 29631
rect 115857 29597 115891 29631
rect 115891 29597 115900 29631
rect 115848 29588 115900 29597
rect 117780 29835 117832 29844
rect 117780 29801 117789 29835
rect 117789 29801 117823 29835
rect 117823 29801 117832 29835
rect 117780 29792 117832 29801
rect 117872 29792 117924 29844
rect 116492 29656 116544 29708
rect 116584 29631 116636 29640
rect 116584 29597 116593 29631
rect 116593 29597 116627 29631
rect 116627 29597 116636 29631
rect 116584 29588 116636 29597
rect 117504 29724 117556 29776
rect 118332 29724 118384 29776
rect 116768 29520 116820 29572
rect 117596 29588 117648 29640
rect 118056 29631 118108 29640
rect 118056 29597 118065 29631
rect 118065 29597 118099 29631
rect 118099 29597 118108 29631
rect 118056 29588 118108 29597
rect 118516 29631 118568 29640
rect 118516 29597 118525 29631
rect 118525 29597 118559 29631
rect 118559 29597 118568 29631
rect 118516 29588 118568 29597
rect 117780 29563 117832 29572
rect 117780 29529 117791 29563
rect 117791 29529 117832 29563
rect 117780 29520 117832 29529
rect 117964 29563 118016 29572
rect 117964 29529 117973 29563
rect 117973 29529 118007 29563
rect 118007 29529 118016 29563
rect 117964 29520 118016 29529
rect 110052 29495 110104 29504
rect 110052 29461 110061 29495
rect 110061 29461 110095 29495
rect 110095 29461 110104 29495
rect 110052 29452 110104 29461
rect 112812 29452 112864 29504
rect 114744 29452 114796 29504
rect 115112 29452 115164 29504
rect 115940 29452 115992 29504
rect 116860 29495 116912 29504
rect 116860 29461 116869 29495
rect 116869 29461 116903 29495
rect 116903 29461 116912 29495
rect 116860 29452 116912 29461
rect 117320 29495 117372 29504
rect 117320 29461 117329 29495
rect 117329 29461 117363 29495
rect 117363 29461 117372 29495
rect 117320 29452 117372 29461
rect 117504 29452 117556 29504
rect 117596 29495 117648 29504
rect 117596 29461 117605 29495
rect 117605 29461 117639 29495
rect 117639 29461 117648 29495
rect 117596 29452 117648 29461
rect 118148 29452 118200 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 113650 29350 113702 29402
rect 113714 29350 113766 29402
rect 113778 29350 113830 29402
rect 113842 29350 113894 29402
rect 113906 29350 113958 29402
rect 109592 29291 109644 29300
rect 109592 29257 109601 29291
rect 109601 29257 109635 29291
rect 109635 29257 109644 29291
rect 109592 29248 109644 29257
rect 109868 29248 109920 29300
rect 110144 29248 110196 29300
rect 110328 29248 110380 29300
rect 110788 29248 110840 29300
rect 113364 29248 113416 29300
rect 109776 29180 109828 29232
rect 109684 29044 109736 29096
rect 110144 29155 110196 29164
rect 110144 29121 110153 29155
rect 110153 29121 110187 29155
rect 110187 29121 110196 29155
rect 110144 29112 110196 29121
rect 110604 29112 110656 29164
rect 110420 29044 110472 29096
rect 111064 28976 111116 29028
rect 113456 29180 113508 29232
rect 116216 29248 116268 29300
rect 116952 29248 117004 29300
rect 117412 29291 117464 29300
rect 117412 29257 117421 29291
rect 117421 29257 117455 29291
rect 117455 29257 117464 29291
rect 117412 29248 117464 29257
rect 111340 29155 111392 29164
rect 111340 29121 111349 29155
rect 111349 29121 111383 29155
rect 111383 29121 111392 29155
rect 111340 29112 111392 29121
rect 111984 29044 112036 29096
rect 111800 28976 111852 29028
rect 113732 29155 113784 29164
rect 113732 29121 113741 29155
rect 113741 29121 113775 29155
rect 113775 29121 113784 29155
rect 113732 29112 113784 29121
rect 114192 29112 114244 29164
rect 114928 29155 114980 29164
rect 114928 29121 114937 29155
rect 114937 29121 114971 29155
rect 114971 29121 114980 29155
rect 114928 29112 114980 29121
rect 115112 29155 115164 29164
rect 115112 29121 115121 29155
rect 115121 29121 115155 29155
rect 115155 29121 115164 29155
rect 115112 29112 115164 29121
rect 114008 29044 114060 29096
rect 115112 28976 115164 29028
rect 115480 29155 115532 29164
rect 115480 29121 115489 29155
rect 115489 29121 115523 29155
rect 115523 29121 115532 29155
rect 115480 29112 115532 29121
rect 115940 29155 115992 29164
rect 115940 29121 115949 29155
rect 115949 29121 115983 29155
rect 115983 29121 115992 29155
rect 115940 29112 115992 29121
rect 116860 29180 116912 29232
rect 117596 29180 117648 29232
rect 110420 28951 110472 28960
rect 110420 28917 110429 28951
rect 110429 28917 110463 28951
rect 110463 28917 110472 28951
rect 110420 28908 110472 28917
rect 115480 28908 115532 28960
rect 116492 29155 116544 29164
rect 116492 29121 116501 29155
rect 116501 29121 116535 29155
rect 116535 29121 116544 29155
rect 116492 29112 116544 29121
rect 116768 29112 116820 29164
rect 117320 29112 117372 29164
rect 117412 29044 117464 29096
rect 117596 29044 117648 29096
rect 117688 28976 117740 29028
rect 118148 29019 118200 29028
rect 118148 28985 118157 29019
rect 118157 28985 118191 29019
rect 118191 28985 118200 29019
rect 118148 28976 118200 28985
rect 118516 29019 118568 29028
rect 118516 28985 118525 29019
rect 118525 28985 118559 29019
rect 118559 28985 118568 29019
rect 118516 28976 118568 28985
rect 116676 28908 116728 28960
rect 116860 28951 116912 28960
rect 116860 28917 116869 28951
rect 116869 28917 116903 28951
rect 116903 28917 116912 28951
rect 116860 28908 116912 28917
rect 116952 28908 117004 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 112914 28806 112966 28858
rect 112978 28806 113030 28858
rect 113042 28806 113094 28858
rect 113106 28806 113158 28858
rect 113170 28806 113222 28858
rect 110052 28704 110104 28756
rect 109776 28568 109828 28620
rect 109868 28543 109920 28552
rect 109868 28509 109877 28543
rect 109877 28509 109911 28543
rect 109911 28509 109920 28543
rect 109868 28500 109920 28509
rect 110144 28568 110196 28620
rect 111708 28704 111760 28756
rect 111984 28747 112036 28756
rect 111984 28713 111993 28747
rect 111993 28713 112027 28747
rect 112027 28713 112036 28747
rect 111984 28704 112036 28713
rect 112444 28704 112496 28756
rect 113456 28704 113508 28756
rect 113732 28704 113784 28756
rect 114100 28704 114152 28756
rect 114928 28704 114980 28756
rect 118056 28747 118108 28756
rect 118056 28713 118065 28747
rect 118065 28713 118099 28747
rect 118099 28713 118108 28747
rect 118056 28704 118108 28713
rect 110604 28636 110656 28688
rect 110236 28500 110288 28552
rect 112260 28500 112312 28552
rect 112444 28543 112496 28552
rect 112444 28509 112453 28543
rect 112453 28509 112487 28543
rect 112487 28509 112496 28543
rect 112444 28500 112496 28509
rect 115940 28636 115992 28688
rect 116124 28636 116176 28688
rect 110420 28432 110472 28484
rect 110788 28432 110840 28484
rect 112628 28364 112680 28416
rect 113548 28543 113600 28552
rect 113548 28509 113557 28543
rect 113557 28509 113591 28543
rect 113591 28509 113600 28543
rect 113548 28500 113600 28509
rect 114744 28611 114796 28620
rect 114744 28577 114753 28611
rect 114753 28577 114787 28611
rect 114787 28577 114796 28611
rect 114744 28568 114796 28577
rect 114836 28611 114888 28620
rect 114836 28577 114845 28611
rect 114845 28577 114879 28611
rect 114879 28577 114888 28611
rect 114836 28568 114888 28577
rect 115020 28568 115072 28620
rect 115480 28568 115532 28620
rect 114376 28543 114428 28552
rect 114376 28509 114385 28543
rect 114385 28509 114419 28543
rect 114419 28509 114428 28543
rect 114376 28500 114428 28509
rect 114468 28500 114520 28552
rect 113456 28475 113508 28484
rect 113456 28441 113465 28475
rect 113465 28441 113499 28475
rect 113499 28441 113508 28475
rect 115112 28543 115164 28552
rect 115112 28509 115121 28543
rect 115121 28509 115155 28543
rect 115155 28509 115164 28543
rect 115112 28500 115164 28509
rect 115296 28543 115348 28552
rect 115296 28509 115305 28543
rect 115305 28509 115339 28543
rect 115339 28509 115348 28543
rect 115296 28500 115348 28509
rect 116216 28543 116268 28552
rect 116216 28509 116225 28543
rect 116225 28509 116259 28543
rect 116259 28509 116268 28543
rect 116216 28500 116268 28509
rect 117136 28500 117188 28552
rect 117780 28500 117832 28552
rect 113456 28432 113508 28441
rect 113548 28364 113600 28416
rect 117044 28432 117096 28484
rect 118240 28543 118292 28552
rect 118240 28509 118249 28543
rect 118249 28509 118283 28543
rect 118283 28509 118292 28543
rect 118240 28500 118292 28509
rect 118608 28500 118660 28552
rect 117964 28432 118016 28484
rect 114928 28364 114980 28416
rect 115572 28364 115624 28416
rect 116952 28364 117004 28416
rect 117596 28407 117648 28416
rect 117596 28373 117605 28407
rect 117605 28373 117639 28407
rect 117639 28373 117648 28407
rect 117596 28364 117648 28373
rect 117780 28407 117832 28416
rect 117780 28373 117789 28407
rect 117789 28373 117823 28407
rect 117823 28373 117832 28407
rect 117780 28364 117832 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 113650 28262 113702 28314
rect 113714 28262 113766 28314
rect 113778 28262 113830 28314
rect 113842 28262 113894 28314
rect 113906 28262 113958 28314
rect 110236 28160 110288 28212
rect 113364 28160 113416 28212
rect 113548 28160 113600 28212
rect 114376 28160 114428 28212
rect 109776 28067 109828 28076
rect 109776 28033 109785 28067
rect 109785 28033 109819 28067
rect 109819 28033 109828 28067
rect 109776 28024 109828 28033
rect 109960 28067 110012 28076
rect 109960 28033 109969 28067
rect 109969 28033 110003 28067
rect 110003 28033 110012 28067
rect 109960 28024 110012 28033
rect 111064 28024 111116 28076
rect 112352 28092 112404 28144
rect 114008 28092 114060 28144
rect 111708 28067 111760 28076
rect 111708 28033 111717 28067
rect 111717 28033 111751 28067
rect 111751 28033 111760 28067
rect 111708 28024 111760 28033
rect 112260 28067 112312 28076
rect 112260 28033 112269 28067
rect 112269 28033 112303 28067
rect 112303 28033 112312 28067
rect 112260 28024 112312 28033
rect 112628 28024 112680 28076
rect 110788 27956 110840 28008
rect 113272 28024 113324 28076
rect 114100 27999 114152 28008
rect 114100 27965 114109 27999
rect 114109 27965 114143 27999
rect 114143 27965 114152 27999
rect 114100 27956 114152 27965
rect 114468 28067 114520 28076
rect 114468 28033 114477 28067
rect 114477 28033 114511 28067
rect 114511 28033 114520 28067
rect 114468 28024 114520 28033
rect 114560 28067 114612 28076
rect 114560 28033 114569 28067
rect 114569 28033 114603 28067
rect 114603 28033 114612 28067
rect 114560 28024 114612 28033
rect 114744 28092 114796 28144
rect 114836 28067 114888 28076
rect 114836 28033 114845 28067
rect 114845 28033 114879 28067
rect 114879 28033 114888 28067
rect 114836 28024 114888 28033
rect 115572 28067 115624 28076
rect 115572 28033 115581 28067
rect 115581 28033 115615 28067
rect 115615 28033 115624 28067
rect 115572 28024 115624 28033
rect 116032 28160 116084 28212
rect 116584 28160 116636 28212
rect 117780 28160 117832 28212
rect 116124 28067 116176 28076
rect 116124 28033 116133 28067
rect 116133 28033 116167 28067
rect 116167 28033 116176 28067
rect 116124 28024 116176 28033
rect 117136 28092 117188 28144
rect 118240 28160 118292 28212
rect 116584 28067 116636 28076
rect 116584 28033 116593 28067
rect 116593 28033 116627 28067
rect 116627 28033 116636 28067
rect 116584 28024 116636 28033
rect 116676 28067 116728 28076
rect 116676 28033 116685 28067
rect 116685 28033 116719 28067
rect 116719 28033 116728 28067
rect 116676 28024 116728 28033
rect 116860 28067 116912 28076
rect 116860 28033 116869 28067
rect 116869 28033 116903 28067
rect 116903 28033 116912 28067
rect 116860 28024 116912 28033
rect 116952 28024 117004 28076
rect 114376 27888 114428 27940
rect 117412 27999 117464 28008
rect 117412 27965 117421 27999
rect 117421 27965 117455 27999
rect 117455 27965 117464 27999
rect 117412 27956 117464 27965
rect 117688 28024 117740 28076
rect 118240 28067 118292 28076
rect 118240 28033 118249 28067
rect 118249 28033 118283 28067
rect 118283 28033 118292 28067
rect 118240 28024 118292 28033
rect 111892 27863 111944 27872
rect 111892 27829 111901 27863
rect 111901 27829 111935 27863
rect 111935 27829 111944 27863
rect 111892 27820 111944 27829
rect 112260 27820 112312 27872
rect 115020 27863 115072 27872
rect 115020 27829 115029 27863
rect 115029 27829 115063 27863
rect 115063 27829 115072 27863
rect 115020 27820 115072 27829
rect 116492 27863 116544 27872
rect 116492 27829 116501 27863
rect 116501 27829 116535 27863
rect 116535 27829 116544 27863
rect 116492 27820 116544 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 112914 27718 112966 27770
rect 112978 27718 113030 27770
rect 113042 27718 113094 27770
rect 113106 27718 113158 27770
rect 113170 27718 113222 27770
rect 109960 27616 110012 27668
rect 110052 27548 110104 27600
rect 111064 27591 111116 27600
rect 111064 27557 111073 27591
rect 111073 27557 111107 27591
rect 111107 27557 111116 27591
rect 111064 27548 111116 27557
rect 109868 27523 109920 27532
rect 109868 27489 109877 27523
rect 109877 27489 109911 27523
rect 109911 27489 109920 27523
rect 109868 27480 109920 27489
rect 112260 27548 112312 27600
rect 114468 27659 114520 27668
rect 114468 27625 114477 27659
rect 114477 27625 114511 27659
rect 114511 27625 114520 27659
rect 114468 27616 114520 27625
rect 116124 27616 116176 27668
rect 117044 27616 117096 27668
rect 118240 27659 118292 27668
rect 118240 27625 118249 27659
rect 118249 27625 118283 27659
rect 118283 27625 118292 27659
rect 118240 27616 118292 27625
rect 111248 27480 111300 27532
rect 110972 27412 111024 27464
rect 111340 27455 111392 27464
rect 111340 27421 111349 27455
rect 111349 27421 111383 27455
rect 111383 27421 111392 27455
rect 111340 27412 111392 27421
rect 111892 27480 111944 27532
rect 112260 27455 112312 27464
rect 112260 27421 112269 27455
rect 112269 27421 112303 27455
rect 112303 27421 112312 27455
rect 112260 27412 112312 27421
rect 113548 27591 113600 27600
rect 113548 27557 113557 27591
rect 113557 27557 113591 27591
rect 113591 27557 113600 27591
rect 113548 27548 113600 27557
rect 113272 27523 113324 27532
rect 113272 27489 113281 27523
rect 113281 27489 113315 27523
rect 113315 27489 113324 27523
rect 113272 27480 113324 27489
rect 114100 27480 114152 27532
rect 114652 27455 114704 27464
rect 114652 27421 114661 27455
rect 114661 27421 114695 27455
rect 114695 27421 114704 27455
rect 114652 27412 114704 27421
rect 115296 27480 115348 27532
rect 114928 27455 114980 27464
rect 114928 27421 114937 27455
rect 114937 27421 114971 27455
rect 114971 27421 114980 27455
rect 114928 27412 114980 27421
rect 115020 27455 115072 27464
rect 115020 27421 115029 27455
rect 115029 27421 115063 27455
rect 115063 27421 115072 27455
rect 115020 27412 115072 27421
rect 112536 27387 112588 27396
rect 112536 27353 112545 27387
rect 112545 27353 112579 27387
rect 112579 27353 112588 27387
rect 112536 27344 112588 27353
rect 112720 27387 112772 27396
rect 112720 27353 112729 27387
rect 112729 27353 112763 27387
rect 112763 27353 112772 27387
rect 112720 27344 112772 27353
rect 111984 27276 112036 27328
rect 112168 27319 112220 27328
rect 112168 27285 112177 27319
rect 112177 27285 112211 27319
rect 112211 27285 112220 27319
rect 115388 27344 115440 27396
rect 115940 27412 115992 27464
rect 116124 27412 116176 27464
rect 117412 27548 117464 27600
rect 118332 27591 118384 27600
rect 118332 27557 118341 27591
rect 118341 27557 118375 27591
rect 118375 27557 118384 27591
rect 118332 27548 118384 27557
rect 116768 27523 116820 27532
rect 116768 27489 116777 27523
rect 116777 27489 116811 27523
rect 116811 27489 116820 27523
rect 116768 27480 116820 27489
rect 117596 27480 117648 27532
rect 116584 27412 116636 27464
rect 116860 27412 116912 27464
rect 118148 27412 118200 27464
rect 118516 27455 118568 27464
rect 118516 27421 118525 27455
rect 118525 27421 118559 27455
rect 118559 27421 118568 27455
rect 118516 27412 118568 27421
rect 116492 27344 116544 27396
rect 112168 27276 112220 27285
rect 114100 27319 114152 27328
rect 114100 27285 114109 27319
rect 114109 27285 114143 27319
rect 114143 27285 114152 27319
rect 114100 27276 114152 27285
rect 115664 27319 115716 27328
rect 115664 27285 115673 27319
rect 115673 27285 115707 27319
rect 115707 27285 115716 27319
rect 115664 27276 115716 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 113650 27174 113702 27226
rect 113714 27174 113766 27226
rect 113778 27174 113830 27226
rect 113842 27174 113894 27226
rect 113906 27174 113958 27226
rect 110788 27115 110840 27124
rect 110788 27081 110797 27115
rect 110797 27081 110831 27115
rect 110831 27081 110840 27115
rect 110788 27072 110840 27081
rect 114008 27072 114060 27124
rect 114836 27072 114888 27124
rect 115296 27115 115348 27124
rect 115296 27081 115305 27115
rect 115305 27081 115339 27115
rect 115339 27081 115348 27115
rect 115296 27072 115348 27081
rect 115388 27115 115440 27124
rect 115388 27081 115397 27115
rect 115397 27081 115431 27115
rect 115431 27081 115440 27115
rect 115388 27072 115440 27081
rect 118516 27115 118568 27124
rect 118516 27081 118525 27115
rect 118525 27081 118559 27115
rect 118559 27081 118568 27115
rect 118516 27072 118568 27081
rect 110972 26979 111024 26988
rect 110972 26945 110981 26979
rect 110981 26945 111015 26979
rect 111015 26945 111024 26979
rect 110972 26936 111024 26945
rect 112168 27004 112220 27056
rect 112536 27004 112588 27056
rect 116124 27047 116176 27056
rect 116124 27013 116133 27047
rect 116133 27013 116167 27047
rect 116167 27013 116176 27047
rect 116124 27004 116176 27013
rect 111248 26979 111300 26988
rect 111248 26945 111257 26979
rect 111257 26945 111291 26979
rect 111291 26945 111300 26979
rect 111248 26936 111300 26945
rect 111340 26979 111392 26988
rect 111340 26945 111349 26979
rect 111349 26945 111383 26979
rect 111383 26945 111392 26979
rect 111340 26936 111392 26945
rect 112076 26979 112128 26988
rect 112076 26945 112085 26979
rect 112085 26945 112119 26979
rect 112119 26945 112128 26979
rect 112076 26936 112128 26945
rect 113548 26979 113600 26988
rect 113548 26945 113557 26979
rect 113557 26945 113591 26979
rect 113591 26945 113600 26979
rect 113548 26936 113600 26945
rect 114744 26936 114796 26988
rect 112352 26868 112404 26920
rect 114652 26911 114704 26920
rect 114652 26877 114661 26911
rect 114661 26877 114695 26911
rect 114695 26877 114704 26911
rect 114652 26868 114704 26877
rect 115664 26979 115716 26988
rect 115664 26945 115673 26979
rect 115673 26945 115707 26979
rect 115707 26945 115716 26979
rect 115664 26936 115716 26945
rect 115848 26979 115900 26988
rect 115848 26945 115857 26979
rect 115857 26945 115891 26979
rect 115891 26945 115900 26979
rect 115848 26936 115900 26945
rect 115848 26775 115900 26784
rect 115848 26741 115857 26775
rect 115857 26741 115891 26775
rect 115891 26741 115900 26775
rect 115848 26732 115900 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 112914 26630 112966 26682
rect 112978 26630 113030 26682
rect 113042 26630 113094 26682
rect 113106 26630 113158 26682
rect 113170 26630 113222 26682
rect 111248 26528 111300 26580
rect 114100 26528 114152 26580
rect 115296 26571 115348 26580
rect 115296 26537 115305 26571
rect 115305 26537 115339 26571
rect 115339 26537 115348 26571
rect 115296 26528 115348 26537
rect 115848 26528 115900 26580
rect 109868 26324 109920 26376
rect 112720 26392 112772 26444
rect 112536 26324 112588 26376
rect 115020 26299 115072 26308
rect 115020 26265 115029 26299
rect 115029 26265 115063 26299
rect 115063 26265 115072 26299
rect 115020 26256 115072 26265
rect 115388 26256 115440 26308
rect 114744 26188 114796 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 113650 26086 113702 26138
rect 113714 26086 113766 26138
rect 113778 26086 113830 26138
rect 113842 26086 113894 26138
rect 113906 26086 113958 26138
rect 115388 25984 115440 26036
rect 114744 25916 114796 25968
rect 115296 25848 115348 25900
rect 115020 25712 115072 25764
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 112914 25542 112966 25594
rect 112978 25542 113030 25594
rect 113042 25542 113094 25594
rect 113106 25542 113158 25594
rect 113170 25542 113222 25594
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 113650 24998 113702 25050
rect 113714 24998 113766 25050
rect 113778 24998 113830 25050
rect 113842 24998 113894 25050
rect 113906 24998 113958 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 112914 24454 112966 24506
rect 112978 24454 113030 24506
rect 113042 24454 113094 24506
rect 113106 24454 113158 24506
rect 113170 24454 113222 24506
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 113650 23910 113702 23962
rect 113714 23910 113766 23962
rect 113778 23910 113830 23962
rect 113842 23910 113894 23962
rect 113906 23910 113958 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 112914 23366 112966 23418
rect 112978 23366 113030 23418
rect 113042 23366 113094 23418
rect 113106 23366 113158 23418
rect 113170 23366 113222 23418
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 113650 22822 113702 22874
rect 113714 22822 113766 22874
rect 113778 22822 113830 22874
rect 113842 22822 113894 22874
rect 113906 22822 113958 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 112914 22278 112966 22330
rect 112978 22278 113030 22330
rect 113042 22278 113094 22330
rect 113106 22278 113158 22330
rect 113170 22278 113222 22330
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 113650 21734 113702 21786
rect 113714 21734 113766 21786
rect 113778 21734 113830 21786
rect 113842 21734 113894 21786
rect 113906 21734 113958 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 112914 21190 112966 21242
rect 112978 21190 113030 21242
rect 113042 21190 113094 21242
rect 113106 21190 113158 21242
rect 113170 21190 113222 21242
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 113650 20646 113702 20698
rect 113714 20646 113766 20698
rect 113778 20646 113830 20698
rect 113842 20646 113894 20698
rect 113906 20646 113958 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 112914 20102 112966 20154
rect 112978 20102 113030 20154
rect 113042 20102 113094 20154
rect 113106 20102 113158 20154
rect 113170 20102 113222 20154
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 113650 19558 113702 19610
rect 113714 19558 113766 19610
rect 113778 19558 113830 19610
rect 113842 19558 113894 19610
rect 113906 19558 113958 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 112914 19014 112966 19066
rect 112978 19014 113030 19066
rect 113042 19014 113094 19066
rect 113106 19014 113158 19066
rect 113170 19014 113222 19066
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 113650 18470 113702 18522
rect 113714 18470 113766 18522
rect 113778 18470 113830 18522
rect 113842 18470 113894 18522
rect 113906 18470 113958 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 112914 17926 112966 17978
rect 112978 17926 113030 17978
rect 113042 17926 113094 17978
rect 113106 17926 113158 17978
rect 113170 17926 113222 17978
rect 9680 17620 9732 17672
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 113650 17382 113702 17434
rect 113714 17382 113766 17434
rect 113778 17382 113830 17434
rect 113842 17382 113894 17434
rect 113906 17382 113958 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 112914 16838 112966 16890
rect 112978 16838 113030 16890
rect 113042 16838 113094 16890
rect 113106 16838 113158 16890
rect 113170 16838 113222 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 113650 16294 113702 16346
rect 113714 16294 113766 16346
rect 113778 16294 113830 16346
rect 113842 16294 113894 16346
rect 113906 16294 113958 16346
rect 1308 16056 1360 16108
rect 9680 15920 9732 15972
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 112914 15750 112966 15802
rect 112978 15750 113030 15802
rect 113042 15750 113094 15802
rect 113106 15750 113158 15802
rect 113170 15750 113222 15802
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 113650 15206 113702 15258
rect 113714 15206 113766 15258
rect 113778 15206 113830 15258
rect 113842 15206 113894 15258
rect 113906 15206 113958 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 112914 14662 112966 14714
rect 112978 14662 113030 14714
rect 113042 14662 113094 14714
rect 113106 14662 113158 14714
rect 113170 14662 113222 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 113650 14118 113702 14170
rect 113714 14118 113766 14170
rect 113778 14118 113830 14170
rect 113842 14118 113894 14170
rect 113906 14118 113958 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 112914 13574 112966 13626
rect 112978 13574 113030 13626
rect 113042 13574 113094 13626
rect 113106 13574 113158 13626
rect 113170 13574 113222 13626
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 113650 13030 113702 13082
rect 113714 13030 113766 13082
rect 113778 13030 113830 13082
rect 113842 13030 113894 13082
rect 113906 13030 113958 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 112914 12486 112966 12538
rect 112978 12486 113030 12538
rect 113042 12486 113094 12538
rect 113106 12486 113158 12538
rect 113170 12486 113222 12538
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 113650 11942 113702 11994
rect 113714 11942 113766 11994
rect 113778 11942 113830 11994
rect 113842 11942 113894 11994
rect 113906 11942 113958 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 112914 11398 112966 11450
rect 112978 11398 113030 11450
rect 113042 11398 113094 11450
rect 113106 11398 113158 11450
rect 113170 11398 113222 11450
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 113650 10854 113702 10906
rect 113714 10854 113766 10906
rect 113778 10854 113830 10906
rect 113842 10854 113894 10906
rect 113906 10854 113958 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 112914 10310 112966 10362
rect 112978 10310 113030 10362
rect 113042 10310 113094 10362
rect 113106 10310 113158 10362
rect 113170 10310 113222 10362
rect 93400 10004 93452 10056
rect 109500 10004 109552 10056
rect 92848 9936 92900 9988
rect 108304 9936 108356 9988
rect 93032 9868 93084 9920
rect 106464 9868 106516 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 113650 9766 113702 9818
rect 113714 9766 113766 9818
rect 113778 9766 113830 9818
rect 113842 9766 113894 9818
rect 113906 9766 113958 9818
rect 8208 9596 8260 9648
rect 15844 9596 15896 9648
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 112914 9222 112966 9274
rect 112978 9222 113030 9274
rect 113042 9222 113094 9274
rect 113106 9222 113158 9274
rect 113170 9222 113222 9274
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 113650 8678 113702 8730
rect 113714 8678 113766 8730
rect 113778 8678 113830 8730
rect 113842 8678 113894 8730
rect 113906 8678 113958 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 112914 8134 112966 8186
rect 112978 8134 113030 8186
rect 113042 8134 113094 8186
rect 113106 8134 113158 8186
rect 113170 8134 113222 8186
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 66314 7590 66366 7642
rect 66378 7590 66430 7642
rect 66442 7590 66494 7642
rect 66506 7590 66558 7642
rect 66570 7590 66622 7642
rect 97034 7590 97086 7642
rect 97098 7590 97150 7642
rect 97162 7590 97214 7642
rect 97226 7590 97278 7642
rect 97290 7590 97342 7642
rect 113650 7590 113702 7642
rect 113714 7590 113766 7642
rect 113778 7590 113830 7642
rect 113842 7590 113894 7642
rect 113906 7590 113958 7642
rect 15844 7488 15896 7540
rect 26976 7531 27028 7540
rect 26976 7497 26985 7531
rect 26985 7497 27019 7531
rect 27019 7497 27028 7531
rect 26976 7488 27028 7497
rect 27804 7488 27856 7540
rect 29552 7531 29604 7540
rect 29552 7497 29561 7531
rect 29561 7497 29595 7531
rect 29595 7497 29604 7531
rect 29552 7488 29604 7497
rect 30196 7531 30248 7540
rect 30196 7497 30205 7531
rect 30205 7497 30239 7531
rect 30239 7497 30248 7531
rect 30196 7488 30248 7497
rect 92848 7531 92900 7540
rect 92848 7497 92857 7531
rect 92857 7497 92891 7531
rect 92891 7497 92900 7531
rect 92848 7488 92900 7497
rect 93032 7531 93084 7540
rect 93032 7497 93041 7531
rect 93041 7497 93075 7531
rect 93075 7497 93084 7531
rect 93032 7488 93084 7497
rect 93216 7531 93268 7540
rect 93216 7497 93225 7531
rect 93225 7497 93259 7531
rect 93259 7497 93268 7531
rect 93216 7488 93268 7497
rect 93400 7531 93452 7540
rect 93400 7497 93409 7531
rect 93409 7497 93443 7531
rect 93443 7497 93452 7531
rect 93400 7488 93452 7497
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 112914 7046 112966 7098
rect 112978 7046 113030 7098
rect 113042 7046 113094 7098
rect 113106 7046 113158 7098
rect 113170 7046 113222 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 66314 6502 66366 6554
rect 66378 6502 66430 6554
rect 66442 6502 66494 6554
rect 66506 6502 66558 6554
rect 66570 6502 66622 6554
rect 97034 6502 97086 6554
rect 97098 6502 97150 6554
rect 97162 6502 97214 6554
rect 97226 6502 97278 6554
rect 97290 6502 97342 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 66314 5414 66366 5466
rect 66378 5414 66430 5466
rect 66442 5414 66494 5466
rect 66506 5414 66558 5466
rect 66570 5414 66622 5466
rect 97034 5414 97086 5466
rect 97098 5414 97150 5466
rect 97162 5414 97214 5466
rect 97226 5414 97278 5466
rect 97290 5414 97342 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 66314 4326 66366 4378
rect 66378 4326 66430 4378
rect 66442 4326 66494 4378
rect 66506 4326 66558 4378
rect 66570 4326 66622 4378
rect 97034 4326 97086 4378
rect 97098 4326 97150 4378
rect 97162 4326 97214 4378
rect 97226 4326 97278 4378
rect 97290 4326 97342 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 66314 3238 66366 3290
rect 66378 3238 66430 3290
rect 66442 3238 66494 3290
rect 66506 3238 66558 3290
rect 66570 3238 66622 3290
rect 97034 3238 97086 3290
rect 97098 3238 97150 3290
rect 97162 3238 97214 3290
rect 97226 3238 97278 3290
rect 97290 3238 97342 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 25872 2635 25924 2644
rect 25872 2601 25881 2635
rect 25881 2601 25915 2635
rect 25915 2601 25924 2635
rect 25872 2592 25924 2601
rect 31668 2635 31720 2644
rect 31668 2601 31677 2635
rect 31677 2601 31711 2635
rect 31711 2601 31720 2635
rect 31668 2592 31720 2601
rect 32956 2635 33008 2644
rect 32956 2601 32965 2635
rect 32965 2601 32999 2635
rect 32999 2601 33008 2635
rect 32956 2592 33008 2601
rect 33784 2635 33836 2644
rect 33784 2601 33793 2635
rect 33793 2601 33827 2635
rect 33827 2601 33836 2635
rect 33784 2592 33836 2601
rect 34796 2592 34848 2644
rect 36176 2635 36228 2644
rect 36176 2601 36185 2635
rect 36185 2601 36219 2635
rect 36219 2601 36228 2635
rect 36176 2592 36228 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 38292 2635 38344 2644
rect 38292 2601 38301 2635
rect 38301 2601 38335 2635
rect 38335 2601 38344 2635
rect 38292 2592 38344 2601
rect 40040 2635 40092 2644
rect 40040 2601 40049 2635
rect 40049 2601 40083 2635
rect 40083 2601 40092 2635
rect 40040 2592 40092 2601
rect 40868 2635 40920 2644
rect 40868 2601 40877 2635
rect 40877 2601 40911 2635
rect 40911 2601 40920 2635
rect 40868 2592 40920 2601
rect 41972 2635 42024 2644
rect 41972 2601 41981 2635
rect 41981 2601 42015 2635
rect 42015 2601 42024 2635
rect 41972 2592 42024 2601
rect 43260 2635 43312 2644
rect 43260 2601 43269 2635
rect 43269 2601 43303 2635
rect 43303 2601 43312 2635
rect 43260 2592 43312 2601
rect 44548 2635 44600 2644
rect 44548 2601 44557 2635
rect 44557 2601 44591 2635
rect 44591 2601 44600 2635
rect 44548 2592 44600 2601
rect 45836 2635 45888 2644
rect 45836 2601 45845 2635
rect 45845 2601 45879 2635
rect 45879 2601 45888 2635
rect 45836 2592 45888 2601
rect 46664 2635 46716 2644
rect 46664 2601 46673 2635
rect 46673 2601 46707 2635
rect 46707 2601 46716 2635
rect 46664 2592 46716 2601
rect 47768 2635 47820 2644
rect 47768 2601 47777 2635
rect 47777 2601 47811 2635
rect 47811 2601 47820 2635
rect 47768 2592 47820 2601
rect 49056 2635 49108 2644
rect 49056 2601 49065 2635
rect 49065 2601 49099 2635
rect 49099 2601 49108 2635
rect 49056 2592 49108 2601
rect 50344 2635 50396 2644
rect 50344 2601 50353 2635
rect 50353 2601 50387 2635
rect 50387 2601 50396 2635
rect 50344 2592 50396 2601
rect 51632 2635 51684 2644
rect 51632 2601 51641 2635
rect 51641 2601 51675 2635
rect 51675 2601 51684 2635
rect 51632 2592 51684 2601
rect 52460 2635 52512 2644
rect 52460 2601 52469 2635
rect 52469 2601 52503 2635
rect 52503 2601 52512 2635
rect 52460 2592 52512 2601
rect 53564 2635 53616 2644
rect 53564 2601 53573 2635
rect 53573 2601 53607 2635
rect 53607 2601 53616 2635
rect 53564 2592 53616 2601
rect 55036 2635 55088 2644
rect 55036 2601 55045 2635
rect 55045 2601 55079 2635
rect 55079 2601 55088 2635
rect 55036 2592 55088 2601
rect 56140 2635 56192 2644
rect 56140 2601 56149 2635
rect 56149 2601 56183 2635
rect 56183 2601 56192 2635
rect 56140 2592 56192 2601
rect 57428 2635 57480 2644
rect 57428 2601 57437 2635
rect 57437 2601 57471 2635
rect 57471 2601 57480 2635
rect 57428 2592 57480 2601
rect 58256 2635 58308 2644
rect 58256 2601 58265 2635
rect 58265 2601 58299 2635
rect 58299 2601 58308 2635
rect 58256 2592 58308 2601
rect 59544 2635 59596 2644
rect 59544 2601 59553 2635
rect 59553 2601 59587 2635
rect 59587 2601 59596 2635
rect 59544 2592 59596 2601
rect 60832 2635 60884 2644
rect 60832 2601 60841 2635
rect 60841 2601 60875 2635
rect 60875 2601 60884 2635
rect 60832 2592 60884 2601
rect 61936 2635 61988 2644
rect 61936 2601 61945 2635
rect 61945 2601 61979 2635
rect 61979 2601 61988 2635
rect 61936 2592 61988 2601
rect 63224 2635 63276 2644
rect 63224 2601 63233 2635
rect 63233 2601 63267 2635
rect 63267 2601 63276 2635
rect 63224 2592 63276 2601
rect 64052 2635 64104 2644
rect 64052 2601 64061 2635
rect 64061 2601 64095 2635
rect 64095 2601 64104 2635
rect 64052 2592 64104 2601
rect 65340 2635 65392 2644
rect 65340 2601 65349 2635
rect 65349 2601 65383 2635
rect 65383 2601 65392 2635
rect 65340 2592 65392 2601
rect 66720 2592 66772 2644
rect 67732 2635 67784 2644
rect 67732 2601 67741 2635
rect 67741 2601 67775 2635
rect 67775 2601 67784 2635
rect 67732 2592 67784 2601
rect 25780 2295 25832 2304
rect 25780 2261 25789 2295
rect 25789 2261 25823 2295
rect 25823 2261 25832 2295
rect 25780 2252 25832 2261
rect 31576 2295 31628 2304
rect 31576 2261 31585 2295
rect 31585 2261 31619 2295
rect 31619 2261 31628 2295
rect 31576 2252 31628 2261
rect 32864 2295 32916 2304
rect 32864 2261 32873 2295
rect 32873 2261 32907 2295
rect 32907 2261 32916 2295
rect 32864 2252 32916 2261
rect 33508 2295 33560 2304
rect 33508 2261 33517 2295
rect 33517 2261 33551 2295
rect 33551 2261 33560 2295
rect 33508 2252 33560 2261
rect 34796 2295 34848 2304
rect 34796 2261 34805 2295
rect 34805 2261 34839 2295
rect 34839 2261 34848 2295
rect 34796 2252 34848 2261
rect 36084 2295 36136 2304
rect 36084 2261 36093 2295
rect 36093 2261 36127 2295
rect 36127 2261 36136 2295
rect 36084 2252 36136 2261
rect 37372 2295 37424 2304
rect 37372 2261 37381 2295
rect 37381 2261 37415 2295
rect 37415 2261 37424 2295
rect 37372 2252 37424 2261
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 39948 2295 40000 2304
rect 39948 2261 39957 2295
rect 39957 2261 39991 2295
rect 39991 2261 40000 2295
rect 39948 2252 40000 2261
rect 40592 2295 40644 2304
rect 40592 2261 40601 2295
rect 40601 2261 40635 2295
rect 40635 2261 40644 2295
rect 40592 2252 40644 2261
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 43168 2295 43220 2304
rect 43168 2261 43177 2295
rect 43177 2261 43211 2295
rect 43211 2261 43220 2295
rect 43168 2252 43220 2261
rect 44456 2295 44508 2304
rect 44456 2261 44465 2295
rect 44465 2261 44499 2295
rect 44499 2261 44508 2295
rect 44456 2252 44508 2261
rect 45744 2295 45796 2304
rect 45744 2261 45753 2295
rect 45753 2261 45787 2295
rect 45787 2261 45796 2295
rect 45744 2252 45796 2261
rect 46388 2295 46440 2304
rect 46388 2261 46397 2295
rect 46397 2261 46431 2295
rect 46431 2261 46440 2295
rect 46388 2252 46440 2261
rect 47676 2295 47728 2304
rect 47676 2261 47685 2295
rect 47685 2261 47719 2295
rect 47719 2261 47728 2295
rect 47676 2252 47728 2261
rect 48964 2295 49016 2304
rect 48964 2261 48973 2295
rect 48973 2261 49007 2295
rect 49007 2261 49016 2295
rect 48964 2252 49016 2261
rect 50252 2295 50304 2304
rect 50252 2261 50261 2295
rect 50261 2261 50295 2295
rect 50295 2261 50304 2295
rect 50252 2252 50304 2261
rect 51540 2295 51592 2304
rect 51540 2261 51549 2295
rect 51549 2261 51583 2295
rect 51583 2261 51592 2295
rect 51540 2252 51592 2261
rect 52184 2295 52236 2304
rect 52184 2261 52193 2295
rect 52193 2261 52227 2295
rect 52227 2261 52236 2295
rect 52184 2252 52236 2261
rect 53472 2295 53524 2304
rect 53472 2261 53481 2295
rect 53481 2261 53515 2295
rect 53515 2261 53524 2295
rect 53472 2252 53524 2261
rect 54760 2295 54812 2304
rect 54760 2261 54769 2295
rect 54769 2261 54803 2295
rect 54803 2261 54812 2295
rect 54760 2252 54812 2261
rect 56048 2295 56100 2304
rect 56048 2261 56057 2295
rect 56057 2261 56091 2295
rect 56091 2261 56100 2295
rect 56048 2252 56100 2261
rect 57336 2295 57388 2304
rect 57336 2261 57345 2295
rect 57345 2261 57379 2295
rect 57379 2261 57388 2295
rect 57336 2252 57388 2261
rect 57980 2295 58032 2304
rect 57980 2261 57989 2295
rect 57989 2261 58023 2295
rect 58023 2261 58032 2295
rect 57980 2252 58032 2261
rect 59268 2295 59320 2304
rect 59268 2261 59277 2295
rect 59277 2261 59311 2295
rect 59311 2261 59320 2295
rect 59268 2252 59320 2261
rect 60556 2295 60608 2304
rect 60556 2261 60565 2295
rect 60565 2261 60599 2295
rect 60599 2261 60608 2295
rect 60556 2252 60608 2261
rect 61844 2295 61896 2304
rect 61844 2261 61853 2295
rect 61853 2261 61887 2295
rect 61887 2261 61896 2295
rect 61844 2252 61896 2261
rect 63132 2295 63184 2304
rect 63132 2261 63141 2295
rect 63141 2261 63175 2295
rect 63175 2261 63184 2295
rect 63132 2252 63184 2261
rect 63776 2295 63828 2304
rect 63776 2261 63785 2295
rect 63785 2261 63819 2295
rect 63819 2261 63828 2295
rect 63776 2252 63828 2261
rect 65064 2295 65116 2304
rect 65064 2261 65073 2295
rect 65073 2261 65107 2295
rect 65107 2261 65116 2295
rect 65064 2252 65116 2261
rect 66720 2252 66772 2304
rect 67640 2295 67692 2304
rect 67640 2261 67649 2295
rect 67649 2261 67683 2295
rect 67683 2261 67692 2295
rect 67640 2252 67692 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 66314 2150 66366 2202
rect 66378 2150 66430 2202
rect 66442 2150 66494 2202
rect 66506 2150 66558 2202
rect 66570 2150 66622 2202
rect 97034 2150 97086 2202
rect 97098 2150 97150 2202
rect 97162 2150 97214 2202
rect 97226 2150 97278 2202
rect 97290 2150 97342 2202
<< metal2 >>
rect 56046 99362 56102 100000
rect 55784 99334 56102 99362
rect 4214 97404 4522 97413
rect 4214 97402 4220 97404
rect 4276 97402 4300 97404
rect 4356 97402 4380 97404
rect 4436 97402 4460 97404
rect 4516 97402 4522 97404
rect 4276 97350 4278 97402
rect 4458 97350 4460 97402
rect 4214 97348 4220 97350
rect 4276 97348 4300 97350
rect 4356 97348 4380 97350
rect 4436 97348 4460 97350
rect 4516 97348 4522 97350
rect 4214 97339 4522 97348
rect 34934 97404 35242 97413
rect 34934 97402 34940 97404
rect 34996 97402 35020 97404
rect 35076 97402 35100 97404
rect 35156 97402 35180 97404
rect 35236 97402 35242 97404
rect 34996 97350 34998 97402
rect 35178 97350 35180 97402
rect 34934 97348 34940 97350
rect 34996 97348 35020 97350
rect 35076 97348 35100 97350
rect 35156 97348 35180 97350
rect 35236 97348 35242 97350
rect 34934 97339 35242 97348
rect 55784 97306 55812 99334
rect 56046 99200 56102 99334
rect 57334 99362 57390 100000
rect 58622 99362 58678 100000
rect 59910 99362 59966 100000
rect 60554 99362 60610 100000
rect 62486 99362 62542 100000
rect 63130 99362 63186 100000
rect 64418 99362 64474 100000
rect 65062 99362 65118 100000
rect 66994 99362 67050 100000
rect 67638 99362 67694 100000
rect 68926 99362 68982 100000
rect 57334 99334 57744 99362
rect 57334 99200 57390 99334
rect 57716 97306 57744 99334
rect 58622 99334 58848 99362
rect 58622 99200 58678 99334
rect 58820 97306 58848 99334
rect 59910 99334 60136 99362
rect 59910 99200 59966 99334
rect 60108 97306 60136 99334
rect 60554 99334 60688 99362
rect 60554 99200 60610 99334
rect 60660 97306 60688 99334
rect 62486 99334 62712 99362
rect 62486 99200 62542 99334
rect 62684 97306 62712 99334
rect 63130 99334 63356 99362
rect 63130 99200 63186 99334
rect 63328 97306 63356 99334
rect 64418 99334 64644 99362
rect 64418 99200 64474 99334
rect 64616 97306 64644 99334
rect 65062 99334 65288 99362
rect 65062 99200 65118 99334
rect 65260 97306 65288 99334
rect 66994 99334 67220 99362
rect 66994 99200 67050 99334
rect 65654 97404 65962 97413
rect 65654 97402 65660 97404
rect 65716 97402 65740 97404
rect 65796 97402 65820 97404
rect 65876 97402 65900 97404
rect 65956 97402 65962 97404
rect 65716 97350 65718 97402
rect 65898 97350 65900 97402
rect 65654 97348 65660 97350
rect 65716 97348 65740 97350
rect 65796 97348 65820 97350
rect 65876 97348 65900 97350
rect 65956 97348 65962 97350
rect 65654 97339 65962 97348
rect 55772 97300 55824 97306
rect 55772 97242 55824 97248
rect 57704 97300 57756 97306
rect 57704 97242 57756 97248
rect 58808 97300 58860 97306
rect 58808 97242 58860 97248
rect 60096 97300 60148 97306
rect 60096 97242 60148 97248
rect 60648 97300 60700 97306
rect 60648 97242 60700 97248
rect 62672 97300 62724 97306
rect 62672 97242 62724 97248
rect 63316 97300 63368 97306
rect 63316 97242 63368 97248
rect 64604 97300 64656 97306
rect 64604 97242 64656 97248
rect 65248 97300 65300 97306
rect 65248 97242 65300 97248
rect 65340 97300 65392 97306
rect 65340 97242 65392 97248
rect 57428 97096 57480 97102
rect 57428 97038 57480 97044
rect 58164 97096 58216 97102
rect 58164 97038 58216 97044
rect 59268 97096 59320 97102
rect 59268 97038 59320 97044
rect 60556 97096 60608 97102
rect 60556 97038 60608 97044
rect 60924 97096 60976 97102
rect 60924 97038 60976 97044
rect 62856 97096 62908 97102
rect 62856 97038 62908 97044
rect 63500 97096 63552 97102
rect 63500 97038 63552 97044
rect 64972 97096 65024 97102
rect 64972 97038 65024 97044
rect 56600 97028 56652 97034
rect 56600 96970 56652 96976
rect 56232 96960 56284 96966
rect 56232 96902 56284 96908
rect 4874 96860 5182 96869
rect 4874 96858 4880 96860
rect 4936 96858 4960 96860
rect 5016 96858 5040 96860
rect 5096 96858 5120 96860
rect 5176 96858 5182 96860
rect 4936 96806 4938 96858
rect 5118 96806 5120 96858
rect 4874 96804 4880 96806
rect 4936 96804 4960 96806
rect 5016 96804 5040 96806
rect 5096 96804 5120 96806
rect 5176 96804 5182 96806
rect 4874 96795 5182 96804
rect 35594 96860 35902 96869
rect 35594 96858 35600 96860
rect 35656 96858 35680 96860
rect 35736 96858 35760 96860
rect 35816 96858 35840 96860
rect 35896 96858 35902 96860
rect 35656 96806 35658 96858
rect 35838 96806 35840 96858
rect 35594 96804 35600 96806
rect 35656 96804 35680 96806
rect 35736 96804 35760 96806
rect 35816 96804 35840 96806
rect 35896 96804 35902 96806
rect 35594 96795 35902 96804
rect 56244 96694 56272 96902
rect 56232 96688 56284 96694
rect 56232 96630 56284 96636
rect 4214 96316 4522 96325
rect 4214 96314 4220 96316
rect 4276 96314 4300 96316
rect 4356 96314 4380 96316
rect 4436 96314 4460 96316
rect 4516 96314 4522 96316
rect 4276 96262 4278 96314
rect 4458 96262 4460 96314
rect 4214 96260 4220 96262
rect 4276 96260 4300 96262
rect 4356 96260 4380 96262
rect 4436 96260 4460 96262
rect 4516 96260 4522 96262
rect 4214 96251 4522 96260
rect 34934 96316 35242 96325
rect 34934 96314 34940 96316
rect 34996 96314 35020 96316
rect 35076 96314 35100 96316
rect 35156 96314 35180 96316
rect 35236 96314 35242 96316
rect 34996 96262 34998 96314
rect 35178 96262 35180 96314
rect 34934 96260 34940 96262
rect 34996 96260 35020 96262
rect 35076 96260 35100 96262
rect 35156 96260 35180 96262
rect 35236 96260 35242 96262
rect 34934 96251 35242 96260
rect 4874 95772 5182 95781
rect 4874 95770 4880 95772
rect 4936 95770 4960 95772
rect 5016 95770 5040 95772
rect 5096 95770 5120 95772
rect 5176 95770 5182 95772
rect 4936 95718 4938 95770
rect 5118 95718 5120 95770
rect 4874 95716 4880 95718
rect 4936 95716 4960 95718
rect 5016 95716 5040 95718
rect 5096 95716 5120 95718
rect 5176 95716 5182 95718
rect 4874 95707 5182 95716
rect 35594 95772 35902 95781
rect 35594 95770 35600 95772
rect 35656 95770 35680 95772
rect 35736 95770 35760 95772
rect 35816 95770 35840 95772
rect 35896 95770 35902 95772
rect 35656 95718 35658 95770
rect 35838 95718 35840 95770
rect 35594 95716 35600 95718
rect 35656 95716 35680 95718
rect 35736 95716 35760 95718
rect 35816 95716 35840 95718
rect 35896 95716 35902 95718
rect 35594 95707 35902 95716
rect 54484 95600 54536 95606
rect 54484 95542 54536 95548
rect 4214 95228 4522 95237
rect 4214 95226 4220 95228
rect 4276 95226 4300 95228
rect 4356 95226 4380 95228
rect 4436 95226 4460 95228
rect 4516 95226 4522 95228
rect 4276 95174 4278 95226
rect 4458 95174 4460 95226
rect 4214 95172 4220 95174
rect 4276 95172 4300 95174
rect 4356 95172 4380 95174
rect 4436 95172 4460 95174
rect 4516 95172 4522 95174
rect 4214 95163 4522 95172
rect 34934 95228 35242 95237
rect 34934 95226 34940 95228
rect 34996 95226 35020 95228
rect 35076 95226 35100 95228
rect 35156 95226 35180 95228
rect 35236 95226 35242 95228
rect 34996 95174 34998 95226
rect 35178 95174 35180 95226
rect 34934 95172 34940 95174
rect 34996 95172 35020 95174
rect 35076 95172 35100 95174
rect 35156 95172 35180 95174
rect 35236 95172 35242 95174
rect 34934 95163 35242 95172
rect 4874 94684 5182 94693
rect 4874 94682 4880 94684
rect 4936 94682 4960 94684
rect 5016 94682 5040 94684
rect 5096 94682 5120 94684
rect 5176 94682 5182 94684
rect 4936 94630 4938 94682
rect 5118 94630 5120 94682
rect 4874 94628 4880 94630
rect 4936 94628 4960 94630
rect 5016 94628 5040 94630
rect 5096 94628 5120 94630
rect 5176 94628 5182 94630
rect 4874 94619 5182 94628
rect 35594 94684 35902 94693
rect 35594 94682 35600 94684
rect 35656 94682 35680 94684
rect 35736 94682 35760 94684
rect 35816 94682 35840 94684
rect 35896 94682 35902 94684
rect 35656 94630 35658 94682
rect 35838 94630 35840 94682
rect 35594 94628 35600 94630
rect 35656 94628 35680 94630
rect 35736 94628 35760 94630
rect 35816 94628 35840 94630
rect 35896 94628 35902 94630
rect 35594 94619 35902 94628
rect 52460 94444 52512 94450
rect 52460 94386 52512 94392
rect 4214 94140 4522 94149
rect 4214 94138 4220 94140
rect 4276 94138 4300 94140
rect 4356 94138 4380 94140
rect 4436 94138 4460 94140
rect 4516 94138 4522 94140
rect 4276 94086 4278 94138
rect 4458 94086 4460 94138
rect 4214 94084 4220 94086
rect 4276 94084 4300 94086
rect 4356 94084 4380 94086
rect 4436 94084 4460 94086
rect 4516 94084 4522 94086
rect 4214 94075 4522 94084
rect 34934 94140 35242 94149
rect 34934 94138 34940 94140
rect 34996 94138 35020 94140
rect 35076 94138 35100 94140
rect 35156 94138 35180 94140
rect 35236 94138 35242 94140
rect 34996 94086 34998 94138
rect 35178 94086 35180 94138
rect 34934 94084 34940 94086
rect 34996 94084 35020 94086
rect 35076 94084 35100 94086
rect 35156 94084 35180 94086
rect 35236 94084 35242 94086
rect 34934 94075 35242 94084
rect 4874 93596 5182 93605
rect 4874 93594 4880 93596
rect 4936 93594 4960 93596
rect 5016 93594 5040 93596
rect 5096 93594 5120 93596
rect 5176 93594 5182 93596
rect 4936 93542 4938 93594
rect 5118 93542 5120 93594
rect 4874 93540 4880 93542
rect 4936 93540 4960 93542
rect 5016 93540 5040 93542
rect 5096 93540 5120 93542
rect 5176 93540 5182 93542
rect 4874 93531 5182 93540
rect 35594 93596 35902 93605
rect 35594 93594 35600 93596
rect 35656 93594 35680 93596
rect 35736 93594 35760 93596
rect 35816 93594 35840 93596
rect 35896 93594 35902 93596
rect 35656 93542 35658 93594
rect 35838 93542 35840 93594
rect 35594 93540 35600 93542
rect 35656 93540 35680 93542
rect 35736 93540 35760 93542
rect 35816 93540 35840 93542
rect 35896 93540 35902 93542
rect 35594 93531 35902 93540
rect 49332 93356 49384 93362
rect 49332 93298 49384 93304
rect 46848 93288 46900 93294
rect 49344 93265 49372 93298
rect 49516 93288 49568 93294
rect 46848 93230 46900 93236
rect 49330 93256 49386 93265
rect 4214 93052 4522 93061
rect 4214 93050 4220 93052
rect 4276 93050 4300 93052
rect 4356 93050 4380 93052
rect 4436 93050 4460 93052
rect 4516 93050 4522 93052
rect 4276 92998 4278 93050
rect 4458 92998 4460 93050
rect 4214 92996 4220 92998
rect 4276 92996 4300 92998
rect 4356 92996 4380 92998
rect 4436 92996 4460 92998
rect 4516 92996 4522 92998
rect 4214 92987 4522 92996
rect 34934 93052 35242 93061
rect 34934 93050 34940 93052
rect 34996 93050 35020 93052
rect 35076 93050 35100 93052
rect 35156 93050 35180 93052
rect 35236 93050 35242 93052
rect 34996 92998 34998 93050
rect 35178 92998 35180 93050
rect 34934 92996 34940 92998
rect 34996 92996 35020 92998
rect 35076 92996 35100 92998
rect 35156 92996 35180 92998
rect 35236 92996 35242 92998
rect 34934 92987 35242 92996
rect 46860 92818 46888 93230
rect 49516 93230 49568 93236
rect 49330 93191 49332 93200
rect 49384 93191 49386 93200
rect 49332 93162 49384 93168
rect 46940 93152 46992 93158
rect 46940 93094 46992 93100
rect 46952 92954 46980 93094
rect 46940 92948 46992 92954
rect 46940 92890 46992 92896
rect 46848 92812 46900 92818
rect 46848 92754 46900 92760
rect 45652 92744 45704 92750
rect 45652 92686 45704 92692
rect 47122 92712 47178 92721
rect 44180 92676 44232 92682
rect 44180 92618 44232 92624
rect 44192 92585 44220 92618
rect 44178 92576 44234 92585
rect 4874 92508 5182 92517
rect 4874 92506 4880 92508
rect 4936 92506 4960 92508
rect 5016 92506 5040 92508
rect 5096 92506 5120 92508
rect 5176 92506 5182 92508
rect 4936 92454 4938 92506
rect 5118 92454 5120 92506
rect 4874 92452 4880 92454
rect 4936 92452 4960 92454
rect 5016 92452 5040 92454
rect 5096 92452 5120 92454
rect 5176 92452 5182 92454
rect 4874 92443 5182 92452
rect 35594 92508 35902 92517
rect 44178 92511 44234 92520
rect 35594 92506 35600 92508
rect 35656 92506 35680 92508
rect 35736 92506 35760 92508
rect 35816 92506 35840 92508
rect 35896 92506 35902 92508
rect 35656 92454 35658 92506
rect 35838 92454 35840 92506
rect 35594 92452 35600 92454
rect 35656 92452 35680 92454
rect 35736 92452 35760 92454
rect 35816 92452 35840 92454
rect 35896 92452 35902 92454
rect 35594 92443 35902 92452
rect 45664 92410 45692 92686
rect 47122 92647 47124 92656
rect 47176 92647 47178 92656
rect 47124 92618 47176 92624
rect 45652 92404 45704 92410
rect 45652 92346 45704 92352
rect 45664 92070 45692 92346
rect 49528 92274 49556 93230
rect 52184 93152 52236 93158
rect 52184 93094 52236 93100
rect 52196 92954 52224 93094
rect 52472 92954 52500 94386
rect 53840 94376 53892 94382
rect 53840 94318 53892 94324
rect 53380 93696 53432 93702
rect 53380 93638 53432 93644
rect 52184 92948 52236 92954
rect 52184 92890 52236 92896
rect 52460 92948 52512 92954
rect 52460 92890 52512 92896
rect 50618 92848 50674 92857
rect 50618 92783 50620 92792
rect 50672 92783 50674 92792
rect 50620 92754 50672 92760
rect 53392 92750 53420 93638
rect 53852 93294 53880 94318
rect 54496 93498 54524 95542
rect 55680 95464 55732 95470
rect 55680 95406 55732 95412
rect 54668 94988 54720 94994
rect 54668 94930 54720 94936
rect 54680 94382 54708 94930
rect 55220 94784 55272 94790
rect 55220 94726 55272 94732
rect 54668 94376 54720 94382
rect 54668 94318 54720 94324
rect 54484 93492 54536 93498
rect 54484 93434 54536 93440
rect 54668 93356 54720 93362
rect 54668 93298 54720 93304
rect 53840 93288 53892 93294
rect 53840 93230 53892 93236
rect 53932 93288 53984 93294
rect 53932 93230 53984 93236
rect 53944 92954 53972 93230
rect 53932 92948 53984 92954
rect 53932 92890 53984 92896
rect 53380 92744 53432 92750
rect 52550 92712 52606 92721
rect 53380 92686 53432 92692
rect 52550 92647 52552 92656
rect 52604 92647 52606 92656
rect 52552 92618 52604 92624
rect 52920 92336 52972 92342
rect 52920 92278 52972 92284
rect 49516 92268 49568 92274
rect 49516 92210 49568 92216
rect 52932 92177 52960 92278
rect 53392 92274 53420 92686
rect 54024 92676 54076 92682
rect 54024 92618 54076 92624
rect 54036 92585 54064 92618
rect 54022 92576 54078 92585
rect 54022 92511 54078 92520
rect 54680 92410 54708 93298
rect 54668 92404 54720 92410
rect 54668 92346 54720 92352
rect 54852 92404 54904 92410
rect 54852 92346 54904 92352
rect 53380 92268 53432 92274
rect 53380 92210 53432 92216
rect 53196 92200 53248 92206
rect 50250 92168 50306 92177
rect 50250 92103 50252 92112
rect 50304 92103 50306 92112
rect 52918 92168 52974 92177
rect 53196 92142 53248 92148
rect 52918 92103 52974 92112
rect 50252 92074 50304 92080
rect 53208 92070 53236 92142
rect 54864 92070 54892 92346
rect 8208 92064 8260 92070
rect 8208 92006 8260 92012
rect 45652 92064 45704 92070
rect 45652 92006 45704 92012
rect 46848 92064 46900 92070
rect 46848 92006 46900 92012
rect 49608 92064 49660 92070
rect 53196 92064 53248 92070
rect 49608 92006 49660 92012
rect 53194 92032 53196 92041
rect 54852 92064 54904 92070
rect 53248 92032 53250 92041
rect 4214 91964 4522 91973
rect 4214 91962 4220 91964
rect 4276 91962 4300 91964
rect 4356 91962 4380 91964
rect 4436 91962 4460 91964
rect 4516 91962 4522 91964
rect 4276 91910 4278 91962
rect 4458 91910 4460 91962
rect 4214 91908 4220 91910
rect 4276 91908 4300 91910
rect 4356 91908 4380 91910
rect 4436 91908 4460 91910
rect 4516 91908 4522 91910
rect 4214 91899 4522 91908
rect 4874 91420 5182 91429
rect 4874 91418 4880 91420
rect 4936 91418 4960 91420
rect 5016 91418 5040 91420
rect 5096 91418 5120 91420
rect 5176 91418 5182 91420
rect 4936 91366 4938 91418
rect 5118 91366 5120 91418
rect 4874 91364 4880 91366
rect 4936 91364 4960 91366
rect 5016 91364 5040 91366
rect 5096 91364 5120 91366
rect 5176 91364 5182 91366
rect 4874 91355 5182 91364
rect 4214 90876 4522 90885
rect 4214 90874 4220 90876
rect 4276 90874 4300 90876
rect 4356 90874 4380 90876
rect 4436 90874 4460 90876
rect 4516 90874 4522 90876
rect 4276 90822 4278 90874
rect 4458 90822 4460 90874
rect 4214 90820 4220 90822
rect 4276 90820 4300 90822
rect 4356 90820 4380 90822
rect 4436 90820 4460 90822
rect 4516 90820 4522 90822
rect 4214 90811 4522 90820
rect 4874 90332 5182 90341
rect 4874 90330 4880 90332
rect 4936 90330 4960 90332
rect 5016 90330 5040 90332
rect 5096 90330 5120 90332
rect 5176 90330 5182 90332
rect 4936 90278 4938 90330
rect 5118 90278 5120 90330
rect 4874 90276 4880 90278
rect 4936 90276 4960 90278
rect 5016 90276 5040 90278
rect 5096 90276 5120 90278
rect 5176 90276 5182 90278
rect 4874 90267 5182 90276
rect 4214 89788 4522 89797
rect 4214 89786 4220 89788
rect 4276 89786 4300 89788
rect 4356 89786 4380 89788
rect 4436 89786 4460 89788
rect 4516 89786 4522 89788
rect 4276 89734 4278 89786
rect 4458 89734 4460 89786
rect 4214 89732 4220 89734
rect 4276 89732 4300 89734
rect 4356 89732 4380 89734
rect 4436 89732 4460 89734
rect 4516 89732 4522 89734
rect 4214 89723 4522 89732
rect 4874 89244 5182 89253
rect 4874 89242 4880 89244
rect 4936 89242 4960 89244
rect 5016 89242 5040 89244
rect 5096 89242 5120 89244
rect 5176 89242 5182 89244
rect 4936 89190 4938 89242
rect 5118 89190 5120 89242
rect 4874 89188 4880 89190
rect 4936 89188 4960 89190
rect 5016 89188 5040 89190
rect 5096 89188 5120 89190
rect 5176 89188 5182 89190
rect 4874 89179 5182 89188
rect 4214 88700 4522 88709
rect 4214 88698 4220 88700
rect 4276 88698 4300 88700
rect 4356 88698 4380 88700
rect 4436 88698 4460 88700
rect 4516 88698 4522 88700
rect 4276 88646 4278 88698
rect 4458 88646 4460 88698
rect 4214 88644 4220 88646
rect 4276 88644 4300 88646
rect 4356 88644 4380 88646
rect 4436 88644 4460 88646
rect 4516 88644 4522 88646
rect 4214 88635 4522 88644
rect 4874 88156 5182 88165
rect 4874 88154 4880 88156
rect 4936 88154 4960 88156
rect 5016 88154 5040 88156
rect 5096 88154 5120 88156
rect 5176 88154 5182 88156
rect 4936 88102 4938 88154
rect 5118 88102 5120 88154
rect 4874 88100 4880 88102
rect 4936 88100 4960 88102
rect 5016 88100 5040 88102
rect 5096 88100 5120 88102
rect 5176 88100 5182 88102
rect 4874 88091 5182 88100
rect 4214 87612 4522 87621
rect 4214 87610 4220 87612
rect 4276 87610 4300 87612
rect 4356 87610 4380 87612
rect 4436 87610 4460 87612
rect 4516 87610 4522 87612
rect 4276 87558 4278 87610
rect 4458 87558 4460 87610
rect 4214 87556 4220 87558
rect 4276 87556 4300 87558
rect 4356 87556 4380 87558
rect 4436 87556 4460 87558
rect 4516 87556 4522 87558
rect 4214 87547 4522 87556
rect 4874 87068 5182 87077
rect 4874 87066 4880 87068
rect 4936 87066 4960 87068
rect 5016 87066 5040 87068
rect 5096 87066 5120 87068
rect 5176 87066 5182 87068
rect 4936 87014 4938 87066
rect 5118 87014 5120 87066
rect 4874 87012 4880 87014
rect 4936 87012 4960 87014
rect 5016 87012 5040 87014
rect 5096 87012 5120 87014
rect 5176 87012 5182 87014
rect 4874 87003 5182 87012
rect 4214 86524 4522 86533
rect 4214 86522 4220 86524
rect 4276 86522 4300 86524
rect 4356 86522 4380 86524
rect 4436 86522 4460 86524
rect 4516 86522 4522 86524
rect 4276 86470 4278 86522
rect 4458 86470 4460 86522
rect 4214 86468 4220 86470
rect 4276 86468 4300 86470
rect 4356 86468 4380 86470
rect 4436 86468 4460 86470
rect 4516 86468 4522 86470
rect 4214 86459 4522 86468
rect 4874 85980 5182 85989
rect 4874 85978 4880 85980
rect 4936 85978 4960 85980
rect 5016 85978 5040 85980
rect 5096 85978 5120 85980
rect 5176 85978 5182 85980
rect 4936 85926 4938 85978
rect 5118 85926 5120 85978
rect 4874 85924 4880 85926
rect 4936 85924 4960 85926
rect 5016 85924 5040 85926
rect 5096 85924 5120 85926
rect 5176 85924 5182 85926
rect 4874 85915 5182 85924
rect 4214 85436 4522 85445
rect 4214 85434 4220 85436
rect 4276 85434 4300 85436
rect 4356 85434 4380 85436
rect 4436 85434 4460 85436
rect 4516 85434 4522 85436
rect 4276 85382 4278 85434
rect 4458 85382 4460 85434
rect 4214 85380 4220 85382
rect 4276 85380 4300 85382
rect 4356 85380 4380 85382
rect 4436 85380 4460 85382
rect 4516 85380 4522 85382
rect 4214 85371 4522 85380
rect 4874 84892 5182 84901
rect 4874 84890 4880 84892
rect 4936 84890 4960 84892
rect 5016 84890 5040 84892
rect 5096 84890 5120 84892
rect 5176 84890 5182 84892
rect 4936 84838 4938 84890
rect 5118 84838 5120 84890
rect 4874 84836 4880 84838
rect 4936 84836 4960 84838
rect 5016 84836 5040 84838
rect 5096 84836 5120 84838
rect 5176 84836 5182 84838
rect 4874 84827 5182 84836
rect 4214 84348 4522 84357
rect 4214 84346 4220 84348
rect 4276 84346 4300 84348
rect 4356 84346 4380 84348
rect 4436 84346 4460 84348
rect 4516 84346 4522 84348
rect 4276 84294 4278 84346
rect 4458 84294 4460 84346
rect 4214 84292 4220 84294
rect 4276 84292 4300 84294
rect 4356 84292 4380 84294
rect 4436 84292 4460 84294
rect 4516 84292 4522 84294
rect 4214 84283 4522 84292
rect 4874 83804 5182 83813
rect 4874 83802 4880 83804
rect 4936 83802 4960 83804
rect 5016 83802 5040 83804
rect 5096 83802 5120 83804
rect 5176 83802 5182 83804
rect 4936 83750 4938 83802
rect 5118 83750 5120 83802
rect 4874 83748 4880 83750
rect 4936 83748 4960 83750
rect 5016 83748 5040 83750
rect 5096 83748 5120 83750
rect 5176 83748 5182 83750
rect 4874 83739 5182 83748
rect 4214 83260 4522 83269
rect 4214 83258 4220 83260
rect 4276 83258 4300 83260
rect 4356 83258 4380 83260
rect 4436 83258 4460 83260
rect 4516 83258 4522 83260
rect 4276 83206 4278 83258
rect 4458 83206 4460 83258
rect 4214 83204 4220 83206
rect 4276 83204 4300 83206
rect 4356 83204 4380 83206
rect 4436 83204 4460 83206
rect 4516 83204 4522 83206
rect 4214 83195 4522 83204
rect 4874 82716 5182 82725
rect 4874 82714 4880 82716
rect 4936 82714 4960 82716
rect 5016 82714 5040 82716
rect 5096 82714 5120 82716
rect 5176 82714 5182 82716
rect 4936 82662 4938 82714
rect 5118 82662 5120 82714
rect 4874 82660 4880 82662
rect 4936 82660 4960 82662
rect 5016 82660 5040 82662
rect 5096 82660 5120 82662
rect 5176 82660 5182 82662
rect 4874 82651 5182 82660
rect 4214 82172 4522 82181
rect 4214 82170 4220 82172
rect 4276 82170 4300 82172
rect 4356 82170 4380 82172
rect 4436 82170 4460 82172
rect 4516 82170 4522 82172
rect 4276 82118 4278 82170
rect 4458 82118 4460 82170
rect 4214 82116 4220 82118
rect 4276 82116 4300 82118
rect 4356 82116 4380 82118
rect 4436 82116 4460 82118
rect 4516 82116 4522 82118
rect 4214 82107 4522 82116
rect 4874 81628 5182 81637
rect 4874 81626 4880 81628
rect 4936 81626 4960 81628
rect 5016 81626 5040 81628
rect 5096 81626 5120 81628
rect 5176 81626 5182 81628
rect 4936 81574 4938 81626
rect 5118 81574 5120 81626
rect 4874 81572 4880 81574
rect 4936 81572 4960 81574
rect 5016 81572 5040 81574
rect 5096 81572 5120 81574
rect 5176 81572 5182 81574
rect 4874 81563 5182 81572
rect 4214 81084 4522 81093
rect 4214 81082 4220 81084
rect 4276 81082 4300 81084
rect 4356 81082 4380 81084
rect 4436 81082 4460 81084
rect 4516 81082 4522 81084
rect 4276 81030 4278 81082
rect 4458 81030 4460 81082
rect 4214 81028 4220 81030
rect 4276 81028 4300 81030
rect 4356 81028 4380 81030
rect 4436 81028 4460 81030
rect 4516 81028 4522 81030
rect 4214 81019 4522 81028
rect 4874 80540 5182 80549
rect 4874 80538 4880 80540
rect 4936 80538 4960 80540
rect 5016 80538 5040 80540
rect 5096 80538 5120 80540
rect 5176 80538 5182 80540
rect 4936 80486 4938 80538
rect 5118 80486 5120 80538
rect 4874 80484 4880 80486
rect 4936 80484 4960 80486
rect 5016 80484 5040 80486
rect 5096 80484 5120 80486
rect 5176 80484 5182 80486
rect 4874 80475 5182 80484
rect 4214 79996 4522 80005
rect 4214 79994 4220 79996
rect 4276 79994 4300 79996
rect 4356 79994 4380 79996
rect 4436 79994 4460 79996
rect 4516 79994 4522 79996
rect 4276 79942 4278 79994
rect 4458 79942 4460 79994
rect 4214 79940 4220 79942
rect 4276 79940 4300 79942
rect 4356 79940 4380 79942
rect 4436 79940 4460 79942
rect 4516 79940 4522 79942
rect 4214 79931 4522 79940
rect 4874 79452 5182 79461
rect 4874 79450 4880 79452
rect 4936 79450 4960 79452
rect 5016 79450 5040 79452
rect 5096 79450 5120 79452
rect 5176 79450 5182 79452
rect 4936 79398 4938 79450
rect 5118 79398 5120 79450
rect 4874 79396 4880 79398
rect 4936 79396 4960 79398
rect 5016 79396 5040 79398
rect 5096 79396 5120 79398
rect 5176 79396 5182 79398
rect 4874 79387 5182 79396
rect 4214 78908 4522 78917
rect 4214 78906 4220 78908
rect 4276 78906 4300 78908
rect 4356 78906 4380 78908
rect 4436 78906 4460 78908
rect 4516 78906 4522 78908
rect 4276 78854 4278 78906
rect 4458 78854 4460 78906
rect 4214 78852 4220 78854
rect 4276 78852 4300 78854
rect 4356 78852 4380 78854
rect 4436 78852 4460 78854
rect 4516 78852 4522 78854
rect 4214 78843 4522 78852
rect 4874 78364 5182 78373
rect 4874 78362 4880 78364
rect 4936 78362 4960 78364
rect 5016 78362 5040 78364
rect 5096 78362 5120 78364
rect 5176 78362 5182 78364
rect 4936 78310 4938 78362
rect 5118 78310 5120 78362
rect 4874 78308 4880 78310
rect 4936 78308 4960 78310
rect 5016 78308 5040 78310
rect 5096 78308 5120 78310
rect 5176 78308 5182 78310
rect 4874 78299 5182 78308
rect 4214 77820 4522 77829
rect 4214 77818 4220 77820
rect 4276 77818 4300 77820
rect 4356 77818 4380 77820
rect 4436 77818 4460 77820
rect 4516 77818 4522 77820
rect 4276 77766 4278 77818
rect 4458 77766 4460 77818
rect 4214 77764 4220 77766
rect 4276 77764 4300 77766
rect 4356 77764 4380 77766
rect 4436 77764 4460 77766
rect 4516 77764 4522 77766
rect 4214 77755 4522 77764
rect 4874 77276 5182 77285
rect 4874 77274 4880 77276
rect 4936 77274 4960 77276
rect 5016 77274 5040 77276
rect 5096 77274 5120 77276
rect 5176 77274 5182 77276
rect 4936 77222 4938 77274
rect 5118 77222 5120 77274
rect 4874 77220 4880 77222
rect 4936 77220 4960 77222
rect 5016 77220 5040 77222
rect 5096 77220 5120 77222
rect 5176 77220 5182 77222
rect 4874 77211 5182 77220
rect 4214 76732 4522 76741
rect 4214 76730 4220 76732
rect 4276 76730 4300 76732
rect 4356 76730 4380 76732
rect 4436 76730 4460 76732
rect 4516 76730 4522 76732
rect 4276 76678 4278 76730
rect 4458 76678 4460 76730
rect 4214 76676 4220 76678
rect 4276 76676 4300 76678
rect 4356 76676 4380 76678
rect 4436 76676 4460 76678
rect 4516 76676 4522 76678
rect 4214 76667 4522 76676
rect 4874 76188 5182 76197
rect 4874 76186 4880 76188
rect 4936 76186 4960 76188
rect 5016 76186 5040 76188
rect 5096 76186 5120 76188
rect 5176 76186 5182 76188
rect 4936 76134 4938 76186
rect 5118 76134 5120 76186
rect 4874 76132 4880 76134
rect 4936 76132 4960 76134
rect 5016 76132 5040 76134
rect 5096 76132 5120 76134
rect 5176 76132 5182 76134
rect 4874 76123 5182 76132
rect 4214 75644 4522 75653
rect 4214 75642 4220 75644
rect 4276 75642 4300 75644
rect 4356 75642 4380 75644
rect 4436 75642 4460 75644
rect 4516 75642 4522 75644
rect 4276 75590 4278 75642
rect 4458 75590 4460 75642
rect 4214 75588 4220 75590
rect 4276 75588 4300 75590
rect 4356 75588 4380 75590
rect 4436 75588 4460 75590
rect 4516 75588 4522 75590
rect 4214 75579 4522 75588
rect 4874 75100 5182 75109
rect 4874 75098 4880 75100
rect 4936 75098 4960 75100
rect 5016 75098 5040 75100
rect 5096 75098 5120 75100
rect 5176 75098 5182 75100
rect 4936 75046 4938 75098
rect 5118 75046 5120 75098
rect 4874 75044 4880 75046
rect 4936 75044 4960 75046
rect 5016 75044 5040 75046
rect 5096 75044 5120 75046
rect 5176 75044 5182 75046
rect 4874 75035 5182 75044
rect 4214 74556 4522 74565
rect 4214 74554 4220 74556
rect 4276 74554 4300 74556
rect 4356 74554 4380 74556
rect 4436 74554 4460 74556
rect 4516 74554 4522 74556
rect 4276 74502 4278 74554
rect 4458 74502 4460 74554
rect 4214 74500 4220 74502
rect 4276 74500 4300 74502
rect 4356 74500 4380 74502
rect 4436 74500 4460 74502
rect 4516 74500 4522 74502
rect 4214 74491 4522 74500
rect 4874 74012 5182 74021
rect 4874 74010 4880 74012
rect 4936 74010 4960 74012
rect 5016 74010 5040 74012
rect 5096 74010 5120 74012
rect 5176 74010 5182 74012
rect 4936 73958 4938 74010
rect 5118 73958 5120 74010
rect 4874 73956 4880 73958
rect 4936 73956 4960 73958
rect 5016 73956 5040 73958
rect 5096 73956 5120 73958
rect 5176 73956 5182 73958
rect 4874 73947 5182 73956
rect 4214 73468 4522 73477
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73403 4522 73412
rect 4874 72924 5182 72933
rect 4874 72922 4880 72924
rect 4936 72922 4960 72924
rect 5016 72922 5040 72924
rect 5096 72922 5120 72924
rect 5176 72922 5182 72924
rect 4936 72870 4938 72922
rect 5118 72870 5120 72922
rect 4874 72868 4880 72870
rect 4936 72868 4960 72870
rect 5016 72868 5040 72870
rect 5096 72868 5120 72870
rect 5176 72868 5182 72870
rect 4874 72859 5182 72868
rect 4214 72380 4522 72389
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 4214 72315 4522 72324
rect 4874 71836 5182 71845
rect 4874 71834 4880 71836
rect 4936 71834 4960 71836
rect 5016 71834 5040 71836
rect 5096 71834 5120 71836
rect 5176 71834 5182 71836
rect 4936 71782 4938 71834
rect 5118 71782 5120 71834
rect 4874 71780 4880 71782
rect 4936 71780 4960 71782
rect 5016 71780 5040 71782
rect 5096 71780 5120 71782
rect 5176 71780 5182 71782
rect 4874 71771 5182 71780
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 4874 70748 5182 70757
rect 4874 70746 4880 70748
rect 4936 70746 4960 70748
rect 5016 70746 5040 70748
rect 5096 70746 5120 70748
rect 5176 70746 5182 70748
rect 4936 70694 4938 70746
rect 5118 70694 5120 70746
rect 4874 70692 4880 70694
rect 4936 70692 4960 70694
rect 5016 70692 5040 70694
rect 5096 70692 5120 70694
rect 5176 70692 5182 70694
rect 4874 70683 5182 70692
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70139 4522 70148
rect 4874 69660 5182 69669
rect 4874 69658 4880 69660
rect 4936 69658 4960 69660
rect 5016 69658 5040 69660
rect 5096 69658 5120 69660
rect 5176 69658 5182 69660
rect 4936 69606 4938 69658
rect 5118 69606 5120 69658
rect 4874 69604 4880 69606
rect 4936 69604 4960 69606
rect 5016 69604 5040 69606
rect 5096 69604 5120 69606
rect 5176 69604 5182 69606
rect 4874 69595 5182 69604
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 4874 68572 5182 68581
rect 4874 68570 4880 68572
rect 4936 68570 4960 68572
rect 5016 68570 5040 68572
rect 5096 68570 5120 68572
rect 5176 68570 5182 68572
rect 4936 68518 4938 68570
rect 5118 68518 5120 68570
rect 4874 68516 4880 68518
rect 4936 68516 4960 68518
rect 5016 68516 5040 68518
rect 5096 68516 5120 68518
rect 5176 68516 5182 68518
rect 4874 68507 5182 68516
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 4874 67484 5182 67493
rect 4874 67482 4880 67484
rect 4936 67482 4960 67484
rect 5016 67482 5040 67484
rect 5096 67482 5120 67484
rect 5176 67482 5182 67484
rect 4936 67430 4938 67482
rect 5118 67430 5120 67482
rect 4874 67428 4880 67430
rect 4936 67428 4960 67430
rect 5016 67428 5040 67430
rect 5096 67428 5120 67430
rect 5176 67428 5182 67430
rect 4874 67419 5182 67428
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 4874 66396 5182 66405
rect 4874 66394 4880 66396
rect 4936 66394 4960 66396
rect 5016 66394 5040 66396
rect 5096 66394 5120 66396
rect 5176 66394 5182 66396
rect 4936 66342 4938 66394
rect 5118 66342 5120 66394
rect 4874 66340 4880 66342
rect 4936 66340 4960 66342
rect 5016 66340 5040 66342
rect 5096 66340 5120 66342
rect 5176 66340 5182 66342
rect 4874 66331 5182 66340
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 4874 65308 5182 65317
rect 4874 65306 4880 65308
rect 4936 65306 4960 65308
rect 5016 65306 5040 65308
rect 5096 65306 5120 65308
rect 5176 65306 5182 65308
rect 4936 65254 4938 65306
rect 5118 65254 5120 65306
rect 4874 65252 4880 65254
rect 4936 65252 4960 65254
rect 5016 65252 5040 65254
rect 5096 65252 5120 65254
rect 5176 65252 5182 65254
rect 4874 65243 5182 65252
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 4874 64220 5182 64229
rect 4874 64218 4880 64220
rect 4936 64218 4960 64220
rect 5016 64218 5040 64220
rect 5096 64218 5120 64220
rect 5176 64218 5182 64220
rect 4936 64166 4938 64218
rect 5118 64166 5120 64218
rect 4874 64164 4880 64166
rect 4936 64164 4960 64166
rect 5016 64164 5040 64166
rect 5096 64164 5120 64166
rect 5176 64164 5182 64166
rect 4874 64155 5182 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 4874 63132 5182 63141
rect 4874 63130 4880 63132
rect 4936 63130 4960 63132
rect 5016 63130 5040 63132
rect 5096 63130 5120 63132
rect 5176 63130 5182 63132
rect 4936 63078 4938 63130
rect 5118 63078 5120 63130
rect 4874 63076 4880 63078
rect 4936 63076 4960 63078
rect 5016 63076 5040 63078
rect 5096 63076 5120 63078
rect 5176 63076 5182 63078
rect 4874 63067 5182 63076
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 4874 62044 5182 62053
rect 4874 62042 4880 62044
rect 4936 62042 4960 62044
rect 5016 62042 5040 62044
rect 5096 62042 5120 62044
rect 5176 62042 5182 62044
rect 4936 61990 4938 62042
rect 5118 61990 5120 62042
rect 4874 61988 4880 61990
rect 4936 61988 4960 61990
rect 5016 61988 5040 61990
rect 5096 61988 5120 61990
rect 5176 61988 5182 61990
rect 4874 61979 5182 61988
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4874 60956 5182 60965
rect 4874 60954 4880 60956
rect 4936 60954 4960 60956
rect 5016 60954 5040 60956
rect 5096 60954 5120 60956
rect 5176 60954 5182 60956
rect 4936 60902 4938 60954
rect 5118 60902 5120 60954
rect 4874 60900 4880 60902
rect 4936 60900 4960 60902
rect 5016 60900 5040 60902
rect 5096 60900 5120 60902
rect 5176 60900 5182 60902
rect 4874 60891 5182 60900
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 4874 59868 5182 59877
rect 4874 59866 4880 59868
rect 4936 59866 4960 59868
rect 5016 59866 5040 59868
rect 5096 59866 5120 59868
rect 5176 59866 5182 59868
rect 4936 59814 4938 59866
rect 5118 59814 5120 59866
rect 4874 59812 4880 59814
rect 4936 59812 4960 59814
rect 5016 59812 5040 59814
rect 5096 59812 5120 59814
rect 5176 59812 5182 59814
rect 4874 59803 5182 59812
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4874 58780 5182 58789
rect 4874 58778 4880 58780
rect 4936 58778 4960 58780
rect 5016 58778 5040 58780
rect 5096 58778 5120 58780
rect 5176 58778 5182 58780
rect 4936 58726 4938 58778
rect 5118 58726 5120 58778
rect 4874 58724 4880 58726
rect 4936 58724 4960 58726
rect 5016 58724 5040 58726
rect 5096 58724 5120 58726
rect 5176 58724 5182 58726
rect 4874 58715 5182 58724
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 1308 44396 1360 44402
rect 1308 44338 1360 44344
rect 1320 44305 1348 44338
rect 1306 44296 1362 44305
rect 1306 44231 1362 44240
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 1308 43308 1360 43314
rect 1308 43250 1360 43256
rect 1320 42945 1348 43250
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 1306 42936 1362 42945
rect 4214 42939 4522 42948
rect 1306 42871 1362 42880
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 1308 41132 1360 41138
rect 1308 41074 1360 41080
rect 1320 40905 1348 41074
rect 1306 40896 1362 40905
rect 1306 40831 1362 40840
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 1308 40520 1360 40526
rect 1308 40462 1360 40468
rect 1320 40225 1348 40462
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 1306 40216 1362 40225
rect 4874 40219 5182 40228
rect 1306 40151 1362 40160
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 1216 38344 1268 38350
rect 1216 38286 1268 38292
rect 1228 38185 1256 38286
rect 1214 38176 1270 38185
rect 1214 38111 1270 38120
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 1308 37868 1360 37874
rect 1308 37810 1360 37816
rect 1320 37505 1348 37810
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 1306 37496 1362 37505
rect 4214 37499 4522 37508
rect 1306 37431 1362 37440
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 1308 35692 1360 35698
rect 1308 35634 1360 35640
rect 1320 35465 1348 35634
rect 1306 35456 1362 35465
rect 1306 35391 1362 35400
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 1320 15745 1348 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 1306 15736 1362 15745
rect 4214 15739 4522 15748
rect 1306 15671 1362 15680
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 8220 9654 8248 92006
rect 34934 91964 35242 91973
rect 34934 91962 34940 91964
rect 34996 91962 35020 91964
rect 35076 91962 35100 91964
rect 35156 91962 35180 91964
rect 35236 91962 35242 91964
rect 34996 91910 34998 91962
rect 35178 91910 35180 91962
rect 34934 91908 34940 91910
rect 34996 91908 35020 91910
rect 35076 91908 35100 91910
rect 35156 91908 35180 91910
rect 35236 91908 35242 91910
rect 34934 91899 35242 91908
rect 46860 89729 46888 92006
rect 49620 91866 49648 92006
rect 54852 92006 54904 92012
rect 53194 91967 53250 91976
rect 55232 91866 55260 94726
rect 55692 94450 55720 95406
rect 55496 94444 55548 94450
rect 55496 94386 55548 94392
rect 55680 94444 55732 94450
rect 55680 94386 55732 94392
rect 55864 94444 55916 94450
rect 55864 94386 55916 94392
rect 55404 94376 55456 94382
rect 55404 94318 55456 94324
rect 55416 92954 55444 94318
rect 55508 93838 55536 94386
rect 55876 94246 55904 94386
rect 55588 94240 55640 94246
rect 55588 94182 55640 94188
rect 55864 94240 55916 94246
rect 55864 94182 55916 94188
rect 55600 93974 55628 94182
rect 55588 93968 55640 93974
rect 55586 93936 55588 93945
rect 55640 93936 55642 93945
rect 55586 93871 55642 93880
rect 55496 93832 55548 93838
rect 55496 93774 55548 93780
rect 56508 93832 56560 93838
rect 56508 93774 56560 93780
rect 55772 93696 55824 93702
rect 55772 93638 55824 93644
rect 55784 93430 55812 93638
rect 55772 93424 55824 93430
rect 55772 93366 55824 93372
rect 56232 93424 56284 93430
rect 56232 93366 56284 93372
rect 56244 93158 56272 93366
rect 56520 93294 56548 93774
rect 56612 93362 56640 96970
rect 56784 96688 56836 96694
rect 56784 96630 56836 96636
rect 56796 96082 56824 96630
rect 56784 96076 56836 96082
rect 56784 96018 56836 96024
rect 56796 94994 56824 96018
rect 57060 95940 57112 95946
rect 57060 95882 57112 95888
rect 56784 94988 56836 94994
rect 56784 94930 56836 94936
rect 56876 94920 56928 94926
rect 56876 94862 56928 94868
rect 56888 94382 56916 94862
rect 57072 94586 57100 95882
rect 57440 95674 57468 97038
rect 58176 96218 58204 97038
rect 58164 96212 58216 96218
rect 58164 96154 58216 96160
rect 59176 95940 59228 95946
rect 59176 95882 59228 95888
rect 57428 95668 57480 95674
rect 57428 95610 57480 95616
rect 57704 95600 57756 95606
rect 57704 95542 57756 95548
rect 57612 95532 57664 95538
rect 57612 95474 57664 95480
rect 57060 94580 57112 94586
rect 57060 94522 57112 94528
rect 56876 94376 56928 94382
rect 56876 94318 56928 94324
rect 56600 93356 56652 93362
rect 56600 93298 56652 93304
rect 56324 93288 56376 93294
rect 56324 93230 56376 93236
rect 56508 93288 56560 93294
rect 56508 93230 56560 93236
rect 56336 93158 56364 93230
rect 56232 93152 56284 93158
rect 56232 93094 56284 93100
rect 56324 93152 56376 93158
rect 56324 93094 56376 93100
rect 55404 92948 55456 92954
rect 55404 92890 55456 92896
rect 56520 92750 56548 93230
rect 56508 92744 56560 92750
rect 56508 92686 56560 92692
rect 56048 92336 56100 92342
rect 56520 92290 56548 92686
rect 56612 92585 56640 93298
rect 56888 93294 56916 94318
rect 57624 93498 57652 95474
rect 57716 94518 57744 95542
rect 57888 95464 57940 95470
rect 57888 95406 57940 95412
rect 57900 94994 57928 95406
rect 57888 94988 57940 94994
rect 57888 94930 57940 94936
rect 57796 94852 57848 94858
rect 57796 94794 57848 94800
rect 57704 94512 57756 94518
rect 57704 94454 57756 94460
rect 57808 94042 57836 94794
rect 58440 94444 58492 94450
rect 58440 94386 58492 94392
rect 57888 94376 57940 94382
rect 57888 94318 57940 94324
rect 57900 94042 57928 94318
rect 57796 94036 57848 94042
rect 57796 93978 57848 93984
rect 57888 94036 57940 94042
rect 57888 93978 57940 93984
rect 58452 93854 58480 94386
rect 58360 93826 58480 93854
rect 59188 93854 59216 95882
rect 59280 95130 59308 97038
rect 59544 95328 59596 95334
rect 59544 95270 59596 95276
rect 59268 95124 59320 95130
rect 59268 95066 59320 95072
rect 59556 94450 59584 95270
rect 60568 94586 60596 97038
rect 60936 95674 60964 97038
rect 62868 95674 62896 97038
rect 60924 95668 60976 95674
rect 60924 95610 60976 95616
rect 62764 95668 62816 95674
rect 62764 95610 62816 95616
rect 62856 95668 62908 95674
rect 62856 95610 62908 95616
rect 60740 95396 60792 95402
rect 60740 95338 60792 95344
rect 60004 94580 60056 94586
rect 60004 94522 60056 94528
rect 60556 94580 60608 94586
rect 60556 94522 60608 94528
rect 59544 94444 59596 94450
rect 59544 94386 59596 94392
rect 59188 93826 59308 93854
rect 59556 93838 59584 94386
rect 58164 93764 58216 93770
rect 58164 93706 58216 93712
rect 57612 93492 57664 93498
rect 57612 93434 57664 93440
rect 56876 93288 56928 93294
rect 56876 93230 56928 93236
rect 57978 92848 58034 92857
rect 57978 92783 57980 92792
rect 58032 92783 58034 92792
rect 57980 92754 58032 92760
rect 56598 92576 56654 92585
rect 56598 92511 56654 92520
rect 56048 92278 56100 92284
rect 56060 91866 56088 92278
rect 56428 92274 56548 92290
rect 56416 92268 56548 92274
rect 56468 92262 56548 92268
rect 56416 92210 56468 92216
rect 49608 91860 49660 91866
rect 49608 91802 49660 91808
rect 55220 91860 55272 91866
rect 55220 91802 55272 91808
rect 56048 91860 56100 91866
rect 56048 91802 56100 91808
rect 58176 90001 58204 93706
rect 58360 92410 58388 93826
rect 59280 93770 59308 93826
rect 59544 93832 59596 93838
rect 59544 93774 59596 93780
rect 59636 93832 59688 93838
rect 59636 93774 59688 93780
rect 59268 93764 59320 93770
rect 59268 93706 59320 93712
rect 59360 93696 59412 93702
rect 59360 93638 59412 93644
rect 58900 93424 58952 93430
rect 58900 93366 58952 93372
rect 58438 92848 58494 92857
rect 58438 92783 58494 92792
rect 58452 92682 58480 92783
rect 58912 92750 58940 93366
rect 58900 92744 58952 92750
rect 58900 92686 58952 92692
rect 58440 92676 58492 92682
rect 58440 92618 58492 92624
rect 58348 92404 58400 92410
rect 58348 92346 58400 92352
rect 58912 92274 58940 92686
rect 59268 92676 59320 92682
rect 59268 92618 59320 92624
rect 58900 92268 58952 92274
rect 58900 92210 58952 92216
rect 58714 92168 58770 92177
rect 58714 92103 58716 92112
rect 58768 92103 58770 92112
rect 58716 92074 58768 92080
rect 58162 89992 58218 90001
rect 58162 89927 58218 89936
rect 59280 89865 59308 92618
rect 59266 89856 59322 89865
rect 59266 89791 59322 89800
rect 59372 89729 59400 93638
rect 59556 93430 59584 93774
rect 59648 93498 59676 93774
rect 60016 93498 60044 94522
rect 60096 94512 60148 94518
rect 60096 94454 60148 94460
rect 60108 94364 60136 94454
rect 60188 94376 60240 94382
rect 60108 94336 60188 94364
rect 60108 93838 60136 94336
rect 60188 94318 60240 94324
rect 60752 94042 60780 95338
rect 62028 95328 62080 95334
rect 62028 95270 62080 95276
rect 62040 94994 62068 95270
rect 62028 94988 62080 94994
rect 62028 94930 62080 94936
rect 61752 94852 61804 94858
rect 61752 94794 61804 94800
rect 62304 94852 62356 94858
rect 62304 94794 62356 94800
rect 61764 94586 61792 94794
rect 61752 94580 61804 94586
rect 61752 94522 61804 94528
rect 60740 94036 60792 94042
rect 60740 93978 60792 93984
rect 60096 93832 60148 93838
rect 60096 93774 60148 93780
rect 61476 93832 61528 93838
rect 61476 93774 61528 93780
rect 61660 93832 61712 93838
rect 61660 93774 61712 93780
rect 60372 93764 60424 93770
rect 60372 93706 60424 93712
rect 59636 93492 59688 93498
rect 59636 93434 59688 93440
rect 60004 93492 60056 93498
rect 60004 93434 60056 93440
rect 59544 93424 59596 93430
rect 59544 93366 59596 93372
rect 59820 93356 59872 93362
rect 59820 93298 59872 93304
rect 59832 92721 59860 93298
rect 60384 93158 60412 93706
rect 60648 93696 60700 93702
rect 60648 93638 60700 93644
rect 61384 93696 61436 93702
rect 61384 93638 61436 93644
rect 60660 93498 60688 93638
rect 60648 93492 60700 93498
rect 60648 93434 60700 93440
rect 60740 93424 60792 93430
rect 60740 93366 60792 93372
rect 60372 93152 60424 93158
rect 60372 93094 60424 93100
rect 60464 93152 60516 93158
rect 60464 93094 60516 93100
rect 60476 92886 60504 93094
rect 60464 92880 60516 92886
rect 60464 92822 60516 92828
rect 59818 92712 59874 92721
rect 59818 92647 59874 92656
rect 59452 92608 59504 92614
rect 59452 92550 59504 92556
rect 59464 90001 59492 92550
rect 60752 92274 60780 93366
rect 61396 92954 61424 93638
rect 61488 93480 61516 93774
rect 61568 93492 61620 93498
rect 61488 93452 61568 93480
rect 61568 93434 61620 93440
rect 61672 93158 61700 93774
rect 62316 93770 62344 94794
rect 62776 93838 62804 95610
rect 63512 95130 63540 97038
rect 64984 95674 65012 97038
rect 64880 95668 64932 95674
rect 64880 95610 64932 95616
rect 64972 95668 65024 95674
rect 64972 95610 65024 95616
rect 63592 95464 63644 95470
rect 63592 95406 63644 95412
rect 63500 95124 63552 95130
rect 63500 95066 63552 95072
rect 63224 94512 63276 94518
rect 63224 94454 63276 94460
rect 62764 93832 62816 93838
rect 62764 93774 62816 93780
rect 62304 93764 62356 93770
rect 62304 93706 62356 93712
rect 61752 93696 61804 93702
rect 61752 93638 61804 93644
rect 62856 93696 62908 93702
rect 62908 93656 62988 93684
rect 62856 93638 62908 93644
rect 61660 93152 61712 93158
rect 61660 93094 61712 93100
rect 61292 92948 61344 92954
rect 61292 92890 61344 92896
rect 61384 92948 61436 92954
rect 61384 92890 61436 92896
rect 61304 92614 61332 92890
rect 61292 92608 61344 92614
rect 61292 92550 61344 92556
rect 60740 92268 60792 92274
rect 60740 92210 60792 92216
rect 60556 92132 60608 92138
rect 60556 92074 60608 92080
rect 59450 89992 59506 90001
rect 59450 89927 59506 89936
rect 46846 89720 46902 89729
rect 46846 89655 46902 89664
rect 59358 89720 59414 89729
rect 59358 89655 59414 89664
rect 60568 89593 60596 92074
rect 61764 91866 61792 93638
rect 62856 93152 62908 93158
rect 62856 93094 62908 93100
rect 61752 91860 61804 91866
rect 61752 91802 61804 91808
rect 62868 91089 62896 93094
rect 62960 92886 62988 93656
rect 63236 93362 63264 94454
rect 63316 94376 63368 94382
rect 63604 94330 63632 95406
rect 64788 95396 64840 95402
rect 64788 95338 64840 95344
rect 64144 94784 64196 94790
rect 64144 94726 64196 94732
rect 63316 94318 63368 94324
rect 63328 93838 63356 94318
rect 63512 94302 63632 94330
rect 63776 94308 63828 94314
rect 63316 93832 63368 93838
rect 63316 93774 63368 93780
rect 63328 93362 63356 93774
rect 63512 93770 63540 94302
rect 63776 94250 63828 94256
rect 63592 94240 63644 94246
rect 63592 94182 63644 94188
rect 63604 93906 63632 94182
rect 63592 93900 63644 93906
rect 63592 93842 63644 93848
rect 63788 93838 63816 94250
rect 64156 94042 64184 94726
rect 64144 94036 64196 94042
rect 64144 93978 64196 93984
rect 63776 93832 63828 93838
rect 63776 93774 63828 93780
rect 64696 93832 64748 93838
rect 64696 93774 64748 93780
rect 63500 93764 63552 93770
rect 63500 93706 63552 93712
rect 64512 93696 64564 93702
rect 64512 93638 64564 93644
rect 64604 93696 64656 93702
rect 64604 93638 64656 93644
rect 63500 93492 63552 93498
rect 63500 93434 63552 93440
rect 63224 93356 63276 93362
rect 63224 93298 63276 93304
rect 63316 93356 63368 93362
rect 63316 93298 63368 93304
rect 63512 93242 63540 93434
rect 63592 93424 63644 93430
rect 63592 93366 63644 93372
rect 63328 93214 63540 93242
rect 62948 92880 63000 92886
rect 62948 92822 63000 92828
rect 63224 92676 63276 92682
rect 63328 92664 63356 93214
rect 63408 93152 63460 93158
rect 63408 93094 63460 93100
rect 63420 92954 63448 93094
rect 63498 92984 63554 92993
rect 63408 92948 63460 92954
rect 63498 92919 63500 92928
rect 63408 92890 63460 92896
rect 63552 92919 63554 92928
rect 63500 92890 63552 92896
rect 63512 92682 63540 92890
rect 63604 92818 63632 93366
rect 63776 93288 63828 93294
rect 63776 93230 63828 93236
rect 63592 92812 63644 92818
rect 63592 92754 63644 92760
rect 63276 92636 63356 92664
rect 63500 92676 63552 92682
rect 63224 92618 63276 92624
rect 63500 92618 63552 92624
rect 63788 92585 63816 93230
rect 64524 92868 64552 93638
rect 64616 92970 64644 93638
rect 64708 93242 64736 93774
rect 64800 93770 64828 95338
rect 64892 93838 64920 95610
rect 65064 95464 65116 95470
rect 65064 95406 65116 95412
rect 65076 94994 65104 95406
rect 65064 94988 65116 94994
rect 65064 94930 65116 94936
rect 65248 94852 65300 94858
rect 65248 94794 65300 94800
rect 65260 94586 65288 94794
rect 65248 94580 65300 94586
rect 65248 94522 65300 94528
rect 64880 93832 64932 93838
rect 64880 93774 64932 93780
rect 64788 93764 64840 93770
rect 64788 93706 64840 93712
rect 65248 93288 65300 93294
rect 64878 93256 64934 93265
rect 64708 93226 64828 93242
rect 64708 93220 64840 93226
rect 64708 93214 64788 93220
rect 65248 93230 65300 93236
rect 64878 93191 64934 93200
rect 64788 93162 64840 93168
rect 64616 92942 64736 92970
rect 64604 92880 64656 92886
rect 64524 92840 64604 92868
rect 64604 92822 64656 92828
rect 63498 92576 63554 92585
rect 63498 92511 63554 92520
rect 63774 92576 63830 92585
rect 63774 92511 63830 92520
rect 63512 92410 63540 92511
rect 63500 92404 63552 92410
rect 63500 92346 63552 92352
rect 64708 92070 64736 92942
rect 64892 92614 64920 93191
rect 64880 92608 64932 92614
rect 64880 92550 64932 92556
rect 64696 92064 64748 92070
rect 64696 92006 64748 92012
rect 62854 91080 62910 91089
rect 62854 91015 62910 91024
rect 65260 89729 65288 93230
rect 65352 92410 65380 97242
rect 67192 97238 67220 99334
rect 67638 99334 67864 99362
rect 67638 99200 67694 99334
rect 67836 97238 67864 99334
rect 68848 99334 68982 99362
rect 67180 97232 67232 97238
rect 67180 97174 67232 97180
rect 67824 97232 67876 97238
rect 67824 97174 67876 97180
rect 67640 97164 67692 97170
rect 67640 97106 67692 97112
rect 66720 97096 66772 97102
rect 66720 97038 66772 97044
rect 67364 97096 67416 97102
rect 67364 97038 67416 97044
rect 66314 96860 66622 96869
rect 66314 96858 66320 96860
rect 66376 96858 66400 96860
rect 66456 96858 66480 96860
rect 66536 96858 66560 96860
rect 66616 96858 66622 96860
rect 66376 96806 66378 96858
rect 66558 96806 66560 96858
rect 66314 96804 66320 96806
rect 66376 96804 66400 96806
rect 66456 96804 66480 96806
rect 66536 96804 66560 96806
rect 66616 96804 66622 96806
rect 66314 96795 66622 96804
rect 65654 96316 65962 96325
rect 65654 96314 65660 96316
rect 65716 96314 65740 96316
rect 65796 96314 65820 96316
rect 65876 96314 65900 96316
rect 65956 96314 65962 96316
rect 65716 96262 65718 96314
rect 65898 96262 65900 96314
rect 65654 96260 65660 96262
rect 65716 96260 65740 96262
rect 65796 96260 65820 96262
rect 65876 96260 65900 96262
rect 65956 96260 65962 96262
rect 65654 96251 65962 96260
rect 66314 95772 66622 95781
rect 66314 95770 66320 95772
rect 66376 95770 66400 95772
rect 66456 95770 66480 95772
rect 66536 95770 66560 95772
rect 66616 95770 66622 95772
rect 66376 95718 66378 95770
rect 66558 95718 66560 95770
rect 66314 95716 66320 95718
rect 66376 95716 66400 95718
rect 66456 95716 66480 95718
rect 66536 95716 66560 95718
rect 66616 95716 66622 95718
rect 66314 95707 66622 95716
rect 66732 95674 66760 97038
rect 66996 95872 67048 95878
rect 66996 95814 67048 95820
rect 66628 95668 66680 95674
rect 66628 95610 66680 95616
rect 66720 95668 66772 95674
rect 66720 95610 66772 95616
rect 65654 95228 65962 95237
rect 65654 95226 65660 95228
rect 65716 95226 65740 95228
rect 65796 95226 65820 95228
rect 65876 95226 65900 95228
rect 65956 95226 65962 95228
rect 65716 95174 65718 95226
rect 65898 95174 65900 95226
rect 65654 95172 65660 95174
rect 65716 95172 65740 95174
rect 65796 95172 65820 95174
rect 65876 95172 65900 95174
rect 65956 95172 65962 95174
rect 65654 95163 65962 95172
rect 66640 94874 66668 95610
rect 67008 95146 67036 95814
rect 67088 95600 67140 95606
rect 67088 95542 67140 95548
rect 66824 95118 67036 95146
rect 66640 94846 66760 94874
rect 66314 94684 66622 94693
rect 66314 94682 66320 94684
rect 66376 94682 66400 94684
rect 66456 94682 66480 94684
rect 66536 94682 66560 94684
rect 66616 94682 66622 94684
rect 66376 94630 66378 94682
rect 66558 94630 66560 94682
rect 66314 94628 66320 94630
rect 66376 94628 66400 94630
rect 66456 94628 66480 94630
rect 66536 94628 66560 94630
rect 66616 94628 66622 94630
rect 66314 94619 66622 94628
rect 65432 94444 65484 94450
rect 65432 94386 65484 94392
rect 65444 93974 65472 94386
rect 65654 94140 65962 94149
rect 65654 94138 65660 94140
rect 65716 94138 65740 94140
rect 65796 94138 65820 94140
rect 65876 94138 65900 94140
rect 65956 94138 65962 94140
rect 65716 94086 65718 94138
rect 65898 94086 65900 94138
rect 65654 94084 65660 94086
rect 65716 94084 65740 94086
rect 65796 94084 65820 94086
rect 65876 94084 65900 94086
rect 65956 94084 65962 94086
rect 65654 94075 65962 94084
rect 65432 93968 65484 93974
rect 65432 93910 65484 93916
rect 65444 93838 65472 93910
rect 66168 93900 66220 93906
rect 66168 93842 66220 93848
rect 65432 93832 65484 93838
rect 65892 93832 65944 93838
rect 65432 93774 65484 93780
rect 65890 93800 65892 93809
rect 65944 93800 65946 93809
rect 65890 93735 65946 93744
rect 65984 93696 66036 93702
rect 65984 93638 66036 93644
rect 65996 93498 66024 93638
rect 65984 93492 66036 93498
rect 65984 93434 66036 93440
rect 66180 93378 66208 93842
rect 66732 93702 66760 94846
rect 66824 93770 66852 95118
rect 66904 94988 66956 94994
rect 66904 94930 66956 94936
rect 66812 93764 66864 93770
rect 66812 93706 66864 93712
rect 66720 93696 66772 93702
rect 66720 93638 66772 93644
rect 66314 93596 66622 93605
rect 66314 93594 66320 93596
rect 66376 93594 66400 93596
rect 66456 93594 66480 93596
rect 66536 93594 66560 93596
rect 66616 93594 66622 93596
rect 66376 93542 66378 93594
rect 66558 93542 66560 93594
rect 66314 93540 66320 93542
rect 66376 93540 66400 93542
rect 66456 93540 66480 93542
rect 66536 93540 66560 93542
rect 66616 93540 66622 93542
rect 66314 93531 66622 93540
rect 66916 93430 66944 94930
rect 66996 94920 67048 94926
rect 66996 94862 67048 94868
rect 67008 93702 67036 94862
rect 67100 93838 67128 95542
rect 67376 95130 67404 97038
rect 67456 97028 67508 97034
rect 67456 96970 67508 96976
rect 67468 96150 67496 96970
rect 67652 96966 67680 97106
rect 68008 97096 68060 97102
rect 68008 97038 68060 97044
rect 67640 96960 67692 96966
rect 67640 96902 67692 96908
rect 67456 96144 67508 96150
rect 67456 96086 67508 96092
rect 67364 95124 67416 95130
rect 67364 95066 67416 95072
rect 67468 94994 67496 96086
rect 67456 94988 67508 94994
rect 67456 94930 67508 94936
rect 67180 94852 67232 94858
rect 67180 94794 67232 94800
rect 67192 94042 67220 94794
rect 67180 94036 67232 94042
rect 67180 93978 67232 93984
rect 67088 93832 67140 93838
rect 67088 93774 67140 93780
rect 67270 93800 67326 93809
rect 67270 93735 67272 93744
rect 67324 93735 67326 93744
rect 67272 93706 67324 93712
rect 66996 93696 67048 93702
rect 66996 93638 67048 93644
rect 66904 93424 66956 93430
rect 66180 93362 66392 93378
rect 66904 93366 66956 93372
rect 66180 93356 66404 93362
rect 66180 93350 66352 93356
rect 66352 93298 66404 93304
rect 66720 93356 66772 93362
rect 66720 93298 66772 93304
rect 65654 93052 65962 93061
rect 65654 93050 65660 93052
rect 65716 93050 65740 93052
rect 65796 93050 65820 93052
rect 65876 93050 65900 93052
rect 65956 93050 65962 93052
rect 65716 92998 65718 93050
rect 65898 92998 65900 93050
rect 65654 92996 65660 92998
rect 65716 92996 65740 92998
rect 65796 92996 65820 92998
rect 65876 92996 65900 92998
rect 65956 92996 65962 92998
rect 65654 92987 65962 92996
rect 66314 92508 66622 92517
rect 66314 92506 66320 92508
rect 66376 92506 66400 92508
rect 66456 92506 66480 92508
rect 66536 92506 66560 92508
rect 66616 92506 66622 92508
rect 66376 92454 66378 92506
rect 66558 92454 66560 92506
rect 66314 92452 66320 92454
rect 66376 92452 66400 92454
rect 66456 92452 66480 92454
rect 66536 92452 66560 92454
rect 66616 92452 66622 92454
rect 66314 92443 66622 92452
rect 65340 92404 65392 92410
rect 65340 92346 65392 92352
rect 66732 92206 66760 93298
rect 66812 93220 66864 93226
rect 66812 93162 66864 93168
rect 66720 92200 66772 92206
rect 66720 92142 66772 92148
rect 65654 91964 65962 91973
rect 65654 91962 65660 91964
rect 65716 91962 65740 91964
rect 65796 91962 65820 91964
rect 65876 91962 65900 91964
rect 65956 91962 65962 91964
rect 65716 91910 65718 91962
rect 65898 91910 65900 91962
rect 65654 91908 65660 91910
rect 65716 91908 65740 91910
rect 65796 91908 65820 91910
rect 65876 91908 65900 91910
rect 65956 91908 65962 91910
rect 65654 91899 65962 91908
rect 66824 89729 66852 93162
rect 67548 92676 67600 92682
rect 67548 92618 67600 92624
rect 67560 89729 67588 92618
rect 67652 92410 67680 96902
rect 68020 96218 68048 97038
rect 68848 96490 68876 99334
rect 68926 99200 68982 99334
rect 70214 99362 70270 100000
rect 71502 99362 71558 100000
rect 72146 99362 72202 100000
rect 74078 99362 74134 100000
rect 107566 99362 107622 100000
rect 108210 99362 108266 100000
rect 70214 99334 70348 99362
rect 70214 99200 70270 99334
rect 70320 97238 70348 99334
rect 71502 99334 71728 99362
rect 71502 99200 71558 99334
rect 71700 97238 71728 99334
rect 72146 99334 72372 99362
rect 72146 99200 72202 99334
rect 72344 97238 72372 99334
rect 74078 99334 74396 99362
rect 74078 99200 74134 99334
rect 74368 97238 74396 99334
rect 107488 99334 107622 99362
rect 96374 97404 96682 97413
rect 96374 97402 96380 97404
rect 96436 97402 96460 97404
rect 96516 97402 96540 97404
rect 96596 97402 96620 97404
rect 96676 97402 96682 97404
rect 96436 97350 96438 97402
rect 96618 97350 96620 97402
rect 96374 97348 96380 97350
rect 96436 97348 96460 97350
rect 96516 97348 96540 97350
rect 96596 97348 96620 97350
rect 96676 97348 96682 97350
rect 96374 97339 96682 97348
rect 107488 97238 107516 99334
rect 107566 99200 107622 99334
rect 107856 99334 108266 99362
rect 107856 97306 107884 99334
rect 108210 99200 108266 99334
rect 107844 97300 107896 97306
rect 107844 97242 107896 97248
rect 70308 97232 70360 97238
rect 70308 97174 70360 97180
rect 71688 97232 71740 97238
rect 71688 97174 71740 97180
rect 72332 97232 72384 97238
rect 72332 97174 72384 97180
rect 74356 97232 74408 97238
rect 74356 97174 74408 97180
rect 107476 97232 107528 97238
rect 107476 97174 107528 97180
rect 70032 97096 70084 97102
rect 70032 97038 70084 97044
rect 71872 97096 71924 97102
rect 71872 97038 71924 97044
rect 72516 97096 72568 97102
rect 72516 97038 72568 97044
rect 74172 97096 74224 97102
rect 74172 97038 74224 97044
rect 69296 96620 69348 96626
rect 69296 96562 69348 96568
rect 68836 96484 68888 96490
rect 68836 96426 68888 96432
rect 68008 96212 68060 96218
rect 68008 96154 68060 96160
rect 69112 95940 69164 95946
rect 69112 95882 69164 95888
rect 67732 95464 67784 95470
rect 67732 95406 67784 95412
rect 69020 95464 69072 95470
rect 69020 95406 69072 95412
rect 67744 93226 67772 95406
rect 68836 94920 68888 94926
rect 68836 94862 68888 94868
rect 68848 94042 68876 94862
rect 68836 94036 68888 94042
rect 68836 93978 68888 93984
rect 68284 93764 68336 93770
rect 68284 93706 68336 93712
rect 67824 93356 67876 93362
rect 67824 93298 67876 93304
rect 67732 93220 67784 93226
rect 67732 93162 67784 93168
rect 67640 92404 67692 92410
rect 67640 92346 67692 92352
rect 67836 92138 67864 93298
rect 68296 92138 68324 93706
rect 68376 93424 68428 93430
rect 68376 93366 68428 93372
rect 68388 93294 68416 93366
rect 68376 93288 68428 93294
rect 68376 93230 68428 93236
rect 69032 93158 69060 95406
rect 69124 93838 69152 95882
rect 69308 95130 69336 96562
rect 69940 95600 69992 95606
rect 69940 95542 69992 95548
rect 69296 95124 69348 95130
rect 69296 95066 69348 95072
rect 69756 94852 69808 94858
rect 69756 94794 69808 94800
rect 69112 93832 69164 93838
rect 69112 93774 69164 93780
rect 69204 93356 69256 93362
rect 69204 93298 69256 93304
rect 69216 93265 69244 93298
rect 69202 93256 69258 93265
rect 69202 93191 69258 93200
rect 69768 93158 69796 94794
rect 69952 93498 69980 95542
rect 70044 95402 70072 97038
rect 70768 96008 70820 96014
rect 70768 95950 70820 95956
rect 70584 95600 70636 95606
rect 70780 95554 70808 95950
rect 71884 95674 71912 97038
rect 71964 95940 72016 95946
rect 71964 95882 72016 95888
rect 71872 95668 71924 95674
rect 71872 95610 71924 95616
rect 70636 95548 70808 95554
rect 70584 95542 70808 95548
rect 71688 95600 71740 95606
rect 71688 95542 71740 95548
rect 70596 95526 70808 95542
rect 70032 95396 70084 95402
rect 70032 95338 70084 95344
rect 70780 94926 70808 95526
rect 70768 94920 70820 94926
rect 70768 94862 70820 94868
rect 70492 94308 70544 94314
rect 70492 94250 70544 94256
rect 70504 93770 70532 94250
rect 70124 93764 70176 93770
rect 70124 93706 70176 93712
rect 70492 93764 70544 93770
rect 70492 93706 70544 93712
rect 69848 93492 69900 93498
rect 69848 93434 69900 93440
rect 69940 93492 69992 93498
rect 69940 93434 69992 93440
rect 69860 93158 69888 93434
rect 70136 93430 70164 93706
rect 70124 93424 70176 93430
rect 70124 93366 70176 93372
rect 70136 93294 70164 93366
rect 70308 93356 70360 93362
rect 70308 93298 70360 93304
rect 69940 93288 69992 93294
rect 69940 93230 69992 93236
rect 70124 93288 70176 93294
rect 70124 93230 70176 93236
rect 68560 93152 68612 93158
rect 68560 93094 68612 93100
rect 69020 93152 69072 93158
rect 69020 93094 69072 93100
rect 69756 93152 69808 93158
rect 69756 93094 69808 93100
rect 69848 93152 69900 93158
rect 69848 93094 69900 93100
rect 68572 92886 68600 93094
rect 69952 92886 69980 93230
rect 70320 92954 70348 93298
rect 70584 93152 70636 93158
rect 70584 93094 70636 93100
rect 70596 92954 70624 93094
rect 70308 92948 70360 92954
rect 70308 92890 70360 92896
rect 70584 92948 70636 92954
rect 70584 92890 70636 92896
rect 68560 92880 68612 92886
rect 68560 92822 68612 92828
rect 69940 92880 69992 92886
rect 69940 92822 69992 92828
rect 69204 92676 69256 92682
rect 69204 92618 69256 92624
rect 69572 92676 69624 92682
rect 69572 92618 69624 92624
rect 70492 92676 70544 92682
rect 70492 92618 70544 92624
rect 69216 92585 69244 92618
rect 69202 92576 69258 92585
rect 69202 92511 69258 92520
rect 69584 92274 69612 92618
rect 70504 92585 70532 92618
rect 70490 92576 70546 92585
rect 70490 92511 70546 92520
rect 69572 92268 69624 92274
rect 69572 92210 69624 92216
rect 70780 92138 70808 94862
rect 70860 93696 70912 93702
rect 70860 93638 70912 93644
rect 71136 93696 71188 93702
rect 71136 93638 71188 93644
rect 70872 93498 70900 93638
rect 70860 93492 70912 93498
rect 70860 93434 70912 93440
rect 67824 92132 67876 92138
rect 67824 92074 67876 92080
rect 68284 92132 68336 92138
rect 68284 92074 68336 92080
rect 70768 92132 70820 92138
rect 70768 92074 70820 92080
rect 71148 90438 71176 93638
rect 71700 93498 71728 95542
rect 71688 93492 71740 93498
rect 71688 93434 71740 93440
rect 71976 93158 72004 95882
rect 72528 95130 72556 97038
rect 74184 96218 74212 97038
rect 107844 96960 107896 96966
rect 107844 96902 107896 96908
rect 97034 96860 97342 96869
rect 97034 96858 97040 96860
rect 97096 96858 97120 96860
rect 97176 96858 97200 96860
rect 97256 96858 97280 96860
rect 97336 96858 97342 96860
rect 97096 96806 97098 96858
rect 97278 96806 97280 96858
rect 97034 96804 97040 96806
rect 97096 96804 97120 96806
rect 97176 96804 97200 96806
rect 97256 96804 97280 96806
rect 97336 96804 97342 96806
rect 97034 96795 97342 96804
rect 96374 96316 96682 96325
rect 96374 96314 96380 96316
rect 96436 96314 96460 96316
rect 96516 96314 96540 96316
rect 96596 96314 96620 96316
rect 96676 96314 96682 96316
rect 96436 96262 96438 96314
rect 96618 96262 96620 96314
rect 96374 96260 96380 96262
rect 96436 96260 96460 96262
rect 96516 96260 96540 96262
rect 96596 96260 96620 96262
rect 96676 96260 96682 96262
rect 96374 96251 96682 96260
rect 74172 96212 74224 96218
rect 74172 96154 74224 96160
rect 74724 95940 74776 95946
rect 74724 95882 74776 95888
rect 72516 95124 72568 95130
rect 72516 95066 72568 95072
rect 72976 94852 73028 94858
rect 72976 94794 73028 94800
rect 72240 93832 72292 93838
rect 72240 93774 72292 93780
rect 72148 93696 72200 93702
rect 72148 93638 72200 93644
rect 72056 93424 72108 93430
rect 72056 93366 72108 93372
rect 71964 93152 72016 93158
rect 71964 93094 72016 93100
rect 71872 92200 71924 92206
rect 71872 92142 71924 92148
rect 71136 90432 71188 90438
rect 71136 90374 71188 90380
rect 71884 89729 71912 92142
rect 72068 92138 72096 93366
rect 72160 93294 72188 93638
rect 72252 93430 72280 93774
rect 72988 93498 73016 94794
rect 74736 93498 74764 95882
rect 97034 95772 97342 95781
rect 97034 95770 97040 95772
rect 97096 95770 97120 95772
rect 97176 95770 97200 95772
rect 97256 95770 97280 95772
rect 97336 95770 97342 95772
rect 97096 95718 97098 95770
rect 97278 95718 97280 95770
rect 97034 95716 97040 95718
rect 97096 95716 97120 95718
rect 97176 95716 97200 95718
rect 97256 95716 97280 95718
rect 97336 95716 97342 95718
rect 97034 95707 97342 95716
rect 96374 95228 96682 95237
rect 96374 95226 96380 95228
rect 96436 95226 96460 95228
rect 96516 95226 96540 95228
rect 96596 95226 96620 95228
rect 96676 95226 96682 95228
rect 96436 95174 96438 95226
rect 96618 95174 96620 95226
rect 96374 95172 96380 95174
rect 96436 95172 96460 95174
rect 96516 95172 96540 95174
rect 96596 95172 96620 95174
rect 96676 95172 96682 95174
rect 96374 95163 96682 95172
rect 97034 94684 97342 94693
rect 97034 94682 97040 94684
rect 97096 94682 97120 94684
rect 97176 94682 97200 94684
rect 97256 94682 97280 94684
rect 97336 94682 97342 94684
rect 97096 94630 97098 94682
rect 97278 94630 97280 94682
rect 97034 94628 97040 94630
rect 97096 94628 97120 94630
rect 97176 94628 97200 94630
rect 97256 94628 97280 94630
rect 97336 94628 97342 94630
rect 97034 94619 97342 94628
rect 96374 94140 96682 94149
rect 96374 94138 96380 94140
rect 96436 94138 96460 94140
rect 96516 94138 96540 94140
rect 96596 94138 96620 94140
rect 96676 94138 96682 94140
rect 96436 94086 96438 94138
rect 96618 94086 96620 94138
rect 96374 94084 96380 94086
rect 96436 94084 96460 94086
rect 96516 94084 96540 94086
rect 96596 94084 96620 94086
rect 96676 94084 96682 94086
rect 96374 94075 96682 94084
rect 97034 93596 97342 93605
rect 97034 93594 97040 93596
rect 97096 93594 97120 93596
rect 97176 93594 97200 93596
rect 97256 93594 97280 93596
rect 97336 93594 97342 93596
rect 97096 93542 97098 93594
rect 97278 93542 97280 93594
rect 97034 93540 97040 93542
rect 97096 93540 97120 93542
rect 97176 93540 97200 93542
rect 97256 93540 97280 93542
rect 97336 93540 97342 93542
rect 97034 93531 97342 93540
rect 72976 93492 73028 93498
rect 72976 93434 73028 93440
rect 74724 93492 74776 93498
rect 74724 93434 74776 93440
rect 72240 93424 72292 93430
rect 72240 93366 72292 93372
rect 72148 93288 72200 93294
rect 72148 93230 72200 93236
rect 74172 93288 74224 93294
rect 74172 93230 74224 93236
rect 72160 92750 72188 93230
rect 72148 92744 72200 92750
rect 72148 92686 72200 92692
rect 72976 92744 73028 92750
rect 72976 92686 73028 92692
rect 72988 92410 73016 92686
rect 73252 92676 73304 92682
rect 73252 92618 73304 92624
rect 73712 92676 73764 92682
rect 73712 92618 73764 92624
rect 72976 92404 73028 92410
rect 72976 92346 73028 92352
rect 72056 92132 72108 92138
rect 72056 92074 72108 92080
rect 73264 91089 73292 92618
rect 73250 91080 73306 91089
rect 73250 91015 73306 91024
rect 73724 89729 73752 92618
rect 74184 91089 74212 93230
rect 107856 93226 107884 96902
rect 107844 93220 107896 93226
rect 107844 93162 107896 93168
rect 108580 93152 108632 93158
rect 108580 93094 108632 93100
rect 96374 93052 96682 93061
rect 96374 93050 96380 93052
rect 96436 93050 96460 93052
rect 96516 93050 96540 93052
rect 96596 93050 96620 93052
rect 96676 93050 96682 93052
rect 96436 92998 96438 93050
rect 96618 92998 96620 93050
rect 96374 92996 96380 92998
rect 96436 92996 96460 92998
rect 96516 92996 96540 92998
rect 96596 92996 96620 92998
rect 96676 92996 96682 92998
rect 96374 92987 96682 92996
rect 77484 92676 77536 92682
rect 77484 92618 77536 92624
rect 74724 92608 74776 92614
rect 74724 92550 74776 92556
rect 74736 92274 74764 92550
rect 77496 92410 77524 92618
rect 79416 92608 79468 92614
rect 79416 92550 79468 92556
rect 77484 92404 77536 92410
rect 77484 92346 77536 92352
rect 74724 92268 74776 92274
rect 74724 92210 74776 92216
rect 75920 92200 75972 92206
rect 75920 92142 75972 92148
rect 74170 91080 74226 91089
rect 74170 91015 74226 91024
rect 75932 89729 75960 92142
rect 77496 91798 77524 92346
rect 79428 92070 79456 92550
rect 97034 92508 97342 92517
rect 97034 92506 97040 92508
rect 97096 92506 97120 92508
rect 97176 92506 97200 92508
rect 97256 92506 97280 92508
rect 97336 92506 97342 92508
rect 97096 92454 97098 92506
rect 97278 92454 97280 92506
rect 97034 92452 97040 92454
rect 97096 92452 97120 92454
rect 97176 92452 97200 92454
rect 97256 92452 97280 92454
rect 97336 92452 97342 92454
rect 97034 92443 97342 92452
rect 100024 92132 100076 92138
rect 100024 92074 100076 92080
rect 79416 92064 79468 92070
rect 79416 92006 79468 92012
rect 89444 92064 89496 92070
rect 89444 92006 89496 92012
rect 77484 91792 77536 91798
rect 77484 91734 77536 91740
rect 89456 89729 89484 92006
rect 96374 91964 96682 91973
rect 96374 91962 96380 91964
rect 96436 91962 96460 91964
rect 96516 91962 96540 91964
rect 96596 91962 96620 91964
rect 96676 91962 96682 91964
rect 96436 91910 96438 91962
rect 96618 91910 96620 91962
rect 96374 91908 96380 91910
rect 96436 91908 96460 91910
rect 96516 91908 96540 91910
rect 96596 91908 96620 91910
rect 96676 91908 96682 91910
rect 96374 91899 96682 91908
rect 100036 91225 100064 92074
rect 108304 91792 108356 91798
rect 108304 91734 108356 91740
rect 100022 91216 100078 91225
rect 100022 91151 100078 91160
rect 65246 89720 65302 89729
rect 65246 89655 65302 89664
rect 66810 89720 66866 89729
rect 66810 89655 66866 89664
rect 67546 89720 67602 89729
rect 67546 89655 67602 89664
rect 71870 89720 71926 89729
rect 71870 89655 71926 89664
rect 73710 89720 73766 89729
rect 73710 89655 73766 89664
rect 75918 89720 75974 89729
rect 75918 89655 75974 89664
rect 89442 89720 89498 89729
rect 89442 89655 89498 89664
rect 60554 89584 60610 89593
rect 60554 89519 60610 89528
rect 106922 89584 106978 89593
rect 106922 89519 106978 89528
rect 106188 86624 106240 86630
rect 106188 86566 106240 86572
rect 106200 86507 106228 86566
rect 106186 86498 106242 86507
rect 106186 86433 106242 86442
rect 106936 52086 106964 89519
rect 108316 54330 108344 91734
rect 108396 90432 108448 90438
rect 108396 90374 108448 90380
rect 108408 67386 108436 90374
rect 108396 67380 108448 67386
rect 108396 67322 108448 67328
rect 108592 54874 108620 93094
rect 113650 92508 113958 92517
rect 113650 92506 113656 92508
rect 113712 92506 113736 92508
rect 113792 92506 113816 92508
rect 113872 92506 113896 92508
rect 113952 92506 113958 92508
rect 113712 92454 113714 92506
rect 113894 92454 113896 92506
rect 113650 92452 113656 92454
rect 113712 92452 113736 92454
rect 113792 92452 113816 92454
rect 113872 92452 113896 92454
rect 113952 92452 113958 92454
rect 113650 92443 113958 92452
rect 112914 91964 113222 91973
rect 112914 91962 112920 91964
rect 112976 91962 113000 91964
rect 113056 91962 113080 91964
rect 113136 91962 113160 91964
rect 113216 91962 113222 91964
rect 112976 91910 112978 91962
rect 113158 91910 113160 91962
rect 112914 91908 112920 91910
rect 112976 91908 113000 91910
rect 113056 91908 113080 91910
rect 113136 91908 113160 91910
rect 113216 91908 113222 91910
rect 112914 91899 113222 91908
rect 113650 91420 113958 91429
rect 113650 91418 113656 91420
rect 113712 91418 113736 91420
rect 113792 91418 113816 91420
rect 113872 91418 113896 91420
rect 113952 91418 113958 91420
rect 113712 91366 113714 91418
rect 113894 91366 113896 91418
rect 113650 91364 113656 91366
rect 113712 91364 113736 91366
rect 113792 91364 113816 91366
rect 113872 91364 113896 91366
rect 113952 91364 113958 91366
rect 113650 91355 113958 91364
rect 112914 90876 113222 90885
rect 112914 90874 112920 90876
rect 112976 90874 113000 90876
rect 113056 90874 113080 90876
rect 113136 90874 113160 90876
rect 113216 90874 113222 90876
rect 112976 90822 112978 90874
rect 113158 90822 113160 90874
rect 112914 90820 112920 90822
rect 112976 90820 113000 90822
rect 113056 90820 113080 90822
rect 113136 90820 113160 90822
rect 113216 90820 113222 90822
rect 112914 90811 113222 90820
rect 113650 90332 113958 90341
rect 113650 90330 113656 90332
rect 113712 90330 113736 90332
rect 113792 90330 113816 90332
rect 113872 90330 113896 90332
rect 113952 90330 113958 90332
rect 113712 90278 113714 90330
rect 113894 90278 113896 90330
rect 113650 90276 113656 90278
rect 113712 90276 113736 90278
rect 113792 90276 113816 90278
rect 113872 90276 113896 90278
rect 113952 90276 113958 90278
rect 113650 90267 113958 90276
rect 112914 89788 113222 89797
rect 112914 89786 112920 89788
rect 112976 89786 113000 89788
rect 113056 89786 113080 89788
rect 113136 89786 113160 89788
rect 113216 89786 113222 89788
rect 112976 89734 112978 89786
rect 113158 89734 113160 89786
rect 112914 89732 112920 89734
rect 112976 89732 113000 89734
rect 113056 89732 113080 89734
rect 113136 89732 113160 89734
rect 113216 89732 113222 89734
rect 112914 89723 113222 89732
rect 113650 89244 113958 89253
rect 113650 89242 113656 89244
rect 113712 89242 113736 89244
rect 113792 89242 113816 89244
rect 113872 89242 113896 89244
rect 113952 89242 113958 89244
rect 113712 89190 113714 89242
rect 113894 89190 113896 89242
rect 113650 89188 113656 89190
rect 113712 89188 113736 89190
rect 113792 89188 113816 89190
rect 113872 89188 113896 89190
rect 113952 89188 113958 89190
rect 113650 89179 113958 89188
rect 112914 88700 113222 88709
rect 112914 88698 112920 88700
rect 112976 88698 113000 88700
rect 113056 88698 113080 88700
rect 113136 88698 113160 88700
rect 113216 88698 113222 88700
rect 112976 88646 112978 88698
rect 113158 88646 113160 88698
rect 112914 88644 112920 88646
rect 112976 88644 113000 88646
rect 113056 88644 113080 88646
rect 113136 88644 113160 88646
rect 113216 88644 113222 88646
rect 112914 88635 113222 88644
rect 113650 88156 113958 88165
rect 113650 88154 113656 88156
rect 113712 88154 113736 88156
rect 113792 88154 113816 88156
rect 113872 88154 113896 88156
rect 113952 88154 113958 88156
rect 113712 88102 113714 88154
rect 113894 88102 113896 88154
rect 113650 88100 113656 88102
rect 113712 88100 113736 88102
rect 113792 88100 113816 88102
rect 113872 88100 113896 88102
rect 113952 88100 113958 88102
rect 113650 88091 113958 88100
rect 112914 87612 113222 87621
rect 112914 87610 112920 87612
rect 112976 87610 113000 87612
rect 113056 87610 113080 87612
rect 113136 87610 113160 87612
rect 113216 87610 113222 87612
rect 112976 87558 112978 87610
rect 113158 87558 113160 87610
rect 112914 87556 112920 87558
rect 112976 87556 113000 87558
rect 113056 87556 113080 87558
rect 113136 87556 113160 87558
rect 113216 87556 113222 87558
rect 112914 87547 113222 87556
rect 113650 87068 113958 87077
rect 113650 87066 113656 87068
rect 113712 87066 113736 87068
rect 113792 87066 113816 87068
rect 113872 87066 113896 87068
rect 113952 87066 113958 87068
rect 113712 87014 113714 87066
rect 113894 87014 113896 87066
rect 113650 87012 113656 87014
rect 113712 87012 113736 87014
rect 113792 87012 113816 87014
rect 113872 87012 113896 87014
rect 113952 87012 113958 87014
rect 113650 87003 113958 87012
rect 112914 86524 113222 86533
rect 112914 86522 112920 86524
rect 112976 86522 113000 86524
rect 113056 86522 113080 86524
rect 113136 86522 113160 86524
rect 113216 86522 113222 86524
rect 112976 86470 112978 86522
rect 113158 86470 113160 86522
rect 112914 86468 112920 86470
rect 112976 86468 113000 86470
rect 113056 86468 113080 86470
rect 113136 86468 113160 86470
rect 113216 86468 113222 86470
rect 112914 86459 113222 86468
rect 113650 85980 113958 85989
rect 113650 85978 113656 85980
rect 113712 85978 113736 85980
rect 113792 85978 113816 85980
rect 113872 85978 113896 85980
rect 113952 85978 113958 85980
rect 113712 85926 113714 85978
rect 113894 85926 113896 85978
rect 113650 85924 113656 85926
rect 113712 85924 113736 85926
rect 113792 85924 113816 85926
rect 113872 85924 113896 85926
rect 113952 85924 113958 85926
rect 113650 85915 113958 85924
rect 112914 85436 113222 85445
rect 112914 85434 112920 85436
rect 112976 85434 113000 85436
rect 113056 85434 113080 85436
rect 113136 85434 113160 85436
rect 113216 85434 113222 85436
rect 112976 85382 112978 85434
rect 113158 85382 113160 85434
rect 112914 85380 112920 85382
rect 112976 85380 113000 85382
rect 113056 85380 113080 85382
rect 113136 85380 113160 85382
rect 113216 85380 113222 85382
rect 112914 85371 113222 85380
rect 113650 84892 113958 84901
rect 113650 84890 113656 84892
rect 113712 84890 113736 84892
rect 113792 84890 113816 84892
rect 113872 84890 113896 84892
rect 113952 84890 113958 84892
rect 113712 84838 113714 84890
rect 113894 84838 113896 84890
rect 113650 84836 113656 84838
rect 113712 84836 113736 84838
rect 113792 84836 113816 84838
rect 113872 84836 113896 84838
rect 113952 84836 113958 84838
rect 113650 84827 113958 84836
rect 112914 84348 113222 84357
rect 112914 84346 112920 84348
rect 112976 84346 113000 84348
rect 113056 84346 113080 84348
rect 113136 84346 113160 84348
rect 113216 84346 113222 84348
rect 112976 84294 112978 84346
rect 113158 84294 113160 84346
rect 112914 84292 112920 84294
rect 112976 84292 113000 84294
rect 113056 84292 113080 84294
rect 113136 84292 113160 84294
rect 113216 84292 113222 84294
rect 112914 84283 113222 84292
rect 113650 83804 113958 83813
rect 113650 83802 113656 83804
rect 113712 83802 113736 83804
rect 113792 83802 113816 83804
rect 113872 83802 113896 83804
rect 113952 83802 113958 83804
rect 113712 83750 113714 83802
rect 113894 83750 113896 83802
rect 113650 83748 113656 83750
rect 113712 83748 113736 83750
rect 113792 83748 113816 83750
rect 113872 83748 113896 83750
rect 113952 83748 113958 83750
rect 113650 83739 113958 83748
rect 112914 83260 113222 83269
rect 112914 83258 112920 83260
rect 112976 83258 113000 83260
rect 113056 83258 113080 83260
rect 113136 83258 113160 83260
rect 113216 83258 113222 83260
rect 112976 83206 112978 83258
rect 113158 83206 113160 83258
rect 112914 83204 112920 83206
rect 112976 83204 113000 83206
rect 113056 83204 113080 83206
rect 113136 83204 113160 83206
rect 113216 83204 113222 83206
rect 112914 83195 113222 83204
rect 113650 82716 113958 82725
rect 113650 82714 113656 82716
rect 113712 82714 113736 82716
rect 113792 82714 113816 82716
rect 113872 82714 113896 82716
rect 113952 82714 113958 82716
rect 113712 82662 113714 82714
rect 113894 82662 113896 82714
rect 113650 82660 113656 82662
rect 113712 82660 113736 82662
rect 113792 82660 113816 82662
rect 113872 82660 113896 82662
rect 113952 82660 113958 82662
rect 113650 82651 113958 82660
rect 112914 82172 113222 82181
rect 112914 82170 112920 82172
rect 112976 82170 113000 82172
rect 113056 82170 113080 82172
rect 113136 82170 113160 82172
rect 113216 82170 113222 82172
rect 112976 82118 112978 82170
rect 113158 82118 113160 82170
rect 112914 82116 112920 82118
rect 112976 82116 113000 82118
rect 113056 82116 113080 82118
rect 113136 82116 113160 82118
rect 113216 82116 113222 82118
rect 112914 82107 113222 82116
rect 113650 81628 113958 81637
rect 113650 81626 113656 81628
rect 113712 81626 113736 81628
rect 113792 81626 113816 81628
rect 113872 81626 113896 81628
rect 113952 81626 113958 81628
rect 113712 81574 113714 81626
rect 113894 81574 113896 81626
rect 113650 81572 113656 81574
rect 113712 81572 113736 81574
rect 113792 81572 113816 81574
rect 113872 81572 113896 81574
rect 113952 81572 113958 81574
rect 113650 81563 113958 81572
rect 112914 81084 113222 81093
rect 112914 81082 112920 81084
rect 112976 81082 113000 81084
rect 113056 81082 113080 81084
rect 113136 81082 113160 81084
rect 113216 81082 113222 81084
rect 112976 81030 112978 81082
rect 113158 81030 113160 81082
rect 112914 81028 112920 81030
rect 112976 81028 113000 81030
rect 113056 81028 113080 81030
rect 113136 81028 113160 81030
rect 113216 81028 113222 81030
rect 112914 81019 113222 81028
rect 113650 80540 113958 80549
rect 113650 80538 113656 80540
rect 113712 80538 113736 80540
rect 113792 80538 113816 80540
rect 113872 80538 113896 80540
rect 113952 80538 113958 80540
rect 113712 80486 113714 80538
rect 113894 80486 113896 80538
rect 113650 80484 113656 80486
rect 113712 80484 113736 80486
rect 113792 80484 113816 80486
rect 113872 80484 113896 80486
rect 113952 80484 113958 80486
rect 113650 80475 113958 80484
rect 112914 79996 113222 80005
rect 112914 79994 112920 79996
rect 112976 79994 113000 79996
rect 113056 79994 113080 79996
rect 113136 79994 113160 79996
rect 113216 79994 113222 79996
rect 112976 79942 112978 79994
rect 113158 79942 113160 79994
rect 112914 79940 112920 79942
rect 112976 79940 113000 79942
rect 113056 79940 113080 79942
rect 113136 79940 113160 79942
rect 113216 79940 113222 79942
rect 112914 79931 113222 79940
rect 113650 79452 113958 79461
rect 113650 79450 113656 79452
rect 113712 79450 113736 79452
rect 113792 79450 113816 79452
rect 113872 79450 113896 79452
rect 113952 79450 113958 79452
rect 113712 79398 113714 79450
rect 113894 79398 113896 79450
rect 113650 79396 113656 79398
rect 113712 79396 113736 79398
rect 113792 79396 113816 79398
rect 113872 79396 113896 79398
rect 113952 79396 113958 79398
rect 113650 79387 113958 79396
rect 112914 78908 113222 78917
rect 112914 78906 112920 78908
rect 112976 78906 113000 78908
rect 113056 78906 113080 78908
rect 113136 78906 113160 78908
rect 113216 78906 113222 78908
rect 112976 78854 112978 78906
rect 113158 78854 113160 78906
rect 112914 78852 112920 78854
rect 112976 78852 113000 78854
rect 113056 78852 113080 78854
rect 113136 78852 113160 78854
rect 113216 78852 113222 78854
rect 112914 78843 113222 78852
rect 113650 78364 113958 78373
rect 113650 78362 113656 78364
rect 113712 78362 113736 78364
rect 113792 78362 113816 78364
rect 113872 78362 113896 78364
rect 113952 78362 113958 78364
rect 113712 78310 113714 78362
rect 113894 78310 113896 78362
rect 113650 78308 113656 78310
rect 113712 78308 113736 78310
rect 113792 78308 113816 78310
rect 113872 78308 113896 78310
rect 113952 78308 113958 78310
rect 113650 78299 113958 78308
rect 112914 77820 113222 77829
rect 112914 77818 112920 77820
rect 112976 77818 113000 77820
rect 113056 77818 113080 77820
rect 113136 77818 113160 77820
rect 113216 77818 113222 77820
rect 112976 77766 112978 77818
rect 113158 77766 113160 77818
rect 112914 77764 112920 77766
rect 112976 77764 113000 77766
rect 113056 77764 113080 77766
rect 113136 77764 113160 77766
rect 113216 77764 113222 77766
rect 112914 77755 113222 77764
rect 113650 77276 113958 77285
rect 113650 77274 113656 77276
rect 113712 77274 113736 77276
rect 113792 77274 113816 77276
rect 113872 77274 113896 77276
rect 113952 77274 113958 77276
rect 113712 77222 113714 77274
rect 113894 77222 113896 77274
rect 113650 77220 113656 77222
rect 113712 77220 113736 77222
rect 113792 77220 113816 77222
rect 113872 77220 113896 77222
rect 113952 77220 113958 77222
rect 113650 77211 113958 77220
rect 112914 76732 113222 76741
rect 112914 76730 112920 76732
rect 112976 76730 113000 76732
rect 113056 76730 113080 76732
rect 113136 76730 113160 76732
rect 113216 76730 113222 76732
rect 112976 76678 112978 76730
rect 113158 76678 113160 76730
rect 112914 76676 112920 76678
rect 112976 76676 113000 76678
rect 113056 76676 113080 76678
rect 113136 76676 113160 76678
rect 113216 76676 113222 76678
rect 112914 76667 113222 76676
rect 113650 76188 113958 76197
rect 113650 76186 113656 76188
rect 113712 76186 113736 76188
rect 113792 76186 113816 76188
rect 113872 76186 113896 76188
rect 113952 76186 113958 76188
rect 113712 76134 113714 76186
rect 113894 76134 113896 76186
rect 113650 76132 113656 76134
rect 113712 76132 113736 76134
rect 113792 76132 113816 76134
rect 113872 76132 113896 76134
rect 113952 76132 113958 76134
rect 113650 76123 113958 76132
rect 112914 75644 113222 75653
rect 112914 75642 112920 75644
rect 112976 75642 113000 75644
rect 113056 75642 113080 75644
rect 113136 75642 113160 75644
rect 113216 75642 113222 75644
rect 112976 75590 112978 75642
rect 113158 75590 113160 75642
rect 112914 75588 112920 75590
rect 112976 75588 113000 75590
rect 113056 75588 113080 75590
rect 113136 75588 113160 75590
rect 113216 75588 113222 75590
rect 112914 75579 113222 75588
rect 113650 75100 113958 75109
rect 113650 75098 113656 75100
rect 113712 75098 113736 75100
rect 113792 75098 113816 75100
rect 113872 75098 113896 75100
rect 113952 75098 113958 75100
rect 113712 75046 113714 75098
rect 113894 75046 113896 75098
rect 113650 75044 113656 75046
rect 113712 75044 113736 75046
rect 113792 75044 113816 75046
rect 113872 75044 113896 75046
rect 113952 75044 113958 75046
rect 113650 75035 113958 75044
rect 112914 74556 113222 74565
rect 112914 74554 112920 74556
rect 112976 74554 113000 74556
rect 113056 74554 113080 74556
rect 113136 74554 113160 74556
rect 113216 74554 113222 74556
rect 112976 74502 112978 74554
rect 113158 74502 113160 74554
rect 112914 74500 112920 74502
rect 112976 74500 113000 74502
rect 113056 74500 113080 74502
rect 113136 74500 113160 74502
rect 113216 74500 113222 74502
rect 112914 74491 113222 74500
rect 113650 74012 113958 74021
rect 113650 74010 113656 74012
rect 113712 74010 113736 74012
rect 113792 74010 113816 74012
rect 113872 74010 113896 74012
rect 113952 74010 113958 74012
rect 113712 73958 113714 74010
rect 113894 73958 113896 74010
rect 113650 73956 113656 73958
rect 113712 73956 113736 73958
rect 113792 73956 113816 73958
rect 113872 73956 113896 73958
rect 113952 73956 113958 73958
rect 113650 73947 113958 73956
rect 112914 73468 113222 73477
rect 112914 73466 112920 73468
rect 112976 73466 113000 73468
rect 113056 73466 113080 73468
rect 113136 73466 113160 73468
rect 113216 73466 113222 73468
rect 112976 73414 112978 73466
rect 113158 73414 113160 73466
rect 112914 73412 112920 73414
rect 112976 73412 113000 73414
rect 113056 73412 113080 73414
rect 113136 73412 113160 73414
rect 113216 73412 113222 73414
rect 112914 73403 113222 73412
rect 113650 72924 113958 72933
rect 113650 72922 113656 72924
rect 113712 72922 113736 72924
rect 113792 72922 113816 72924
rect 113872 72922 113896 72924
rect 113952 72922 113958 72924
rect 113712 72870 113714 72922
rect 113894 72870 113896 72922
rect 113650 72868 113656 72870
rect 113712 72868 113736 72870
rect 113792 72868 113816 72870
rect 113872 72868 113896 72870
rect 113952 72868 113958 72870
rect 113650 72859 113958 72868
rect 112914 72380 113222 72389
rect 112914 72378 112920 72380
rect 112976 72378 113000 72380
rect 113056 72378 113080 72380
rect 113136 72378 113160 72380
rect 113216 72378 113222 72380
rect 112976 72326 112978 72378
rect 113158 72326 113160 72378
rect 112914 72324 112920 72326
rect 112976 72324 113000 72326
rect 113056 72324 113080 72326
rect 113136 72324 113160 72326
rect 113216 72324 113222 72326
rect 112914 72315 113222 72324
rect 113650 71836 113958 71845
rect 113650 71834 113656 71836
rect 113712 71834 113736 71836
rect 113792 71834 113816 71836
rect 113872 71834 113896 71836
rect 113952 71834 113958 71836
rect 113712 71782 113714 71834
rect 113894 71782 113896 71834
rect 113650 71780 113656 71782
rect 113712 71780 113736 71782
rect 113792 71780 113816 71782
rect 113872 71780 113896 71782
rect 113952 71780 113958 71782
rect 113650 71771 113958 71780
rect 112914 71292 113222 71301
rect 112914 71290 112920 71292
rect 112976 71290 113000 71292
rect 113056 71290 113080 71292
rect 113136 71290 113160 71292
rect 113216 71290 113222 71292
rect 112976 71238 112978 71290
rect 113158 71238 113160 71290
rect 112914 71236 112920 71238
rect 112976 71236 113000 71238
rect 113056 71236 113080 71238
rect 113136 71236 113160 71238
rect 113216 71236 113222 71238
rect 112914 71227 113222 71236
rect 113650 70748 113958 70757
rect 113650 70746 113656 70748
rect 113712 70746 113736 70748
rect 113792 70746 113816 70748
rect 113872 70746 113896 70748
rect 113952 70746 113958 70748
rect 113712 70694 113714 70746
rect 113894 70694 113896 70746
rect 113650 70692 113656 70694
rect 113712 70692 113736 70694
rect 113792 70692 113816 70694
rect 113872 70692 113896 70694
rect 113952 70692 113958 70694
rect 113650 70683 113958 70692
rect 112914 70204 113222 70213
rect 112914 70202 112920 70204
rect 112976 70202 113000 70204
rect 113056 70202 113080 70204
rect 113136 70202 113160 70204
rect 113216 70202 113222 70204
rect 112976 70150 112978 70202
rect 113158 70150 113160 70202
rect 112914 70148 112920 70150
rect 112976 70148 113000 70150
rect 113056 70148 113080 70150
rect 113136 70148 113160 70150
rect 113216 70148 113222 70150
rect 112914 70139 113222 70148
rect 113650 69660 113958 69669
rect 113650 69658 113656 69660
rect 113712 69658 113736 69660
rect 113792 69658 113816 69660
rect 113872 69658 113896 69660
rect 113952 69658 113958 69660
rect 113712 69606 113714 69658
rect 113894 69606 113896 69658
rect 113650 69604 113656 69606
rect 113712 69604 113736 69606
rect 113792 69604 113816 69606
rect 113872 69604 113896 69606
rect 113952 69604 113958 69606
rect 113650 69595 113958 69604
rect 112914 69116 113222 69125
rect 112914 69114 112920 69116
rect 112976 69114 113000 69116
rect 113056 69114 113080 69116
rect 113136 69114 113160 69116
rect 113216 69114 113222 69116
rect 112976 69062 112978 69114
rect 113158 69062 113160 69114
rect 112914 69060 112920 69062
rect 112976 69060 113000 69062
rect 113056 69060 113080 69062
rect 113136 69060 113160 69062
rect 113216 69060 113222 69062
rect 112914 69051 113222 69060
rect 113650 68572 113958 68581
rect 113650 68570 113656 68572
rect 113712 68570 113736 68572
rect 113792 68570 113816 68572
rect 113872 68570 113896 68572
rect 113952 68570 113958 68572
rect 113712 68518 113714 68570
rect 113894 68518 113896 68570
rect 113650 68516 113656 68518
rect 113712 68516 113736 68518
rect 113792 68516 113816 68518
rect 113872 68516 113896 68518
rect 113952 68516 113958 68518
rect 113650 68507 113958 68516
rect 112914 68028 113222 68037
rect 112914 68026 112920 68028
rect 112976 68026 113000 68028
rect 113056 68026 113080 68028
rect 113136 68026 113160 68028
rect 113216 68026 113222 68028
rect 112976 67974 112978 68026
rect 113158 67974 113160 68026
rect 112914 67972 112920 67974
rect 112976 67972 113000 67974
rect 113056 67972 113080 67974
rect 113136 67972 113160 67974
rect 113216 67972 113222 67974
rect 112914 67963 113222 67972
rect 113650 67484 113958 67493
rect 113650 67482 113656 67484
rect 113712 67482 113736 67484
rect 113792 67482 113816 67484
rect 113872 67482 113896 67484
rect 113952 67482 113958 67484
rect 113712 67430 113714 67482
rect 113894 67430 113896 67482
rect 113650 67428 113656 67430
rect 113712 67428 113736 67430
rect 113792 67428 113816 67430
rect 113872 67428 113896 67430
rect 113952 67428 113958 67430
rect 113650 67419 113958 67428
rect 109684 67244 109736 67250
rect 109684 67186 109736 67192
rect 108672 57860 108724 57866
rect 108672 57802 108724 57808
rect 108684 55214 108712 57802
rect 109696 57798 109724 67186
rect 109960 67040 110012 67046
rect 109960 66982 110012 66988
rect 109972 57934 110000 66982
rect 112914 66940 113222 66949
rect 112914 66938 112920 66940
rect 112976 66938 113000 66940
rect 113056 66938 113080 66940
rect 113136 66938 113160 66940
rect 113216 66938 113222 66940
rect 112976 66886 112978 66938
rect 113158 66886 113160 66938
rect 112914 66884 112920 66886
rect 112976 66884 113000 66886
rect 113056 66884 113080 66886
rect 113136 66884 113160 66886
rect 113216 66884 113222 66886
rect 112914 66875 113222 66884
rect 113650 66396 113958 66405
rect 113650 66394 113656 66396
rect 113712 66394 113736 66396
rect 113792 66394 113816 66396
rect 113872 66394 113896 66396
rect 113952 66394 113958 66396
rect 113712 66342 113714 66394
rect 113894 66342 113896 66394
rect 113650 66340 113656 66342
rect 113712 66340 113736 66342
rect 113792 66340 113816 66342
rect 113872 66340 113896 66342
rect 113952 66340 113958 66342
rect 113650 66331 113958 66340
rect 112914 65852 113222 65861
rect 112914 65850 112920 65852
rect 112976 65850 113000 65852
rect 113056 65850 113080 65852
rect 113136 65850 113160 65852
rect 113216 65850 113222 65852
rect 112976 65798 112978 65850
rect 113158 65798 113160 65850
rect 112914 65796 112920 65798
rect 112976 65796 113000 65798
rect 113056 65796 113080 65798
rect 113136 65796 113160 65798
rect 113216 65796 113222 65798
rect 112914 65787 113222 65796
rect 113650 65308 113958 65317
rect 113650 65306 113656 65308
rect 113712 65306 113736 65308
rect 113792 65306 113816 65308
rect 113872 65306 113896 65308
rect 113952 65306 113958 65308
rect 113712 65254 113714 65306
rect 113894 65254 113896 65306
rect 113650 65252 113656 65254
rect 113712 65252 113736 65254
rect 113792 65252 113816 65254
rect 113872 65252 113896 65254
rect 113952 65252 113958 65254
rect 113650 65243 113958 65252
rect 112914 64764 113222 64773
rect 112914 64762 112920 64764
rect 112976 64762 113000 64764
rect 113056 64762 113080 64764
rect 113136 64762 113160 64764
rect 113216 64762 113222 64764
rect 112976 64710 112978 64762
rect 113158 64710 113160 64762
rect 112914 64708 112920 64710
rect 112976 64708 113000 64710
rect 113056 64708 113080 64710
rect 113136 64708 113160 64710
rect 113216 64708 113222 64710
rect 112914 64699 113222 64708
rect 113650 64220 113958 64229
rect 113650 64218 113656 64220
rect 113712 64218 113736 64220
rect 113792 64218 113816 64220
rect 113872 64218 113896 64220
rect 113952 64218 113958 64220
rect 113712 64166 113714 64218
rect 113894 64166 113896 64218
rect 113650 64164 113656 64166
rect 113712 64164 113736 64166
rect 113792 64164 113816 64166
rect 113872 64164 113896 64166
rect 113952 64164 113958 64166
rect 113650 64155 113958 64164
rect 112914 63676 113222 63685
rect 112914 63674 112920 63676
rect 112976 63674 113000 63676
rect 113056 63674 113080 63676
rect 113136 63674 113160 63676
rect 113216 63674 113222 63676
rect 112976 63622 112978 63674
rect 113158 63622 113160 63674
rect 112914 63620 112920 63622
rect 112976 63620 113000 63622
rect 113056 63620 113080 63622
rect 113136 63620 113160 63622
rect 113216 63620 113222 63622
rect 112914 63611 113222 63620
rect 113650 63132 113958 63141
rect 113650 63130 113656 63132
rect 113712 63130 113736 63132
rect 113792 63130 113816 63132
rect 113872 63130 113896 63132
rect 113952 63130 113958 63132
rect 113712 63078 113714 63130
rect 113894 63078 113896 63130
rect 113650 63076 113656 63078
rect 113712 63076 113736 63078
rect 113792 63076 113816 63078
rect 113872 63076 113896 63078
rect 113952 63076 113958 63078
rect 113650 63067 113958 63076
rect 112914 62588 113222 62597
rect 112914 62586 112920 62588
rect 112976 62586 113000 62588
rect 113056 62586 113080 62588
rect 113136 62586 113160 62588
rect 113216 62586 113222 62588
rect 112976 62534 112978 62586
rect 113158 62534 113160 62586
rect 112914 62532 112920 62534
rect 112976 62532 113000 62534
rect 113056 62532 113080 62534
rect 113136 62532 113160 62534
rect 113216 62532 113222 62534
rect 112914 62523 113222 62532
rect 113650 62044 113958 62053
rect 113650 62042 113656 62044
rect 113712 62042 113736 62044
rect 113792 62042 113816 62044
rect 113872 62042 113896 62044
rect 113952 62042 113958 62044
rect 113712 61990 113714 62042
rect 113894 61990 113896 62042
rect 113650 61988 113656 61990
rect 113712 61988 113736 61990
rect 113792 61988 113816 61990
rect 113872 61988 113896 61990
rect 113952 61988 113958 61990
rect 113650 61979 113958 61988
rect 112914 61500 113222 61509
rect 112914 61498 112920 61500
rect 112976 61498 113000 61500
rect 113056 61498 113080 61500
rect 113136 61498 113160 61500
rect 113216 61498 113222 61500
rect 112976 61446 112978 61498
rect 113158 61446 113160 61498
rect 112914 61444 112920 61446
rect 112976 61444 113000 61446
rect 113056 61444 113080 61446
rect 113136 61444 113160 61446
rect 113216 61444 113222 61446
rect 112914 61435 113222 61444
rect 113650 60956 113958 60965
rect 113650 60954 113656 60956
rect 113712 60954 113736 60956
rect 113792 60954 113816 60956
rect 113872 60954 113896 60956
rect 113952 60954 113958 60956
rect 113712 60902 113714 60954
rect 113894 60902 113896 60954
rect 113650 60900 113656 60902
rect 113712 60900 113736 60902
rect 113792 60900 113816 60902
rect 113872 60900 113896 60902
rect 113952 60900 113958 60902
rect 113650 60891 113958 60900
rect 112914 60412 113222 60421
rect 112914 60410 112920 60412
rect 112976 60410 113000 60412
rect 113056 60410 113080 60412
rect 113136 60410 113160 60412
rect 113216 60410 113222 60412
rect 112976 60358 112978 60410
rect 113158 60358 113160 60410
rect 112914 60356 112920 60358
rect 112976 60356 113000 60358
rect 113056 60356 113080 60358
rect 113136 60356 113160 60358
rect 113216 60356 113222 60358
rect 112914 60347 113222 60356
rect 113650 59868 113958 59877
rect 113650 59866 113656 59868
rect 113712 59866 113736 59868
rect 113792 59866 113816 59868
rect 113872 59866 113896 59868
rect 113952 59866 113958 59868
rect 113712 59814 113714 59866
rect 113894 59814 113896 59866
rect 113650 59812 113656 59814
rect 113712 59812 113736 59814
rect 113792 59812 113816 59814
rect 113872 59812 113896 59814
rect 113952 59812 113958 59814
rect 113650 59803 113958 59812
rect 112914 59324 113222 59333
rect 112914 59322 112920 59324
rect 112976 59322 113000 59324
rect 113056 59322 113080 59324
rect 113136 59322 113160 59324
rect 113216 59322 113222 59324
rect 112976 59270 112978 59322
rect 113158 59270 113160 59322
rect 112914 59268 112920 59270
rect 112976 59268 113000 59270
rect 113056 59268 113080 59270
rect 113136 59268 113160 59270
rect 113216 59268 113222 59270
rect 112914 59259 113222 59268
rect 113650 58780 113958 58789
rect 113650 58778 113656 58780
rect 113712 58778 113736 58780
rect 113792 58778 113816 58780
rect 113872 58778 113896 58780
rect 113952 58778 113958 58780
rect 113712 58726 113714 58778
rect 113894 58726 113896 58778
rect 113650 58724 113656 58726
rect 113712 58724 113736 58726
rect 113792 58724 113816 58726
rect 113872 58724 113896 58726
rect 113952 58724 113958 58726
rect 113650 58715 113958 58724
rect 112914 58236 113222 58245
rect 112914 58234 112920 58236
rect 112976 58234 113000 58236
rect 113056 58234 113080 58236
rect 113136 58234 113160 58236
rect 113216 58234 113222 58236
rect 112976 58182 112978 58234
rect 113158 58182 113160 58234
rect 112914 58180 112920 58182
rect 112976 58180 113000 58182
rect 113056 58180 113080 58182
rect 113136 58180 113160 58182
rect 113216 58180 113222 58182
rect 112914 58171 113222 58180
rect 109960 57928 110012 57934
rect 109960 57870 110012 57876
rect 109684 57792 109736 57798
rect 109684 57734 109736 57740
rect 108684 55186 108804 55214
rect 108580 54868 108632 54874
rect 108580 54810 108632 54816
rect 108592 54670 108620 54810
rect 108580 54664 108632 54670
rect 108580 54606 108632 54612
rect 108304 54324 108356 54330
rect 108304 54266 108356 54272
rect 108316 53582 108344 54266
rect 108304 53576 108356 53582
rect 108304 53518 108356 53524
rect 108316 52154 108344 53518
rect 108592 52578 108620 54606
rect 108592 52550 108712 52578
rect 108580 52420 108632 52426
rect 108580 52362 108632 52368
rect 108304 52148 108356 52154
rect 108304 52090 108356 52096
rect 106924 52080 106976 52086
rect 106924 52022 106976 52028
rect 108316 51406 108344 52090
rect 108304 51400 108356 51406
rect 108304 51342 108356 51348
rect 108592 49434 108620 52362
rect 108684 50930 108712 52550
rect 108672 50924 108724 50930
rect 108672 50866 108724 50872
rect 108684 50522 108712 50866
rect 108672 50516 108724 50522
rect 108672 50458 108724 50464
rect 108684 50318 108712 50458
rect 108672 50312 108724 50318
rect 108672 50254 108724 50260
rect 108580 49428 108632 49434
rect 108580 49370 108632 49376
rect 108684 49366 108712 50254
rect 108672 49360 108724 49366
rect 108672 49302 108724 49308
rect 108304 49224 108356 49230
rect 108304 49166 108356 49172
rect 108316 45966 108344 49166
rect 108580 48000 108632 48006
rect 108580 47942 108632 47948
rect 108592 46578 108620 47942
rect 108776 47258 108804 55186
rect 109132 54596 109184 54602
rect 109132 54538 109184 54544
rect 109040 53440 109092 53446
rect 109040 53382 109092 53388
rect 109052 53242 109080 53382
rect 109040 53236 109092 53242
rect 109040 53178 109092 53184
rect 109052 52562 109080 53178
rect 109040 52556 109092 52562
rect 109040 52498 109092 52504
rect 109144 52426 109172 54538
rect 109972 53446 110000 57870
rect 113650 57692 113958 57701
rect 113650 57690 113656 57692
rect 113712 57690 113736 57692
rect 113792 57690 113816 57692
rect 113872 57690 113896 57692
rect 113952 57690 113958 57692
rect 113712 57638 113714 57690
rect 113894 57638 113896 57690
rect 113650 57636 113656 57638
rect 113712 57636 113736 57638
rect 113792 57636 113816 57638
rect 113872 57636 113896 57638
rect 113952 57636 113958 57638
rect 113650 57627 113958 57636
rect 112914 57148 113222 57157
rect 112914 57146 112920 57148
rect 112976 57146 113000 57148
rect 113056 57146 113080 57148
rect 113136 57146 113160 57148
rect 113216 57146 113222 57148
rect 112976 57094 112978 57146
rect 113158 57094 113160 57146
rect 112914 57092 112920 57094
rect 112976 57092 113000 57094
rect 113056 57092 113080 57094
rect 113136 57092 113160 57094
rect 113216 57092 113222 57094
rect 112914 57083 113222 57092
rect 113650 56604 113958 56613
rect 113650 56602 113656 56604
rect 113712 56602 113736 56604
rect 113792 56602 113816 56604
rect 113872 56602 113896 56604
rect 113952 56602 113958 56604
rect 113712 56550 113714 56602
rect 113894 56550 113896 56602
rect 113650 56548 113656 56550
rect 113712 56548 113736 56550
rect 113792 56548 113816 56550
rect 113872 56548 113896 56550
rect 113952 56548 113958 56550
rect 113650 56539 113958 56548
rect 112914 56060 113222 56069
rect 112914 56058 112920 56060
rect 112976 56058 113000 56060
rect 113056 56058 113080 56060
rect 113136 56058 113160 56060
rect 113216 56058 113222 56060
rect 112976 56006 112978 56058
rect 113158 56006 113160 56058
rect 112914 56004 112920 56006
rect 112976 56004 113000 56006
rect 113056 56004 113080 56006
rect 113136 56004 113160 56006
rect 113216 56004 113222 56006
rect 112914 55995 113222 56004
rect 113650 55516 113958 55525
rect 113650 55514 113656 55516
rect 113712 55514 113736 55516
rect 113792 55514 113816 55516
rect 113872 55514 113896 55516
rect 113952 55514 113958 55516
rect 113712 55462 113714 55514
rect 113894 55462 113896 55514
rect 113650 55460 113656 55462
rect 113712 55460 113736 55462
rect 113792 55460 113816 55462
rect 113872 55460 113896 55462
rect 113952 55460 113958 55462
rect 113650 55451 113958 55460
rect 112914 54972 113222 54981
rect 112914 54970 112920 54972
rect 112976 54970 113000 54972
rect 113056 54970 113080 54972
rect 113136 54970 113160 54972
rect 113216 54970 113222 54972
rect 112976 54918 112978 54970
rect 113158 54918 113160 54970
rect 112914 54916 112920 54918
rect 112976 54916 113000 54918
rect 113056 54916 113080 54918
rect 113136 54916 113160 54918
rect 113216 54916 113222 54918
rect 112914 54907 113222 54916
rect 113650 54428 113958 54437
rect 113650 54426 113656 54428
rect 113712 54426 113736 54428
rect 113792 54426 113816 54428
rect 113872 54426 113896 54428
rect 113952 54426 113958 54428
rect 113712 54374 113714 54426
rect 113894 54374 113896 54426
rect 113650 54372 113656 54374
rect 113712 54372 113736 54374
rect 113792 54372 113816 54374
rect 113872 54372 113896 54374
rect 113952 54372 113958 54374
rect 113650 54363 113958 54372
rect 112914 53884 113222 53893
rect 112914 53882 112920 53884
rect 112976 53882 113000 53884
rect 113056 53882 113080 53884
rect 113136 53882 113160 53884
rect 113216 53882 113222 53884
rect 112976 53830 112978 53882
rect 113158 53830 113160 53882
rect 112914 53828 112920 53830
rect 112976 53828 113000 53830
rect 113056 53828 113080 53830
rect 113136 53828 113160 53830
rect 113216 53828 113222 53830
rect 112914 53819 113222 53828
rect 109960 53440 110012 53446
rect 109960 53382 110012 53388
rect 110696 53440 110748 53446
rect 110696 53382 110748 53388
rect 110708 52494 110736 53382
rect 113650 53340 113958 53349
rect 113650 53338 113656 53340
rect 113712 53338 113736 53340
rect 113792 53338 113816 53340
rect 113872 53338 113896 53340
rect 113952 53338 113958 53340
rect 113712 53286 113714 53338
rect 113894 53286 113896 53338
rect 113650 53284 113656 53286
rect 113712 53284 113736 53286
rect 113792 53284 113816 53286
rect 113872 53284 113896 53286
rect 113952 53284 113958 53286
rect 113650 53275 113958 53284
rect 112914 52796 113222 52805
rect 112914 52794 112920 52796
rect 112976 52794 113000 52796
rect 113056 52794 113080 52796
rect 113136 52794 113160 52796
rect 113216 52794 113222 52796
rect 112976 52742 112978 52794
rect 113158 52742 113160 52794
rect 112914 52740 112920 52742
rect 112976 52740 113000 52742
rect 113056 52740 113080 52742
rect 113136 52740 113160 52742
rect 113216 52740 113222 52742
rect 112914 52731 113222 52740
rect 110696 52488 110748 52494
rect 110696 52430 110748 52436
rect 109132 52420 109184 52426
rect 109132 52362 109184 52368
rect 109408 52352 109460 52358
rect 109408 52294 109460 52300
rect 109420 52018 109448 52294
rect 109408 52012 109460 52018
rect 109408 51954 109460 51960
rect 108948 50720 109000 50726
rect 108948 50662 109000 50668
rect 108960 48142 108988 50662
rect 109132 50244 109184 50250
rect 109132 50186 109184 50192
rect 109040 49156 109092 49162
rect 109040 49098 109092 49104
rect 108948 48136 109000 48142
rect 108948 48078 109000 48084
rect 108764 47252 108816 47258
rect 108764 47194 108816 47200
rect 108580 46572 108632 46578
rect 108580 46514 108632 46520
rect 108304 45960 108356 45966
rect 108304 45902 108356 45908
rect 108316 45626 108344 45902
rect 108488 45824 108540 45830
rect 108488 45766 108540 45772
rect 108304 45620 108356 45626
rect 108304 45562 108356 45568
rect 108316 44402 108344 45562
rect 108304 44396 108356 44402
rect 108304 44338 108356 44344
rect 9678 44202 9734 44211
rect 9678 44140 9680 44146
rect 9732 44140 9734 44146
rect 9678 44137 9734 44140
rect 9680 44134 9732 44137
rect 108316 43994 108344 44338
rect 108304 43988 108356 43994
rect 108304 43930 108356 43936
rect 108316 43790 108344 43930
rect 108500 43874 108528 45766
rect 108592 45490 108620 46514
rect 109052 45966 109080 49098
rect 109144 46986 109172 50186
rect 109420 49162 109448 51954
rect 109592 51264 109644 51270
rect 109592 51206 109644 51212
rect 109604 50998 109632 51206
rect 109592 50992 109644 50998
rect 109592 50934 109644 50940
rect 109500 49360 109552 49366
rect 109500 49302 109552 49308
rect 109408 49156 109460 49162
rect 109408 49098 109460 49104
rect 109132 46980 109184 46986
rect 109132 46922 109184 46928
rect 109040 45960 109092 45966
rect 109040 45902 109092 45908
rect 109224 45824 109276 45830
rect 109224 45766 109276 45772
rect 108580 45484 108632 45490
rect 108580 45426 108632 45432
rect 109132 45280 109184 45286
rect 109132 45222 109184 45228
rect 108856 44260 108908 44266
rect 108856 44202 108908 44208
rect 108500 43846 108620 43874
rect 108304 43784 108356 43790
rect 108304 43726 108356 43732
rect 9680 43172 9732 43178
rect 9680 43114 9732 43120
rect 9692 42987 9720 43114
rect 9678 42978 9734 42987
rect 9678 42913 9734 42922
rect 108316 42906 108344 43726
rect 108304 42900 108356 42906
rect 108304 42842 108356 42848
rect 108316 41818 108344 42842
rect 108488 42560 108540 42566
rect 108488 42502 108540 42508
rect 108304 41812 108356 41818
rect 108304 41754 108356 41760
rect 108316 41614 108344 41754
rect 108304 41608 108356 41614
rect 108304 41550 108356 41556
rect 108396 41472 108448 41478
rect 108396 41414 108448 41420
rect 9678 41210 9734 41219
rect 9678 41145 9734 41154
rect 9692 41002 9720 41145
rect 9680 40996 9732 41002
rect 9680 40938 9732 40944
rect 9680 40452 9732 40458
rect 9680 40394 9732 40400
rect 9692 40131 9720 40394
rect 9678 40122 9734 40131
rect 9678 40057 9734 40066
rect 106924 39364 106976 39370
rect 106924 39306 106976 39312
rect 9678 38490 9734 38499
rect 9678 38425 9734 38434
rect 9692 38282 9720 38425
rect 9680 38276 9732 38282
rect 9680 38218 9732 38224
rect 9496 37732 9548 37738
rect 9496 37674 9548 37680
rect 9508 37547 9536 37674
rect 9494 37538 9550 37547
rect 9494 37473 9550 37482
rect 9494 35770 9550 35779
rect 9494 35708 9496 35714
rect 9548 35708 9550 35714
rect 9494 35705 9550 35708
rect 9496 35702 9548 35705
rect 106936 26625 106964 39306
rect 108212 39296 108264 39302
rect 108212 39238 108264 39244
rect 107016 37324 107068 37330
rect 107016 37266 107068 37272
rect 106922 26616 106978 26625
rect 106922 26551 106978 26560
rect 107028 24993 107056 37266
rect 107108 36168 107160 36174
rect 107108 36110 107160 36116
rect 107014 24984 107070 24993
rect 107014 24919 107070 24928
rect 107120 23633 107148 36110
rect 108224 34678 108252 39238
rect 108408 36854 108436 41414
rect 108500 38282 108528 42502
rect 108592 42294 108620 43846
rect 108672 43716 108724 43722
rect 108672 43658 108724 43664
rect 108580 42288 108632 42294
rect 108580 42230 108632 42236
rect 108580 40452 108632 40458
rect 108580 40394 108632 40400
rect 108488 38276 108540 38282
rect 108488 38218 108540 38224
rect 108592 38010 108620 40394
rect 108684 39370 108712 43658
rect 108764 41132 108816 41138
rect 108764 41074 108816 41080
rect 108672 39364 108724 39370
rect 108672 39306 108724 39312
rect 108672 38208 108724 38214
rect 108672 38150 108724 38156
rect 108580 38004 108632 38010
rect 108580 37946 108632 37952
rect 108488 37460 108540 37466
rect 108488 37402 108540 37408
rect 108396 36848 108448 36854
rect 108396 36790 108448 36796
rect 108304 36576 108356 36582
rect 108304 36518 108356 36524
rect 108212 34672 108264 34678
rect 108212 34614 108264 34620
rect 108316 33522 108344 36518
rect 108396 35556 108448 35562
rect 108396 35498 108448 35504
rect 108304 33516 108356 33522
rect 108304 33458 108356 33464
rect 108316 33046 108344 33458
rect 108304 33040 108356 33046
rect 108304 32982 108356 32988
rect 108304 32904 108356 32910
rect 108408 32892 108436 35498
rect 108500 34746 108528 37402
rect 108684 34762 108712 38150
rect 108776 37890 108804 41074
rect 108868 40458 108896 44202
rect 109144 43382 109172 45222
rect 109132 43376 109184 43382
rect 109132 43318 109184 43324
rect 109236 43314 109264 45766
rect 109420 45642 109448 49098
rect 109512 45778 109540 49302
rect 109604 48210 109632 50934
rect 109592 48204 109644 48210
rect 109592 48146 109644 48152
rect 110328 48204 110380 48210
rect 110328 48146 110380 48152
rect 110052 48068 110104 48074
rect 110052 48010 110104 48016
rect 109684 46368 109736 46374
rect 109684 46310 109736 46316
rect 109512 45750 109632 45778
rect 109420 45614 109540 45642
rect 109512 45558 109540 45614
rect 109316 45552 109368 45558
rect 109316 45494 109368 45500
rect 109408 45552 109460 45558
rect 109408 45494 109460 45500
rect 109500 45552 109552 45558
rect 109500 45494 109552 45500
rect 109328 45082 109356 45494
rect 109316 45076 109368 45082
rect 109316 45018 109368 45024
rect 109420 43722 109448 45494
rect 109512 44878 109540 45494
rect 109604 45490 109632 45750
rect 109696 45490 109724 46310
rect 109592 45484 109644 45490
rect 109592 45426 109644 45432
rect 109684 45484 109736 45490
rect 109684 45426 109736 45432
rect 110064 45422 110092 48010
rect 110340 47138 110368 48146
rect 110512 47252 110564 47258
rect 110512 47194 110564 47200
rect 110340 47122 110460 47138
rect 110340 47116 110472 47122
rect 110340 47110 110420 47116
rect 110144 46980 110196 46986
rect 110144 46922 110196 46928
rect 110052 45416 110104 45422
rect 110052 45358 110104 45364
rect 109592 45280 109644 45286
rect 109592 45222 109644 45228
rect 109604 44878 109632 45222
rect 109500 44872 109552 44878
rect 109500 44814 109552 44820
rect 109592 44872 109644 44878
rect 109592 44814 109644 44820
rect 109408 43716 109460 43722
rect 109408 43658 109460 43664
rect 109224 43308 109276 43314
rect 109224 43250 109276 43256
rect 108948 41676 109000 41682
rect 108948 41618 109000 41624
rect 108960 41138 108988 41618
rect 108948 41132 109000 41138
rect 108948 41074 109000 41080
rect 108948 40996 109000 41002
rect 108948 40938 109000 40944
rect 108960 40594 108988 40938
rect 108948 40588 109000 40594
rect 108948 40530 109000 40536
rect 108856 40452 108908 40458
rect 108856 40394 108908 40400
rect 108960 38486 108988 40530
rect 108948 38480 109000 38486
rect 108948 38422 109000 38428
rect 109420 37942 109448 43658
rect 109512 43330 109540 44814
rect 110156 43994 110184 46922
rect 110340 46170 110368 47110
rect 110420 47058 110472 47064
rect 110328 46164 110380 46170
rect 110328 46106 110380 46112
rect 110144 43988 110196 43994
rect 110144 43930 110196 43936
rect 110236 43988 110288 43994
rect 110236 43930 110288 43936
rect 109684 43852 109736 43858
rect 109684 43794 109736 43800
rect 109512 43314 109632 43330
rect 109512 43308 109644 43314
rect 109512 43302 109592 43308
rect 109512 42702 109540 43302
rect 109592 43250 109644 43256
rect 109592 43104 109644 43110
rect 109592 43046 109644 43052
rect 109500 42696 109552 42702
rect 109500 42638 109552 42644
rect 109512 42106 109540 42638
rect 109604 42634 109632 43046
rect 109592 42628 109644 42634
rect 109592 42570 109644 42576
rect 109512 42078 109632 42106
rect 109500 42016 109552 42022
rect 109500 41958 109552 41964
rect 109512 40050 109540 41958
rect 109604 41546 109632 42078
rect 109592 41540 109644 41546
rect 109592 41482 109644 41488
rect 109604 40050 109632 41482
rect 109696 41414 109724 43794
rect 109776 43784 109828 43790
rect 109776 43726 109828 43732
rect 109788 41818 109816 43726
rect 109868 43648 109920 43654
rect 109868 43590 109920 43596
rect 109880 42906 109908 43590
rect 110248 43450 110276 43930
rect 110236 43444 110288 43450
rect 110236 43386 110288 43392
rect 110144 43308 110196 43314
rect 110144 43250 110196 43256
rect 109960 43172 110012 43178
rect 109960 43114 110012 43120
rect 109868 42900 109920 42906
rect 109868 42842 109920 42848
rect 109868 42628 109920 42634
rect 109868 42570 109920 42576
rect 109776 41812 109828 41818
rect 109776 41754 109828 41760
rect 109696 41386 109816 41414
rect 109684 41132 109736 41138
rect 109684 41074 109736 41080
rect 109696 40662 109724 41074
rect 109684 40656 109736 40662
rect 109684 40598 109736 40604
rect 109788 40610 109816 41386
rect 109880 41138 109908 42570
rect 109868 41132 109920 41138
rect 109868 41074 109920 41080
rect 109696 40050 109724 40598
rect 109788 40582 109908 40610
rect 109880 40526 109908 40582
rect 109868 40520 109920 40526
rect 109868 40462 109920 40468
rect 109500 40044 109552 40050
rect 109500 39986 109552 39992
rect 109592 40044 109644 40050
rect 109592 39986 109644 39992
rect 109684 40044 109736 40050
rect 109684 39986 109736 39992
rect 109512 39098 109540 39986
rect 109604 39098 109632 39986
rect 109776 39636 109828 39642
rect 109776 39578 109828 39584
rect 109684 39364 109736 39370
rect 109684 39306 109736 39312
rect 109500 39092 109552 39098
rect 109500 39034 109552 39040
rect 109592 39092 109644 39098
rect 109592 39034 109644 39040
rect 109592 38820 109644 38826
rect 109592 38762 109644 38768
rect 109316 37936 109368 37942
rect 108776 37862 108896 37890
rect 109316 37878 109368 37884
rect 109408 37936 109460 37942
rect 109408 37878 109460 37884
rect 108764 37732 108816 37738
rect 108764 37674 108816 37680
rect 108776 35834 108804 37674
rect 108868 37466 108896 37862
rect 108856 37460 108908 37466
rect 108856 37402 108908 37408
rect 108856 37120 108908 37126
rect 108856 37062 108908 37068
rect 108764 35828 108816 35834
rect 108764 35770 108816 35776
rect 108764 35080 108816 35086
rect 108764 35022 108816 35028
rect 108488 34740 108540 34746
rect 108488 34682 108540 34688
rect 108592 34734 108712 34762
rect 108592 34610 108620 34734
rect 108776 34610 108804 35022
rect 108488 34604 108540 34610
rect 108488 34546 108540 34552
rect 108580 34604 108632 34610
rect 108764 34604 108816 34610
rect 108580 34546 108632 34552
rect 108684 34564 108764 34592
rect 108500 33998 108528 34546
rect 108592 33998 108620 34546
rect 108488 33992 108540 33998
rect 108488 33934 108540 33940
rect 108580 33992 108632 33998
rect 108580 33934 108632 33940
rect 108500 33658 108528 33934
rect 108488 33652 108540 33658
rect 108488 33594 108540 33600
rect 108684 33522 108712 34564
rect 108764 34546 108816 34552
rect 108868 34202 108896 37062
rect 109040 36100 109092 36106
rect 109040 36042 109092 36048
rect 109052 35850 109080 36042
rect 109224 36032 109276 36038
rect 109224 35974 109276 35980
rect 108960 35834 109080 35850
rect 108948 35828 109080 35834
rect 109000 35822 109080 35828
rect 108948 35770 109000 35776
rect 109040 35760 109092 35766
rect 108960 35708 109040 35714
rect 108960 35702 109092 35708
rect 108960 35686 109080 35702
rect 108856 34196 108908 34202
rect 108856 34138 108908 34144
rect 108764 33924 108816 33930
rect 108764 33866 108816 33872
rect 108672 33516 108724 33522
rect 108672 33458 108724 33464
rect 108356 32864 108436 32892
rect 108304 32846 108356 32852
rect 108408 32570 108436 32864
rect 108684 32570 108712 33458
rect 108396 32564 108448 32570
rect 108396 32506 108448 32512
rect 108672 32564 108724 32570
rect 108672 32506 108724 32512
rect 108488 32224 108540 32230
rect 108488 32166 108540 32172
rect 108500 31822 108528 32166
rect 108776 31890 108804 33866
rect 108960 33402 108988 35686
rect 109040 35488 109092 35494
rect 109040 35430 109092 35436
rect 109052 35290 109080 35430
rect 109040 35284 109092 35290
rect 109040 35226 109092 35232
rect 109236 34746 109264 35974
rect 109328 35834 109356 37878
rect 109420 37262 109448 37878
rect 109408 37256 109460 37262
rect 109408 37198 109460 37204
rect 109408 36372 109460 36378
rect 109408 36314 109460 36320
rect 109316 35828 109368 35834
rect 109316 35770 109368 35776
rect 109420 34746 109448 36314
rect 109604 35698 109632 38762
rect 109696 36378 109724 39306
rect 109788 39030 109816 39578
rect 109776 39024 109828 39030
rect 109776 38966 109828 38972
rect 109880 38010 109908 40462
rect 109972 40050 110000 43114
rect 110156 43110 110184 43250
rect 110144 43104 110196 43110
rect 110144 43046 110196 43052
rect 110156 42702 110184 43046
rect 110144 42696 110196 42702
rect 110144 42638 110196 42644
rect 110340 42226 110368 46106
rect 110420 45892 110472 45898
rect 110420 45834 110472 45840
rect 110432 43994 110460 45834
rect 110420 43988 110472 43994
rect 110420 43930 110472 43936
rect 110328 42220 110380 42226
rect 110328 42162 110380 42168
rect 110052 42152 110104 42158
rect 110052 42094 110104 42100
rect 110064 40730 110092 42094
rect 110236 41608 110288 41614
rect 110236 41550 110288 41556
rect 110248 41138 110276 41550
rect 110236 41132 110288 41138
rect 110236 41074 110288 41080
rect 110340 41002 110368 42162
rect 110524 41682 110552 47194
rect 110512 41676 110564 41682
rect 110512 41618 110564 41624
rect 110524 41414 110552 41618
rect 110604 41540 110656 41546
rect 110604 41482 110656 41488
rect 110432 41386 110552 41414
rect 110328 40996 110380 41002
rect 110328 40938 110380 40944
rect 110236 40928 110288 40934
rect 110236 40870 110288 40876
rect 110052 40724 110104 40730
rect 110052 40666 110104 40672
rect 110144 40384 110196 40390
rect 110144 40326 110196 40332
rect 110156 40186 110184 40326
rect 110144 40180 110196 40186
rect 110144 40122 110196 40128
rect 109960 40044 110012 40050
rect 109960 39986 110012 39992
rect 109972 38962 110000 39986
rect 110144 39840 110196 39846
rect 110144 39782 110196 39788
rect 109960 38956 110012 38962
rect 109960 38898 110012 38904
rect 110156 38842 110184 39782
rect 110248 39642 110276 40870
rect 110328 40724 110380 40730
rect 110328 40666 110380 40672
rect 110236 39636 110288 39642
rect 110236 39578 110288 39584
rect 110248 39370 110276 39578
rect 110236 39364 110288 39370
rect 110236 39306 110288 39312
rect 110340 39098 110368 40666
rect 110432 40186 110460 41386
rect 110616 41138 110644 41482
rect 110604 41132 110656 41138
rect 110604 41074 110656 41080
rect 110512 40928 110564 40934
rect 110512 40870 110564 40876
rect 110420 40180 110472 40186
rect 110420 40122 110472 40128
rect 110432 39982 110460 40122
rect 110524 40118 110552 40870
rect 110616 40662 110644 41074
rect 110604 40656 110656 40662
rect 110604 40598 110656 40604
rect 110604 40384 110656 40390
rect 110604 40326 110656 40332
rect 110512 40112 110564 40118
rect 110512 40054 110564 40060
rect 110420 39976 110472 39982
rect 110420 39918 110472 39924
rect 110432 39658 110460 39918
rect 110432 39630 110552 39658
rect 110420 39500 110472 39506
rect 110420 39442 110472 39448
rect 110328 39092 110380 39098
rect 110328 39034 110380 39040
rect 110156 38814 110276 38842
rect 110144 38752 110196 38758
rect 110144 38694 110196 38700
rect 110052 38276 110104 38282
rect 110052 38218 110104 38224
rect 109868 38004 109920 38010
rect 109868 37946 109920 37952
rect 109776 36712 109828 36718
rect 109776 36654 109828 36660
rect 109684 36372 109736 36378
rect 109684 36314 109736 36320
rect 109788 35766 109816 36654
rect 109880 36106 109908 37946
rect 109960 37664 110012 37670
rect 109960 37606 110012 37612
rect 109972 37346 110000 37606
rect 110064 37466 110092 38218
rect 110156 37942 110184 38694
rect 110144 37936 110196 37942
rect 110144 37878 110196 37884
rect 110052 37460 110104 37466
rect 110052 37402 110104 37408
rect 109972 37318 110092 37346
rect 109960 37188 110012 37194
rect 109960 37130 110012 37136
rect 109868 36100 109920 36106
rect 109868 36042 109920 36048
rect 109776 35760 109828 35766
rect 109776 35702 109828 35708
rect 109592 35692 109644 35698
rect 109592 35634 109644 35640
rect 109604 35562 109632 35634
rect 109592 35556 109644 35562
rect 109592 35498 109644 35504
rect 109500 35488 109552 35494
rect 109500 35430 109552 35436
rect 109224 34740 109276 34746
rect 109224 34682 109276 34688
rect 109408 34740 109460 34746
rect 109408 34682 109460 34688
rect 109040 34604 109092 34610
rect 109040 34546 109092 34552
rect 109052 33998 109080 34546
rect 109040 33992 109092 33998
rect 109040 33934 109092 33940
rect 109224 33856 109276 33862
rect 109224 33798 109276 33804
rect 109236 33590 109264 33798
rect 109224 33584 109276 33590
rect 109224 33526 109276 33532
rect 109132 33516 109184 33522
rect 109132 33458 109184 33464
rect 108868 33374 108988 33402
rect 108868 33114 108896 33374
rect 108948 33312 109000 33318
rect 108948 33254 109000 33260
rect 108856 33108 108908 33114
rect 108856 33050 108908 33056
rect 108960 32434 108988 33254
rect 109144 33114 109172 33458
rect 109132 33108 109184 33114
rect 109132 33050 109184 33056
rect 109236 32910 109264 33526
rect 109408 33312 109460 33318
rect 109406 33280 109408 33289
rect 109460 33280 109462 33289
rect 109406 33215 109462 33224
rect 109224 32904 109276 32910
rect 109224 32846 109276 32852
rect 109408 32768 109460 32774
rect 109512 32722 109540 35430
rect 109972 34678 110000 37130
rect 110064 35306 110092 37318
rect 110156 37262 110184 37878
rect 110144 37256 110196 37262
rect 110144 37198 110196 37204
rect 110248 36174 110276 38814
rect 110328 37800 110380 37806
rect 110328 37742 110380 37748
rect 110236 36168 110288 36174
rect 110236 36110 110288 36116
rect 110064 35278 110184 35306
rect 109960 34672 110012 34678
rect 109960 34614 110012 34620
rect 109960 34536 110012 34542
rect 109960 34478 110012 34484
rect 109868 34400 109920 34406
rect 109868 34342 109920 34348
rect 109592 34196 109644 34202
rect 109592 34138 109644 34144
rect 109604 33386 109632 34138
rect 109880 33998 109908 34342
rect 109972 34082 110000 34478
rect 110156 34406 110184 35278
rect 110340 34542 110368 37742
rect 110432 36922 110460 39442
rect 110524 39098 110552 39630
rect 110512 39092 110564 39098
rect 110512 39034 110564 39040
rect 110616 37992 110644 40326
rect 110708 39642 110736 52430
rect 113650 52252 113958 52261
rect 113650 52250 113656 52252
rect 113712 52250 113736 52252
rect 113792 52250 113816 52252
rect 113872 52250 113896 52252
rect 113952 52250 113958 52252
rect 113712 52198 113714 52250
rect 113894 52198 113896 52250
rect 113650 52196 113656 52198
rect 113712 52196 113736 52198
rect 113792 52196 113816 52198
rect 113872 52196 113896 52198
rect 113952 52196 113958 52198
rect 113650 52187 113958 52196
rect 112914 51708 113222 51717
rect 112914 51706 112920 51708
rect 112976 51706 113000 51708
rect 113056 51706 113080 51708
rect 113136 51706 113160 51708
rect 113216 51706 113222 51708
rect 112976 51654 112978 51706
rect 113158 51654 113160 51706
rect 112914 51652 112920 51654
rect 112976 51652 113000 51654
rect 113056 51652 113080 51654
rect 113136 51652 113160 51654
rect 113216 51652 113222 51654
rect 112914 51643 113222 51652
rect 113650 51164 113958 51173
rect 113650 51162 113656 51164
rect 113712 51162 113736 51164
rect 113792 51162 113816 51164
rect 113872 51162 113896 51164
rect 113952 51162 113958 51164
rect 113712 51110 113714 51162
rect 113894 51110 113896 51162
rect 113650 51108 113656 51110
rect 113712 51108 113736 51110
rect 113792 51108 113816 51110
rect 113872 51108 113896 51110
rect 113952 51108 113958 51110
rect 113650 51099 113958 51108
rect 112914 50620 113222 50629
rect 112914 50618 112920 50620
rect 112976 50618 113000 50620
rect 113056 50618 113080 50620
rect 113136 50618 113160 50620
rect 113216 50618 113222 50620
rect 112976 50566 112978 50618
rect 113158 50566 113160 50618
rect 112914 50564 112920 50566
rect 112976 50564 113000 50566
rect 113056 50564 113080 50566
rect 113136 50564 113160 50566
rect 113216 50564 113222 50566
rect 112914 50555 113222 50564
rect 113650 50076 113958 50085
rect 113650 50074 113656 50076
rect 113712 50074 113736 50076
rect 113792 50074 113816 50076
rect 113872 50074 113896 50076
rect 113952 50074 113958 50076
rect 113712 50022 113714 50074
rect 113894 50022 113896 50074
rect 113650 50020 113656 50022
rect 113712 50020 113736 50022
rect 113792 50020 113816 50022
rect 113872 50020 113896 50022
rect 113952 50020 113958 50022
rect 113650 50011 113958 50020
rect 112914 49532 113222 49541
rect 112914 49530 112920 49532
rect 112976 49530 113000 49532
rect 113056 49530 113080 49532
rect 113136 49530 113160 49532
rect 113216 49530 113222 49532
rect 112976 49478 112978 49530
rect 113158 49478 113160 49530
rect 112914 49476 112920 49478
rect 112976 49476 113000 49478
rect 113056 49476 113080 49478
rect 113136 49476 113160 49478
rect 113216 49476 113222 49478
rect 112914 49467 113222 49476
rect 113650 48988 113958 48997
rect 113650 48986 113656 48988
rect 113712 48986 113736 48988
rect 113792 48986 113816 48988
rect 113872 48986 113896 48988
rect 113952 48986 113958 48988
rect 113712 48934 113714 48986
rect 113894 48934 113896 48986
rect 113650 48932 113656 48934
rect 113712 48932 113736 48934
rect 113792 48932 113816 48934
rect 113872 48932 113896 48934
rect 113952 48932 113958 48934
rect 113650 48923 113958 48932
rect 112914 48444 113222 48453
rect 112914 48442 112920 48444
rect 112976 48442 113000 48444
rect 113056 48442 113080 48444
rect 113136 48442 113160 48444
rect 113216 48442 113222 48444
rect 112976 48390 112978 48442
rect 113158 48390 113160 48442
rect 112914 48388 112920 48390
rect 112976 48388 113000 48390
rect 113056 48388 113080 48390
rect 113136 48388 113160 48390
rect 113216 48388 113222 48390
rect 112914 48379 113222 48388
rect 113650 47900 113958 47909
rect 113650 47898 113656 47900
rect 113712 47898 113736 47900
rect 113792 47898 113816 47900
rect 113872 47898 113896 47900
rect 113952 47898 113958 47900
rect 113712 47846 113714 47898
rect 113894 47846 113896 47898
rect 113650 47844 113656 47846
rect 113712 47844 113736 47846
rect 113792 47844 113816 47846
rect 113872 47844 113896 47846
rect 113952 47844 113958 47846
rect 113650 47835 113958 47844
rect 112914 47356 113222 47365
rect 112914 47354 112920 47356
rect 112976 47354 113000 47356
rect 113056 47354 113080 47356
rect 113136 47354 113160 47356
rect 113216 47354 113222 47356
rect 112976 47302 112978 47354
rect 113158 47302 113160 47354
rect 112914 47300 112920 47302
rect 112976 47300 113000 47302
rect 113056 47300 113080 47302
rect 113136 47300 113160 47302
rect 113216 47300 113222 47302
rect 112914 47291 113222 47300
rect 113650 46812 113958 46821
rect 113650 46810 113656 46812
rect 113712 46810 113736 46812
rect 113792 46810 113816 46812
rect 113872 46810 113896 46812
rect 113952 46810 113958 46812
rect 113712 46758 113714 46810
rect 113894 46758 113896 46810
rect 113650 46756 113656 46758
rect 113712 46756 113736 46758
rect 113792 46756 113816 46758
rect 113872 46756 113896 46758
rect 113952 46756 113958 46758
rect 113650 46747 113958 46756
rect 112914 46268 113222 46277
rect 112914 46266 112920 46268
rect 112976 46266 113000 46268
rect 113056 46266 113080 46268
rect 113136 46266 113160 46268
rect 113216 46266 113222 46268
rect 112976 46214 112978 46266
rect 113158 46214 113160 46266
rect 112914 46212 112920 46214
rect 112976 46212 113000 46214
rect 113056 46212 113080 46214
rect 113136 46212 113160 46214
rect 113216 46212 113222 46214
rect 112914 46203 113222 46212
rect 113650 45724 113958 45733
rect 113650 45722 113656 45724
rect 113712 45722 113736 45724
rect 113792 45722 113816 45724
rect 113872 45722 113896 45724
rect 113952 45722 113958 45724
rect 113712 45670 113714 45722
rect 113894 45670 113896 45722
rect 113650 45668 113656 45670
rect 113712 45668 113736 45670
rect 113792 45668 113816 45670
rect 113872 45668 113896 45670
rect 113952 45668 113958 45670
rect 113650 45659 113958 45668
rect 112914 45180 113222 45189
rect 112914 45178 112920 45180
rect 112976 45178 113000 45180
rect 113056 45178 113080 45180
rect 113136 45178 113160 45180
rect 113216 45178 113222 45180
rect 112976 45126 112978 45178
rect 113158 45126 113160 45178
rect 112914 45124 112920 45126
rect 112976 45124 113000 45126
rect 113056 45124 113080 45126
rect 113136 45124 113160 45126
rect 113216 45124 113222 45126
rect 112914 45115 113222 45124
rect 113650 44636 113958 44645
rect 113650 44634 113656 44636
rect 113712 44634 113736 44636
rect 113792 44634 113816 44636
rect 113872 44634 113896 44636
rect 113952 44634 113958 44636
rect 113712 44582 113714 44634
rect 113894 44582 113896 44634
rect 113650 44580 113656 44582
rect 113712 44580 113736 44582
rect 113792 44580 113816 44582
rect 113872 44580 113896 44582
rect 113952 44580 113958 44582
rect 113650 44571 113958 44580
rect 112914 44092 113222 44101
rect 112914 44090 112920 44092
rect 112976 44090 113000 44092
rect 113056 44090 113080 44092
rect 113136 44090 113160 44092
rect 113216 44090 113222 44092
rect 112976 44038 112978 44090
rect 113158 44038 113160 44090
rect 112914 44036 112920 44038
rect 112976 44036 113000 44038
rect 113056 44036 113080 44038
rect 113136 44036 113160 44038
rect 113216 44036 113222 44038
rect 112914 44027 113222 44036
rect 113650 43548 113958 43557
rect 113650 43546 113656 43548
rect 113712 43546 113736 43548
rect 113792 43546 113816 43548
rect 113872 43546 113896 43548
rect 113952 43546 113958 43548
rect 113712 43494 113714 43546
rect 113894 43494 113896 43546
rect 113650 43492 113656 43494
rect 113712 43492 113736 43494
rect 113792 43492 113816 43494
rect 113872 43492 113896 43494
rect 113952 43492 113958 43494
rect 113650 43483 113958 43492
rect 112914 43004 113222 43013
rect 112914 43002 112920 43004
rect 112976 43002 113000 43004
rect 113056 43002 113080 43004
rect 113136 43002 113160 43004
rect 113216 43002 113222 43004
rect 112976 42950 112978 43002
rect 113158 42950 113160 43002
rect 112914 42948 112920 42950
rect 112976 42948 113000 42950
rect 113056 42948 113080 42950
rect 113136 42948 113160 42950
rect 113216 42948 113222 42950
rect 112914 42939 113222 42948
rect 113650 42460 113958 42469
rect 113650 42458 113656 42460
rect 113712 42458 113736 42460
rect 113792 42458 113816 42460
rect 113872 42458 113896 42460
rect 113952 42458 113958 42460
rect 113712 42406 113714 42458
rect 113894 42406 113896 42458
rect 113650 42404 113656 42406
rect 113712 42404 113736 42406
rect 113792 42404 113816 42406
rect 113872 42404 113896 42406
rect 113952 42404 113958 42406
rect 113650 42395 113958 42404
rect 112914 41916 113222 41925
rect 112914 41914 112920 41916
rect 112976 41914 113000 41916
rect 113056 41914 113080 41916
rect 113136 41914 113160 41916
rect 113216 41914 113222 41916
rect 112976 41862 112978 41914
rect 113158 41862 113160 41914
rect 112914 41860 112920 41862
rect 112976 41860 113000 41862
rect 113056 41860 113080 41862
rect 113136 41860 113160 41862
rect 113216 41860 113222 41862
rect 112914 41851 113222 41860
rect 110788 41472 110840 41478
rect 110788 41414 110840 41420
rect 110800 40186 110828 41414
rect 113650 41372 113958 41381
rect 113650 41370 113656 41372
rect 113712 41370 113736 41372
rect 113792 41370 113816 41372
rect 113872 41370 113896 41372
rect 113952 41370 113958 41372
rect 113712 41318 113714 41370
rect 113894 41318 113896 41370
rect 113650 41316 113656 41318
rect 113712 41316 113736 41318
rect 113792 41316 113816 41318
rect 113872 41316 113896 41318
rect 113952 41316 113958 41318
rect 113650 41307 113958 41316
rect 110880 41132 110932 41138
rect 110880 41074 110932 41080
rect 110788 40180 110840 40186
rect 110788 40122 110840 40128
rect 110892 40118 110920 41074
rect 112914 40828 113222 40837
rect 112914 40826 112920 40828
rect 112976 40826 113000 40828
rect 113056 40826 113080 40828
rect 113136 40826 113160 40828
rect 113216 40826 113222 40828
rect 112976 40774 112978 40826
rect 113158 40774 113160 40826
rect 112914 40772 112920 40774
rect 112976 40772 113000 40774
rect 113056 40772 113080 40774
rect 113136 40772 113160 40774
rect 113216 40772 113222 40774
rect 112914 40763 113222 40772
rect 113456 40520 113508 40526
rect 113456 40462 113508 40468
rect 110880 40112 110932 40118
rect 110880 40054 110932 40060
rect 110696 39636 110748 39642
rect 110696 39578 110748 39584
rect 110892 38554 110920 40054
rect 111340 40044 111392 40050
rect 111340 39986 111392 39992
rect 111156 39840 111208 39846
rect 111156 39782 111208 39788
rect 110972 38752 111024 38758
rect 110972 38694 111024 38700
rect 110880 38548 110932 38554
rect 110880 38490 110932 38496
rect 110524 37964 110644 37992
rect 110524 37754 110552 37964
rect 110616 37874 110736 37890
rect 110604 37868 110736 37874
rect 110656 37862 110736 37868
rect 110604 37810 110656 37816
rect 110524 37726 110644 37754
rect 110512 37664 110564 37670
rect 110512 37606 110564 37612
rect 110420 36916 110472 36922
rect 110420 36858 110472 36864
rect 110420 35692 110472 35698
rect 110420 35634 110472 35640
rect 110328 34536 110380 34542
rect 110328 34478 110380 34484
rect 110144 34400 110196 34406
rect 110144 34342 110196 34348
rect 110052 34128 110104 34134
rect 109972 34076 110052 34082
rect 109972 34070 110104 34076
rect 109972 34054 110092 34070
rect 109868 33992 109920 33998
rect 109868 33934 109920 33940
rect 109684 33652 109736 33658
rect 109684 33594 109736 33600
rect 109592 33380 109644 33386
rect 109592 33322 109644 33328
rect 109696 33114 109724 33594
rect 109776 33516 109828 33522
rect 109776 33458 109828 33464
rect 109684 33108 109736 33114
rect 109684 33050 109736 33056
rect 109788 32842 109816 33458
rect 109776 32836 109828 32842
rect 109776 32778 109828 32784
rect 109460 32716 109540 32722
rect 109408 32710 109540 32716
rect 109868 32768 109920 32774
rect 109868 32710 109920 32716
rect 109420 32694 109540 32710
rect 109512 32434 109540 32694
rect 108948 32428 109000 32434
rect 108948 32370 109000 32376
rect 109500 32428 109552 32434
rect 109500 32370 109552 32376
rect 109880 32366 109908 32710
rect 109868 32360 109920 32366
rect 109868 32302 109920 32308
rect 109408 32224 109460 32230
rect 109408 32166 109460 32172
rect 108764 31884 108816 31890
rect 108764 31826 108816 31832
rect 108304 31816 108356 31822
rect 108304 31758 108356 31764
rect 108488 31816 108540 31822
rect 108488 31758 108540 31764
rect 108856 31816 108908 31822
rect 108856 31758 108908 31764
rect 108316 31210 108344 31758
rect 108868 31414 108896 31758
rect 109420 31754 109448 32166
rect 109972 31890 110000 34054
rect 110052 33040 110104 33046
rect 110052 32982 110104 32988
rect 109960 31884 110012 31890
rect 109960 31826 110012 31832
rect 110064 31770 110092 32982
rect 110156 32570 110184 34342
rect 110236 33992 110288 33998
rect 110236 33934 110288 33940
rect 110248 33114 110276 33934
rect 110236 33108 110288 33114
rect 110236 33050 110288 33056
rect 110144 32564 110196 32570
rect 110144 32506 110196 32512
rect 110340 31958 110368 34478
rect 110432 33998 110460 35634
rect 110524 34474 110552 37606
rect 110616 35698 110644 37726
rect 110708 36582 110736 37862
rect 110788 37800 110840 37806
rect 110788 37742 110840 37748
rect 110800 37466 110828 37742
rect 110788 37460 110840 37466
rect 110788 37402 110840 37408
rect 110788 36712 110840 36718
rect 110788 36654 110840 36660
rect 110696 36576 110748 36582
rect 110696 36518 110748 36524
rect 110604 35692 110656 35698
rect 110604 35634 110656 35640
rect 110616 35086 110644 35634
rect 110604 35080 110656 35086
rect 110604 35022 110656 35028
rect 110604 34944 110656 34950
rect 110604 34886 110656 34892
rect 110616 34610 110644 34886
rect 110708 34678 110736 36518
rect 110800 36378 110828 36654
rect 110880 36576 110932 36582
rect 110880 36518 110932 36524
rect 110788 36372 110840 36378
rect 110788 36314 110840 36320
rect 110892 35222 110920 36518
rect 110984 36394 111012 38694
rect 111064 37732 111116 37738
rect 111064 37674 111116 37680
rect 111076 36854 111104 37674
rect 111064 36848 111116 36854
rect 111064 36790 111116 36796
rect 111168 36718 111196 39782
rect 111352 38962 111380 39986
rect 112914 39740 113222 39749
rect 112914 39738 112920 39740
rect 112976 39738 113000 39740
rect 113056 39738 113080 39740
rect 113136 39738 113160 39740
rect 113216 39738 113222 39740
rect 112976 39686 112978 39738
rect 113158 39686 113160 39738
rect 112914 39684 112920 39686
rect 112976 39684 113000 39686
rect 113056 39684 113080 39686
rect 113136 39684 113160 39686
rect 113216 39684 113222 39686
rect 112914 39675 113222 39684
rect 111340 38956 111392 38962
rect 111340 38898 111392 38904
rect 111248 37664 111300 37670
rect 111248 37606 111300 37612
rect 111260 37398 111288 37606
rect 111248 37392 111300 37398
rect 111248 37334 111300 37340
rect 111156 36712 111208 36718
rect 111156 36654 111208 36660
rect 110984 36366 111104 36394
rect 110972 36236 111024 36242
rect 110972 36178 111024 36184
rect 110984 35630 111012 36178
rect 110972 35624 111024 35630
rect 110972 35566 111024 35572
rect 110880 35216 110932 35222
rect 110880 35158 110932 35164
rect 111076 34950 111104 36366
rect 111248 35148 111300 35154
rect 111248 35090 111300 35096
rect 111064 34944 111116 34950
rect 111064 34886 111116 34892
rect 111076 34678 111104 34886
rect 111260 34746 111288 35090
rect 111248 34740 111300 34746
rect 111248 34682 111300 34688
rect 111352 34678 111380 38898
rect 112914 38652 113222 38661
rect 112914 38650 112920 38652
rect 112976 38650 113000 38652
rect 113056 38650 113080 38652
rect 113136 38650 113160 38652
rect 113216 38650 113222 38652
rect 112976 38598 112978 38650
rect 113158 38598 113160 38650
rect 112914 38596 112920 38598
rect 112976 38596 113000 38598
rect 113056 38596 113080 38598
rect 113136 38596 113160 38598
rect 113216 38596 113222 38598
rect 112914 38587 113222 38596
rect 111892 38344 111944 38350
rect 111892 38286 111944 38292
rect 112352 38344 112404 38350
rect 112352 38286 112404 38292
rect 111904 37806 111932 38286
rect 112364 37806 112392 38286
rect 113468 37874 113496 40462
rect 113650 40284 113958 40293
rect 113650 40282 113656 40284
rect 113712 40282 113736 40284
rect 113792 40282 113816 40284
rect 113872 40282 113896 40284
rect 113952 40282 113958 40284
rect 113712 40230 113714 40282
rect 113894 40230 113896 40282
rect 113650 40228 113656 40230
rect 113712 40228 113736 40230
rect 113792 40228 113816 40230
rect 113872 40228 113896 40230
rect 113952 40228 113958 40230
rect 113650 40219 113958 40228
rect 113650 39196 113958 39205
rect 113650 39194 113656 39196
rect 113712 39194 113736 39196
rect 113792 39194 113816 39196
rect 113872 39194 113896 39196
rect 113952 39194 113958 39196
rect 113712 39142 113714 39194
rect 113894 39142 113896 39194
rect 113650 39140 113656 39142
rect 113712 39140 113736 39142
rect 113792 39140 113816 39142
rect 113872 39140 113896 39142
rect 113952 39140 113958 39142
rect 113650 39131 113958 39140
rect 113650 38108 113958 38117
rect 113650 38106 113656 38108
rect 113712 38106 113736 38108
rect 113792 38106 113816 38108
rect 113872 38106 113896 38108
rect 113952 38106 113958 38108
rect 113712 38054 113714 38106
rect 113894 38054 113896 38106
rect 113650 38052 113656 38054
rect 113712 38052 113736 38054
rect 113792 38052 113816 38054
rect 113872 38052 113896 38054
rect 113952 38052 113958 38054
rect 113650 38043 113958 38052
rect 112812 37868 112864 37874
rect 112812 37810 112864 37816
rect 113456 37868 113508 37874
rect 113456 37810 113508 37816
rect 114560 37868 114612 37874
rect 114560 37810 114612 37816
rect 111892 37800 111944 37806
rect 111892 37742 111944 37748
rect 112352 37800 112404 37806
rect 112404 37748 112576 37754
rect 112352 37742 112576 37748
rect 112364 37726 112576 37742
rect 112444 37664 112496 37670
rect 112444 37606 112496 37612
rect 111708 37188 111760 37194
rect 111708 37130 111760 37136
rect 111720 35766 111748 37130
rect 112456 37126 112484 37606
rect 112548 37126 112576 37726
rect 112824 37398 112852 37810
rect 112914 37564 113222 37573
rect 112914 37562 112920 37564
rect 112976 37562 113000 37564
rect 113056 37562 113080 37564
rect 113136 37562 113160 37564
rect 113216 37562 113222 37564
rect 112976 37510 112978 37562
rect 113158 37510 113160 37562
rect 112914 37508 112920 37510
rect 112976 37508 113000 37510
rect 113056 37508 113080 37510
rect 113136 37508 113160 37510
rect 113216 37508 113222 37510
rect 112914 37499 113222 37508
rect 113468 37398 113496 37810
rect 113824 37800 113876 37806
rect 113824 37742 113876 37748
rect 113548 37460 113600 37466
rect 113548 37402 113600 37408
rect 112812 37392 112864 37398
rect 112812 37334 112864 37340
rect 113456 37392 113508 37398
rect 113456 37334 113508 37340
rect 113180 37256 113232 37262
rect 113180 37198 113232 37204
rect 112444 37120 112496 37126
rect 112444 37062 112496 37068
rect 112536 37120 112588 37126
rect 112536 37062 112588 37068
rect 112456 36922 112484 37062
rect 112444 36916 112496 36922
rect 112444 36858 112496 36864
rect 111892 36780 111944 36786
rect 111892 36722 111944 36728
rect 111904 35834 111932 36722
rect 112168 36576 112220 36582
rect 112168 36518 112220 36524
rect 112180 36106 112208 36518
rect 112548 36378 112576 37062
rect 112812 36848 112864 36854
rect 112812 36790 112864 36796
rect 112536 36372 112588 36378
rect 112536 36314 112588 36320
rect 112352 36304 112404 36310
rect 112352 36246 112404 36252
rect 112364 36174 112392 36246
rect 112824 36174 112852 36790
rect 113192 36786 113220 37198
rect 113454 36816 113510 36825
rect 113180 36780 113232 36786
rect 113180 36722 113232 36728
rect 113364 36780 113416 36786
rect 113454 36751 113510 36760
rect 113364 36722 113416 36728
rect 113192 36666 113220 36722
rect 113192 36638 113312 36666
rect 113376 36650 113404 36722
rect 112914 36476 113222 36485
rect 112914 36474 112920 36476
rect 112976 36474 113000 36476
rect 113056 36474 113080 36476
rect 113136 36474 113160 36476
rect 113216 36474 113222 36476
rect 112976 36422 112978 36474
rect 113158 36422 113160 36474
rect 112914 36420 112920 36422
rect 112976 36420 113000 36422
rect 113056 36420 113080 36422
rect 113136 36420 113160 36422
rect 113216 36420 113222 36422
rect 112914 36411 113222 36420
rect 113284 36174 113312 36638
rect 113364 36644 113416 36650
rect 113364 36586 113416 36592
rect 113376 36378 113404 36586
rect 113364 36372 113416 36378
rect 113364 36314 113416 36320
rect 112352 36168 112404 36174
rect 112352 36110 112404 36116
rect 112444 36168 112496 36174
rect 112444 36110 112496 36116
rect 112536 36168 112588 36174
rect 112536 36110 112588 36116
rect 112812 36168 112864 36174
rect 112812 36110 112864 36116
rect 113088 36168 113140 36174
rect 113088 36110 113140 36116
rect 113272 36168 113324 36174
rect 113272 36110 113324 36116
rect 112076 36100 112128 36106
rect 112076 36042 112128 36048
rect 112168 36100 112220 36106
rect 112168 36042 112220 36048
rect 111892 35828 111944 35834
rect 111892 35770 111944 35776
rect 111708 35760 111760 35766
rect 111708 35702 111760 35708
rect 111616 35624 111668 35630
rect 111616 35566 111668 35572
rect 111628 35290 111656 35566
rect 111616 35284 111668 35290
rect 111616 35226 111668 35232
rect 110696 34672 110748 34678
rect 110696 34614 110748 34620
rect 111064 34672 111116 34678
rect 111064 34614 111116 34620
rect 111340 34672 111392 34678
rect 111340 34614 111392 34620
rect 111720 34610 111748 35702
rect 112088 35222 112116 36042
rect 112456 35290 112484 36110
rect 112548 35698 112576 36110
rect 112824 35698 112852 36110
rect 113100 35698 113128 36110
rect 113272 36032 113324 36038
rect 113272 35974 113324 35980
rect 112536 35692 112588 35698
rect 112536 35634 112588 35640
rect 112812 35692 112864 35698
rect 112812 35634 112864 35640
rect 113088 35692 113140 35698
rect 113088 35634 113140 35640
rect 112536 35556 112588 35562
rect 112536 35498 112588 35504
rect 112548 35290 112576 35498
rect 112444 35284 112496 35290
rect 112444 35226 112496 35232
rect 112536 35284 112588 35290
rect 112536 35226 112588 35232
rect 112076 35216 112128 35222
rect 112076 35158 112128 35164
rect 111984 35012 112036 35018
rect 111984 34954 112036 34960
rect 111996 34728 112024 34954
rect 112076 34740 112128 34746
rect 111996 34700 112076 34728
rect 110604 34604 110656 34610
rect 110604 34546 110656 34552
rect 111708 34604 111760 34610
rect 111708 34546 111760 34552
rect 110512 34468 110564 34474
rect 110512 34410 110564 34416
rect 110524 34202 110552 34410
rect 110788 34400 110840 34406
rect 110788 34342 110840 34348
rect 110972 34400 111024 34406
rect 110972 34342 111024 34348
rect 111616 34400 111668 34406
rect 111616 34342 111668 34348
rect 110512 34196 110564 34202
rect 110512 34138 110564 34144
rect 110800 34066 110828 34342
rect 110984 34134 111012 34342
rect 110972 34128 111024 34134
rect 110972 34070 111024 34076
rect 110788 34060 110840 34066
rect 110788 34002 110840 34008
rect 110420 33992 110472 33998
rect 110420 33934 110472 33940
rect 111340 33992 111392 33998
rect 111628 33946 111656 34342
rect 111720 34066 111748 34546
rect 111892 34468 111944 34474
rect 111892 34410 111944 34416
rect 111708 34060 111760 34066
rect 111708 34002 111760 34008
rect 111340 33934 111392 33940
rect 110972 33856 111024 33862
rect 110972 33798 111024 33804
rect 110604 33448 110656 33454
rect 110604 33390 110656 33396
rect 110616 31958 110644 33390
rect 110984 32978 111012 33798
rect 111352 33522 111380 33934
rect 111444 33930 111748 33946
rect 111432 33924 111748 33930
rect 111484 33918 111748 33924
rect 111432 33866 111484 33872
rect 111444 33522 111472 33866
rect 111720 33862 111748 33918
rect 111616 33856 111668 33862
rect 111616 33798 111668 33804
rect 111708 33856 111760 33862
rect 111708 33798 111760 33804
rect 111800 33856 111852 33862
rect 111800 33798 111852 33804
rect 111340 33516 111392 33522
rect 111340 33458 111392 33464
rect 111432 33516 111484 33522
rect 111432 33458 111484 33464
rect 111628 33454 111656 33798
rect 111812 33522 111840 33798
rect 111800 33516 111852 33522
rect 111800 33458 111852 33464
rect 111616 33448 111668 33454
rect 111616 33390 111668 33396
rect 111628 32978 111656 33390
rect 110972 32972 111024 32978
rect 110972 32914 111024 32920
rect 111616 32972 111668 32978
rect 111616 32914 111668 32920
rect 111812 32910 111840 33458
rect 111800 32904 111852 32910
rect 111800 32846 111852 32852
rect 110972 32428 111024 32434
rect 110972 32370 111024 32376
rect 111432 32428 111484 32434
rect 111432 32370 111484 32376
rect 110880 32224 110932 32230
rect 110880 32166 110932 32172
rect 110328 31952 110380 31958
rect 110328 31894 110380 31900
rect 110604 31952 110656 31958
rect 110604 31894 110656 31900
rect 109420 31726 109540 31754
rect 108856 31408 108908 31414
rect 108856 31350 108908 31356
rect 108304 31204 108356 31210
rect 108304 31146 108356 31152
rect 107106 23624 107162 23633
rect 107106 23559 107162 23568
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9692 17283 9720 17614
rect 9678 17274 9734 17283
rect 9678 17209 9734 17218
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9692 15651 9720 15914
rect 9678 15642 9734 15651
rect 9678 15577 9734 15586
rect 106462 11928 106518 11937
rect 106462 11863 106518 11872
rect 93400 10056 93452 10062
rect 93400 9998 93452 10004
rect 92848 9988 92900 9994
rect 92848 9930 92900 9936
rect 15842 9888 15898 9897
rect 15842 9823 15898 9832
rect 92754 9888 92810 9897
rect 92860 9874 92888 9930
rect 92810 9846 92888 9874
rect 93032 9920 93084 9926
rect 93412 9897 93440 9998
rect 106476 9926 106504 11863
rect 108316 9994 108344 31146
rect 108764 31136 108816 31142
rect 108764 31078 108816 31084
rect 108776 10033 108804 31078
rect 109224 30728 109276 30734
rect 109224 30670 109276 30676
rect 109236 30394 109264 30670
rect 109224 30388 109276 30394
rect 109224 30330 109276 30336
rect 109512 10062 109540 31726
rect 109972 31742 110092 31770
rect 110420 31816 110472 31822
rect 110420 31758 110472 31764
rect 109592 31340 109644 31346
rect 109592 31282 109644 31288
rect 109604 30938 109632 31282
rect 109592 30932 109644 30938
rect 109592 30874 109644 30880
rect 109684 30728 109736 30734
rect 109684 30670 109736 30676
rect 109592 30320 109644 30326
rect 109592 30262 109644 30268
rect 109604 29646 109632 30262
rect 109696 29850 109724 30670
rect 109972 30376 110000 31742
rect 110052 31408 110104 31414
rect 110052 31350 110104 31356
rect 110064 30870 110092 31350
rect 110052 30864 110104 30870
rect 110052 30806 110104 30812
rect 110328 30728 110380 30734
rect 110328 30670 110380 30676
rect 109788 30348 110000 30376
rect 109788 30258 109816 30348
rect 109776 30252 109828 30258
rect 109776 30194 109828 30200
rect 109868 30252 109920 30258
rect 109868 30194 109920 30200
rect 109684 29844 109736 29850
rect 109684 29786 109736 29792
rect 109776 29844 109828 29850
rect 109776 29786 109828 29792
rect 109788 29646 109816 29786
rect 109880 29714 109908 30194
rect 109868 29708 109920 29714
rect 109868 29650 109920 29656
rect 109972 29696 110000 30348
rect 110144 30252 110196 30258
rect 110144 30194 110196 30200
rect 110156 29850 110184 30194
rect 110144 29844 110196 29850
rect 110144 29786 110196 29792
rect 110052 29708 110104 29714
rect 109972 29668 110052 29696
rect 109592 29640 109644 29646
rect 109592 29582 109644 29588
rect 109776 29640 109828 29646
rect 109776 29582 109828 29588
rect 109604 29306 109632 29582
rect 109592 29300 109644 29306
rect 109592 29242 109644 29248
rect 109788 29238 109816 29582
rect 109880 29306 109908 29650
rect 109868 29300 109920 29306
rect 109868 29242 109920 29248
rect 109776 29232 109828 29238
rect 109776 29174 109828 29180
rect 109684 29096 109736 29102
rect 109736 29044 109816 29050
rect 109684 29038 109816 29044
rect 109696 29022 109816 29038
rect 109788 28626 109816 29022
rect 109972 28642 110000 29668
rect 110052 29650 110104 29656
rect 110144 29640 110196 29646
rect 110196 29588 110276 29594
rect 110144 29582 110276 29588
rect 110156 29566 110276 29582
rect 110052 29504 110104 29510
rect 110052 29446 110104 29452
rect 110064 28762 110092 29446
rect 110144 29300 110196 29306
rect 110144 29242 110196 29248
rect 110156 29170 110184 29242
rect 110144 29164 110196 29170
rect 110144 29106 110196 29112
rect 110052 28756 110104 28762
rect 110052 28698 110104 28704
rect 109776 28620 109828 28626
rect 109972 28614 110092 28642
rect 110156 28626 110184 29106
rect 109776 28562 109828 28568
rect 109788 28082 109816 28562
rect 109868 28552 109920 28558
rect 109868 28494 109920 28500
rect 109776 28076 109828 28082
rect 109776 28018 109828 28024
rect 109880 27538 109908 28494
rect 109960 28076 110012 28082
rect 109960 28018 110012 28024
rect 109972 27674 110000 28018
rect 109960 27668 110012 27674
rect 109960 27610 110012 27616
rect 110064 27606 110092 28614
rect 110144 28620 110196 28626
rect 110144 28562 110196 28568
rect 110248 28558 110276 29566
rect 110340 29306 110368 30670
rect 110432 30326 110460 31758
rect 110512 31272 110564 31278
rect 110512 31214 110564 31220
rect 110524 30938 110552 31214
rect 110616 31210 110644 31894
rect 110892 31890 110920 32166
rect 110880 31884 110932 31890
rect 110880 31826 110932 31832
rect 110984 31482 111012 32370
rect 111340 32360 111392 32366
rect 111340 32302 111392 32308
rect 111352 31634 111380 32302
rect 111444 31754 111472 32370
rect 111708 31952 111760 31958
rect 111708 31894 111760 31900
rect 111444 31726 111564 31754
rect 111536 31686 111564 31726
rect 111432 31680 111484 31686
rect 111352 31628 111432 31634
rect 111352 31622 111484 31628
rect 111524 31680 111576 31686
rect 111524 31622 111576 31628
rect 111352 31606 111472 31622
rect 110972 31476 111024 31482
rect 110972 31418 111024 31424
rect 111338 31240 111394 31249
rect 110604 31204 110656 31210
rect 111338 31175 111394 31184
rect 110604 31146 110656 31152
rect 111352 31142 111380 31175
rect 111340 31136 111392 31142
rect 111340 31078 111392 31084
rect 111444 30938 111472 31606
rect 110512 30932 110564 30938
rect 110512 30874 110564 30880
rect 111432 30932 111484 30938
rect 111432 30874 111484 30880
rect 110880 30796 110932 30802
rect 110880 30738 110932 30744
rect 110512 30728 110564 30734
rect 110512 30670 110564 30676
rect 110420 30320 110472 30326
rect 110420 30262 110472 30268
rect 110432 29782 110460 30262
rect 110420 29776 110472 29782
rect 110420 29718 110472 29724
rect 110524 29322 110552 30670
rect 110892 30394 110920 30738
rect 111340 30728 111392 30734
rect 111340 30670 111392 30676
rect 110880 30388 110932 30394
rect 110880 30330 110932 30336
rect 110892 30258 110920 30330
rect 110604 30252 110656 30258
rect 110604 30194 110656 30200
rect 110880 30252 110932 30258
rect 110880 30194 110932 30200
rect 111248 30252 111300 30258
rect 111248 30194 111300 30200
rect 110616 29850 110644 30194
rect 111156 30048 111208 30054
rect 111156 29990 111208 29996
rect 111168 29850 111196 29990
rect 110604 29844 110656 29850
rect 110604 29786 110656 29792
rect 111156 29844 111208 29850
rect 111156 29786 111208 29792
rect 111260 29782 111288 30194
rect 110972 29776 111024 29782
rect 110972 29718 111024 29724
rect 111248 29776 111300 29782
rect 111248 29718 111300 29724
rect 110984 29646 111012 29718
rect 110788 29640 110840 29646
rect 110788 29582 110840 29588
rect 110972 29640 111024 29646
rect 110972 29582 111024 29588
rect 111064 29640 111116 29646
rect 111064 29582 111116 29588
rect 110328 29300 110380 29306
rect 110328 29242 110380 29248
rect 110432 29294 110552 29322
rect 110800 29306 110828 29582
rect 110788 29300 110840 29306
rect 110432 29102 110460 29294
rect 110788 29242 110840 29248
rect 110604 29164 110656 29170
rect 110604 29106 110656 29112
rect 110420 29096 110472 29102
rect 110420 29038 110472 29044
rect 110432 28966 110460 29038
rect 110420 28960 110472 28966
rect 110420 28902 110472 28908
rect 110236 28552 110288 28558
rect 110236 28494 110288 28500
rect 110248 28218 110276 28494
rect 110432 28490 110460 28902
rect 110616 28694 110644 29106
rect 111076 29034 111104 29582
rect 111352 29170 111380 30670
rect 111536 30394 111564 31622
rect 111616 31136 111668 31142
rect 111616 31078 111668 31084
rect 111628 30734 111656 31078
rect 111720 30938 111748 31894
rect 111904 31890 111932 34410
rect 111996 33522 112024 34700
rect 112076 34682 112128 34688
rect 111984 33516 112036 33522
rect 111984 33458 112036 33464
rect 111996 33046 112024 33458
rect 111984 33040 112036 33046
rect 111984 32982 112036 32988
rect 112548 32842 112576 35226
rect 112824 35018 112852 35634
rect 112914 35388 113222 35397
rect 112914 35386 112920 35388
rect 112976 35386 113000 35388
rect 113056 35386 113080 35388
rect 113136 35386 113160 35388
rect 113216 35386 113222 35388
rect 112976 35334 112978 35386
rect 113158 35334 113160 35386
rect 112914 35332 112920 35334
rect 112976 35332 113000 35334
rect 113056 35332 113080 35334
rect 113136 35332 113160 35334
rect 113216 35332 113222 35334
rect 112914 35323 113222 35332
rect 112996 35284 113048 35290
rect 112996 35226 113048 35232
rect 112904 35080 112956 35086
rect 112904 35022 112956 35028
rect 112812 35012 112864 35018
rect 112812 34954 112864 34960
rect 112916 34388 112944 35022
rect 113008 34950 113036 35226
rect 113284 35222 113312 35974
rect 113364 35828 113416 35834
rect 113364 35770 113416 35776
rect 113272 35216 113324 35222
rect 113272 35158 113324 35164
rect 113376 35086 113404 35770
rect 113468 35630 113496 36751
rect 113560 36530 113588 37402
rect 113836 37330 113864 37742
rect 114100 37664 114152 37670
rect 114100 37606 114152 37612
rect 114468 37664 114520 37670
rect 114468 37606 114520 37612
rect 113824 37324 113876 37330
rect 113824 37266 113876 37272
rect 114008 37256 114060 37262
rect 114008 37198 114060 37204
rect 113650 37020 113958 37029
rect 113650 37018 113656 37020
rect 113712 37018 113736 37020
rect 113792 37018 113816 37020
rect 113872 37018 113896 37020
rect 113952 37018 113958 37020
rect 113712 36966 113714 37018
rect 113894 36966 113896 37018
rect 113650 36964 113656 36966
rect 113712 36964 113736 36966
rect 113792 36964 113816 36966
rect 113872 36964 113896 36966
rect 113952 36964 113958 36966
rect 113650 36955 113958 36964
rect 114020 36825 114048 37198
rect 114112 36854 114140 37606
rect 114284 37256 114336 37262
rect 114284 37198 114336 37204
rect 114376 37256 114428 37262
rect 114376 37198 114428 37204
rect 114192 37188 114244 37194
rect 114192 37130 114244 37136
rect 114100 36848 114152 36854
rect 114006 36816 114062 36825
rect 113916 36780 113968 36786
rect 114100 36790 114152 36796
rect 114006 36751 114008 36760
rect 113916 36722 113968 36728
rect 114060 36751 114062 36760
rect 114008 36722 114060 36728
rect 113928 36582 113956 36722
rect 113916 36576 113968 36582
rect 113560 36502 113864 36530
rect 113916 36518 113968 36524
rect 113548 36304 113600 36310
rect 113548 36246 113600 36252
rect 113560 35698 113588 36246
rect 113836 36174 113864 36502
rect 114100 36236 114152 36242
rect 114100 36178 114152 36184
rect 113824 36168 113876 36174
rect 113824 36110 113876 36116
rect 114008 36168 114060 36174
rect 114008 36110 114060 36116
rect 113836 36038 113864 36110
rect 113824 36032 113876 36038
rect 113824 35974 113876 35980
rect 113650 35932 113958 35941
rect 113650 35930 113656 35932
rect 113712 35930 113736 35932
rect 113792 35930 113816 35932
rect 113872 35930 113896 35932
rect 113952 35930 113958 35932
rect 113712 35878 113714 35930
rect 113894 35878 113896 35930
rect 113650 35876 113656 35878
rect 113712 35876 113736 35878
rect 113792 35876 113816 35878
rect 113872 35876 113896 35878
rect 113952 35876 113958 35878
rect 113650 35867 113958 35876
rect 114020 35834 114048 36110
rect 114008 35828 114060 35834
rect 114008 35770 114060 35776
rect 113548 35692 113600 35698
rect 113548 35634 113600 35640
rect 113456 35624 113508 35630
rect 113456 35566 113508 35572
rect 114112 35290 114140 36178
rect 114204 35630 114232 37130
rect 114296 36786 114324 37198
rect 114388 36786 114416 37198
rect 114480 36854 114508 37606
rect 114572 37194 114600 37810
rect 116400 37324 116452 37330
rect 116400 37266 116452 37272
rect 115020 37256 115072 37262
rect 115020 37198 115072 37204
rect 116308 37256 116360 37262
rect 116308 37198 116360 37204
rect 114560 37188 114612 37194
rect 114560 37130 114612 37136
rect 114836 37188 114888 37194
rect 114836 37130 114888 37136
rect 114848 36922 114876 37130
rect 114652 36916 114704 36922
rect 114652 36858 114704 36864
rect 114836 36916 114888 36922
rect 114836 36858 114888 36864
rect 114468 36848 114520 36854
rect 114468 36790 114520 36796
rect 114664 36786 114692 36858
rect 115032 36786 115060 37198
rect 116216 37120 116268 37126
rect 116216 37062 116268 37068
rect 116228 36922 116256 37062
rect 116124 36916 116176 36922
rect 116124 36858 116176 36864
rect 116216 36916 116268 36922
rect 116216 36858 116268 36864
rect 115112 36848 115164 36854
rect 115110 36816 115112 36825
rect 115572 36848 115624 36854
rect 115164 36816 115166 36825
rect 114284 36780 114336 36786
rect 114284 36722 114336 36728
rect 114376 36780 114428 36786
rect 114376 36722 114428 36728
rect 114652 36780 114704 36786
rect 114652 36722 114704 36728
rect 114928 36780 114980 36786
rect 114928 36722 114980 36728
rect 115020 36780 115072 36786
rect 115572 36790 115624 36796
rect 115110 36751 115166 36760
rect 115020 36722 115072 36728
rect 114296 35766 114324 36722
rect 114388 36310 114416 36722
rect 114940 36310 114968 36722
rect 115032 36378 115060 36722
rect 115204 36576 115256 36582
rect 115204 36518 115256 36524
rect 115020 36372 115072 36378
rect 115020 36314 115072 36320
rect 114376 36304 114428 36310
rect 114376 36246 114428 36252
rect 114928 36304 114980 36310
rect 114928 36246 114980 36252
rect 115216 36242 115244 36518
rect 115584 36378 115612 36790
rect 116136 36786 116164 36858
rect 115848 36780 115900 36786
rect 115848 36722 115900 36728
rect 116124 36780 116176 36786
rect 116124 36722 116176 36728
rect 115572 36372 115624 36378
rect 115572 36314 115624 36320
rect 115388 36304 115440 36310
rect 115388 36246 115440 36252
rect 115204 36236 115256 36242
rect 115204 36178 115256 36184
rect 114468 36100 114520 36106
rect 115204 36100 115256 36106
rect 114520 36060 114600 36088
rect 114468 36042 114520 36048
rect 114284 35760 114336 35766
rect 114284 35702 114336 35708
rect 114376 35692 114428 35698
rect 114376 35634 114428 35640
rect 114192 35624 114244 35630
rect 114192 35566 114244 35572
rect 114100 35284 114152 35290
rect 114100 35226 114152 35232
rect 113640 35216 113692 35222
rect 113640 35158 113692 35164
rect 113456 35148 113508 35154
rect 113456 35090 113508 35096
rect 113364 35080 113416 35086
rect 113364 35022 113416 35028
rect 112996 34944 113048 34950
rect 112996 34886 113048 34892
rect 112824 34360 112944 34388
rect 112824 34134 112852 34360
rect 112914 34300 113222 34309
rect 112914 34298 112920 34300
rect 112976 34298 113000 34300
rect 113056 34298 113080 34300
rect 113136 34298 113160 34300
rect 113216 34298 113222 34300
rect 112976 34246 112978 34298
rect 113158 34246 113160 34298
rect 112914 34244 112920 34246
rect 112976 34244 113000 34246
rect 113056 34244 113080 34246
rect 113136 34244 113160 34246
rect 113216 34244 113222 34246
rect 112914 34235 113222 34244
rect 113468 34202 113496 35090
rect 113652 35086 113680 35158
rect 114192 35148 114244 35154
rect 114192 35090 114244 35096
rect 113640 35080 113692 35086
rect 113640 35022 113692 35028
rect 114008 34944 114060 34950
rect 114008 34886 114060 34892
rect 114100 34944 114152 34950
rect 114100 34886 114152 34892
rect 113650 34844 113958 34853
rect 113650 34842 113656 34844
rect 113712 34842 113736 34844
rect 113792 34842 113816 34844
rect 113872 34842 113896 34844
rect 113952 34842 113958 34844
rect 113712 34790 113714 34842
rect 113894 34790 113896 34842
rect 113650 34788 113656 34790
rect 113712 34788 113736 34790
rect 113792 34788 113816 34790
rect 113872 34788 113896 34790
rect 113952 34788 113958 34790
rect 113650 34779 113958 34788
rect 113548 34536 113600 34542
rect 113548 34478 113600 34484
rect 113456 34196 113508 34202
rect 113456 34138 113508 34144
rect 112812 34128 112864 34134
rect 112812 34070 112864 34076
rect 112628 33516 112680 33522
rect 112628 33458 112680 33464
rect 112720 33516 112772 33522
rect 112720 33458 112772 33464
rect 112536 32836 112588 32842
rect 112536 32778 112588 32784
rect 112640 32570 112668 33458
rect 112732 32910 112760 33458
rect 112914 33212 113222 33221
rect 112914 33210 112920 33212
rect 112976 33210 113000 33212
rect 113056 33210 113080 33212
rect 113136 33210 113160 33212
rect 113216 33210 113222 33212
rect 112976 33158 112978 33210
rect 113158 33158 113160 33210
rect 112914 33156 112920 33158
rect 112976 33156 113000 33158
rect 113056 33156 113080 33158
rect 113136 33156 113160 33158
rect 113216 33156 113222 33158
rect 112914 33147 113222 33156
rect 112720 32904 112772 32910
rect 112720 32846 112772 32852
rect 112628 32564 112680 32570
rect 112628 32506 112680 32512
rect 112732 32434 112760 32846
rect 112996 32836 113048 32842
rect 112996 32778 113048 32784
rect 113008 32434 113036 32778
rect 113180 32768 113232 32774
rect 113180 32710 113232 32716
rect 112168 32428 112220 32434
rect 112168 32370 112220 32376
rect 112720 32428 112772 32434
rect 112720 32370 112772 32376
rect 112996 32428 113048 32434
rect 112996 32370 113048 32376
rect 112076 32360 112128 32366
rect 112076 32302 112128 32308
rect 111984 32224 112036 32230
rect 111984 32166 112036 32172
rect 111892 31884 111944 31890
rect 111892 31826 111944 31832
rect 111800 31816 111852 31822
rect 111800 31758 111852 31764
rect 111812 31414 111840 31758
rect 111904 31482 111932 31826
rect 111892 31476 111944 31482
rect 111892 31418 111944 31424
rect 111800 31408 111852 31414
rect 111800 31350 111852 31356
rect 111996 31346 112024 32166
rect 112088 32026 112116 32302
rect 112076 32020 112128 32026
rect 112076 31962 112128 31968
rect 112180 31482 112208 32370
rect 112444 32360 112496 32366
rect 112444 32302 112496 32308
rect 113192 32314 113220 32710
rect 112260 32224 112312 32230
rect 112260 32166 112312 32172
rect 112352 32224 112404 32230
rect 112352 32166 112404 32172
rect 112168 31476 112220 31482
rect 112168 31418 112220 31424
rect 112272 31346 112300 32166
rect 112364 31754 112392 32166
rect 112352 31748 112404 31754
rect 112352 31690 112404 31696
rect 111892 31340 111944 31346
rect 111892 31282 111944 31288
rect 111984 31340 112036 31346
rect 111984 31282 112036 31288
rect 112260 31340 112312 31346
rect 112260 31282 112312 31288
rect 111904 31249 111932 31282
rect 112364 31278 112392 31690
rect 112456 31482 112484 32302
rect 113192 32286 113312 32314
rect 112914 32124 113222 32133
rect 112914 32122 112920 32124
rect 112976 32122 113000 32124
rect 113056 32122 113080 32124
rect 113136 32122 113160 32124
rect 113216 32122 113222 32124
rect 112976 32070 112978 32122
rect 113158 32070 113160 32122
rect 112914 32068 112920 32070
rect 112976 32068 113000 32070
rect 113056 32068 113080 32070
rect 113136 32068 113160 32070
rect 113216 32068 113222 32070
rect 112914 32059 113222 32068
rect 113180 31952 113232 31958
rect 113180 31894 113232 31900
rect 112444 31476 112496 31482
rect 112444 31418 112496 31424
rect 112812 31340 112864 31346
rect 112812 31282 112864 31288
rect 112352 31272 112404 31278
rect 111890 31240 111946 31249
rect 112352 31214 112404 31220
rect 112536 31272 112588 31278
rect 112536 31214 112588 31220
rect 111890 31175 111946 31184
rect 111708 30932 111760 30938
rect 111708 30874 111760 30880
rect 112548 30841 112576 31214
rect 112534 30832 112590 30841
rect 111904 30802 112024 30818
rect 111892 30796 112024 30802
rect 111944 30790 112024 30796
rect 111892 30738 111944 30744
rect 111616 30728 111668 30734
rect 111616 30670 111668 30676
rect 111892 30660 111944 30666
rect 111892 30602 111944 30608
rect 111524 30388 111576 30394
rect 111524 30330 111576 30336
rect 111904 30190 111932 30602
rect 111996 30258 112024 30790
rect 112534 30767 112590 30776
rect 112076 30592 112128 30598
rect 112076 30534 112128 30540
rect 112088 30394 112116 30534
rect 112076 30388 112128 30394
rect 112076 30330 112128 30336
rect 112548 30326 112576 30767
rect 112536 30320 112588 30326
rect 112536 30262 112588 30268
rect 112824 30258 112852 31282
rect 113192 31124 113220 31894
rect 113284 31822 113312 32286
rect 113456 32292 113508 32298
rect 113456 32234 113508 32240
rect 113272 31816 113324 31822
rect 113272 31758 113324 31764
rect 113284 31414 113312 31758
rect 113468 31754 113496 32234
rect 113456 31748 113508 31754
rect 113456 31690 113508 31696
rect 113272 31408 113324 31414
rect 113272 31350 113324 31356
rect 113468 31346 113496 31690
rect 113456 31340 113508 31346
rect 113456 31282 113508 31288
rect 113364 31204 113416 31210
rect 113364 31146 113416 31152
rect 113192 31096 113312 31124
rect 112914 31036 113222 31045
rect 112914 31034 112920 31036
rect 112976 31034 113000 31036
rect 113056 31034 113080 31036
rect 113136 31034 113160 31036
rect 113216 31034 113222 31036
rect 112976 30982 112978 31034
rect 113158 30982 113160 31034
rect 112914 30980 112920 30982
rect 112976 30980 113000 30982
rect 113056 30980 113080 30982
rect 113136 30980 113160 30982
rect 113216 30980 113222 30982
rect 112914 30971 113222 30980
rect 113086 30832 113142 30841
rect 113284 30802 113312 31096
rect 113086 30767 113142 30776
rect 113272 30796 113324 30802
rect 113100 30734 113128 30767
rect 113272 30738 113324 30744
rect 113088 30728 113140 30734
rect 113088 30670 113140 30676
rect 113100 30598 113128 30670
rect 113376 30666 113404 31146
rect 113560 30818 113588 34478
rect 113732 34400 113784 34406
rect 113732 34342 113784 34348
rect 113744 33930 113772 34342
rect 114020 34202 114048 34886
rect 114112 34746 114140 34886
rect 114100 34740 114152 34746
rect 114100 34682 114152 34688
rect 114098 34640 114154 34649
rect 114098 34575 114100 34584
rect 114152 34575 114154 34584
rect 114100 34546 114152 34552
rect 114008 34196 114060 34202
rect 114008 34138 114060 34144
rect 113732 33924 113784 33930
rect 113732 33866 113784 33872
rect 113650 33756 113958 33765
rect 113650 33754 113656 33756
rect 113712 33754 113736 33756
rect 113792 33754 113816 33756
rect 113872 33754 113896 33756
rect 113952 33754 113958 33756
rect 113712 33702 113714 33754
rect 113894 33702 113896 33754
rect 113650 33700 113656 33702
rect 113712 33700 113736 33702
rect 113792 33700 113816 33702
rect 113872 33700 113896 33702
rect 113952 33700 113958 33702
rect 113650 33691 113958 33700
rect 114008 33448 114060 33454
rect 114008 33390 114060 33396
rect 113650 32668 113958 32677
rect 113650 32666 113656 32668
rect 113712 32666 113736 32668
rect 113792 32666 113816 32668
rect 113872 32666 113896 32668
rect 113952 32666 113958 32668
rect 113712 32614 113714 32666
rect 113894 32614 113896 32666
rect 113650 32612 113656 32614
rect 113712 32612 113736 32614
rect 113792 32612 113816 32614
rect 113872 32612 113896 32614
rect 113952 32612 113958 32614
rect 113650 32603 113958 32612
rect 114020 32552 114048 33390
rect 113928 32524 114048 32552
rect 113928 32230 113956 32524
rect 113916 32224 113968 32230
rect 113916 32166 113968 32172
rect 113928 31754 113956 32166
rect 114112 31958 114140 34546
rect 114204 34406 114232 35090
rect 114388 34950 114416 35634
rect 114468 35624 114520 35630
rect 114468 35566 114520 35572
rect 114480 35086 114508 35566
rect 114572 35222 114600 36060
rect 115204 36042 115256 36048
rect 114836 36032 114888 36038
rect 114836 35974 114888 35980
rect 114928 36032 114980 36038
rect 114928 35974 114980 35980
rect 114848 35834 114876 35974
rect 114836 35828 114888 35834
rect 114836 35770 114888 35776
rect 114560 35216 114612 35222
rect 114560 35158 114612 35164
rect 114652 35148 114704 35154
rect 114652 35090 114704 35096
rect 114468 35080 114520 35086
rect 114468 35022 114520 35028
rect 114376 34944 114428 34950
rect 114376 34886 114428 34892
rect 114480 34746 114508 35022
rect 114664 34950 114692 35090
rect 114652 34944 114704 34950
rect 114652 34886 114704 34892
rect 114468 34740 114520 34746
rect 114468 34682 114520 34688
rect 114940 34678 114968 35974
rect 115216 35698 115244 36042
rect 115296 36032 115348 36038
rect 115296 35974 115348 35980
rect 115308 35698 115336 35974
rect 115204 35692 115256 35698
rect 115124 35652 115204 35680
rect 115124 35290 115152 35652
rect 115204 35634 115256 35640
rect 115296 35692 115348 35698
rect 115296 35634 115348 35640
rect 115204 35488 115256 35494
rect 115204 35430 115256 35436
rect 115112 35284 115164 35290
rect 115112 35226 115164 35232
rect 115216 35086 115244 35430
rect 115204 35080 115256 35086
rect 115204 35022 115256 35028
rect 115296 35080 115348 35086
rect 115296 35022 115348 35028
rect 115308 34950 115336 35022
rect 115296 34944 115348 34950
rect 115296 34886 115348 34892
rect 114928 34672 114980 34678
rect 114928 34614 114980 34620
rect 114284 34604 114336 34610
rect 114284 34546 114336 34552
rect 115020 34604 115072 34610
rect 115020 34546 115072 34552
rect 114192 34400 114244 34406
rect 114192 34342 114244 34348
rect 114296 34202 114324 34546
rect 114560 34468 114612 34474
rect 114560 34410 114612 34416
rect 114284 34196 114336 34202
rect 114284 34138 114336 34144
rect 114192 33992 114244 33998
rect 114192 33934 114244 33940
rect 114204 32298 114232 33934
rect 114376 33856 114428 33862
rect 114376 33798 114428 33804
rect 114284 32768 114336 32774
rect 114284 32710 114336 32716
rect 114296 32434 114324 32710
rect 114284 32428 114336 32434
rect 114284 32370 114336 32376
rect 114192 32292 114244 32298
rect 114192 32234 114244 32240
rect 114100 31952 114152 31958
rect 114098 31920 114100 31929
rect 114152 31920 114154 31929
rect 114098 31855 114154 31864
rect 114008 31816 114060 31822
rect 114008 31758 114060 31764
rect 114100 31816 114152 31822
rect 114100 31758 114152 31764
rect 113916 31748 113968 31754
rect 113916 31690 113968 31696
rect 113650 31580 113958 31589
rect 113650 31578 113656 31580
rect 113712 31578 113736 31580
rect 113792 31578 113816 31580
rect 113872 31578 113896 31580
rect 113952 31578 113958 31580
rect 113712 31526 113714 31578
rect 113894 31526 113896 31578
rect 113650 31524 113656 31526
rect 113712 31524 113736 31526
rect 113792 31524 113816 31526
rect 113872 31524 113896 31526
rect 113952 31524 113958 31526
rect 113650 31515 113958 31524
rect 113824 31340 113876 31346
rect 114020 31328 114048 31758
rect 114112 31346 114140 31758
rect 114284 31748 114336 31754
rect 114284 31690 114336 31696
rect 114296 31498 114324 31690
rect 114388 31686 114416 33798
rect 114572 33522 114600 34410
rect 115032 34202 115060 34546
rect 115112 34536 115164 34542
rect 115112 34478 115164 34484
rect 115020 34196 115072 34202
rect 115020 34138 115072 34144
rect 114928 33992 114980 33998
rect 114926 33960 114928 33969
rect 114980 33960 114982 33969
rect 114926 33895 114982 33904
rect 114560 33516 114612 33522
rect 114560 33458 114612 33464
rect 114836 33516 114888 33522
rect 114836 33458 114888 33464
rect 114572 33114 114600 33458
rect 114560 33108 114612 33114
rect 114560 33050 114612 33056
rect 114468 32564 114520 32570
rect 114468 32506 114520 32512
rect 114480 31890 114508 32506
rect 114468 31884 114520 31890
rect 114468 31826 114520 31832
rect 114376 31680 114428 31686
rect 114376 31622 114428 31628
rect 114296 31470 114416 31498
rect 114480 31482 114508 31826
rect 113876 31300 114048 31328
rect 114100 31340 114152 31346
rect 113824 31282 113876 31288
rect 114100 31282 114152 31288
rect 114284 31340 114336 31346
rect 114284 31282 114336 31288
rect 113468 30790 113588 30818
rect 113364 30660 113416 30666
rect 113364 30602 113416 30608
rect 113088 30592 113140 30598
rect 113088 30534 113140 30540
rect 111984 30252 112036 30258
rect 111984 30194 112036 30200
rect 112076 30252 112128 30258
rect 112076 30194 112128 30200
rect 112260 30252 112312 30258
rect 112260 30194 112312 30200
rect 112812 30252 112864 30258
rect 112812 30194 112864 30200
rect 111892 30184 111944 30190
rect 111892 30126 111944 30132
rect 111996 29730 112024 30194
rect 111904 29702 112024 29730
rect 112088 29714 112116 30194
rect 112076 29708 112128 29714
rect 111904 29646 111932 29702
rect 112076 29650 112128 29656
rect 111708 29640 111760 29646
rect 111708 29582 111760 29588
rect 111892 29640 111944 29646
rect 111892 29582 111944 29588
rect 111340 29164 111392 29170
rect 111340 29106 111392 29112
rect 111064 29028 111116 29034
rect 111064 28970 111116 28976
rect 111720 28762 111748 29582
rect 111800 29028 111852 29034
rect 111800 28970 111852 28976
rect 111708 28756 111760 28762
rect 111708 28698 111760 28704
rect 110604 28688 110656 28694
rect 110604 28630 110656 28636
rect 110420 28484 110472 28490
rect 110420 28426 110472 28432
rect 110788 28484 110840 28490
rect 110788 28426 110840 28432
rect 110236 28212 110288 28218
rect 110236 28154 110288 28160
rect 110800 28014 110828 28426
rect 111812 28098 111840 28970
rect 111904 28642 111932 29582
rect 111984 29096 112036 29102
rect 111984 29038 112036 29044
rect 111996 28762 112024 29038
rect 111984 28756 112036 28762
rect 111984 28698 112036 28704
rect 111904 28614 112024 28642
rect 111720 28082 111840 28098
rect 111064 28076 111116 28082
rect 111064 28018 111116 28024
rect 111708 28076 111840 28082
rect 111760 28070 111840 28076
rect 111708 28018 111760 28024
rect 110788 28008 110840 28014
rect 110788 27950 110840 27956
rect 110052 27600 110104 27606
rect 110052 27542 110104 27548
rect 109868 27532 109920 27538
rect 109868 27474 109920 27480
rect 109880 26382 109908 27474
rect 110800 27130 110828 27950
rect 111076 27606 111104 28018
rect 111892 27872 111944 27878
rect 111892 27814 111944 27820
rect 111064 27600 111116 27606
rect 111064 27542 111116 27548
rect 111904 27538 111932 27814
rect 111248 27532 111300 27538
rect 111248 27474 111300 27480
rect 111892 27532 111944 27538
rect 111892 27474 111944 27480
rect 110972 27464 111024 27470
rect 110972 27406 111024 27412
rect 110788 27124 110840 27130
rect 110788 27066 110840 27072
rect 110984 26994 111012 27406
rect 111260 26994 111288 27474
rect 111340 27464 111392 27470
rect 111340 27406 111392 27412
rect 111352 26994 111380 27406
rect 111996 27334 112024 28614
rect 111984 27328 112036 27334
rect 111984 27270 112036 27276
rect 112088 26994 112116 29650
rect 112272 29578 112300 30194
rect 112260 29572 112312 29578
rect 112260 29514 112312 29520
rect 112824 29510 112852 30194
rect 112914 29948 113222 29957
rect 112914 29946 112920 29948
rect 112976 29946 113000 29948
rect 113056 29946 113080 29948
rect 113136 29946 113160 29948
rect 113216 29946 113222 29948
rect 112976 29894 112978 29946
rect 113158 29894 113160 29946
rect 112914 29892 112920 29894
rect 112976 29892 113000 29894
rect 113056 29892 113080 29894
rect 113136 29892 113160 29894
rect 113216 29892 113222 29894
rect 112914 29883 113222 29892
rect 112812 29504 112864 29510
rect 112812 29446 112864 29452
rect 113364 29300 113416 29306
rect 113364 29242 113416 29248
rect 112914 28860 113222 28869
rect 112914 28858 112920 28860
rect 112976 28858 113000 28860
rect 113056 28858 113080 28860
rect 113136 28858 113160 28860
rect 113216 28858 113222 28860
rect 112976 28806 112978 28858
rect 113158 28806 113160 28858
rect 112914 28804 112920 28806
rect 112976 28804 113000 28806
rect 113056 28804 113080 28806
rect 113136 28804 113160 28806
rect 113216 28804 113222 28806
rect 112914 28795 113222 28804
rect 112444 28756 112496 28762
rect 112444 28698 112496 28704
rect 112456 28558 112484 28698
rect 112260 28552 112312 28558
rect 112260 28494 112312 28500
rect 112444 28552 112496 28558
rect 112444 28494 112496 28500
rect 112272 28082 112300 28494
rect 112628 28416 112680 28422
rect 112628 28358 112680 28364
rect 112352 28144 112404 28150
rect 112352 28086 112404 28092
rect 112260 28076 112312 28082
rect 112260 28018 112312 28024
rect 112260 27872 112312 27878
rect 112260 27814 112312 27820
rect 112272 27606 112300 27814
rect 112260 27600 112312 27606
rect 112260 27542 112312 27548
rect 112272 27470 112300 27542
rect 112260 27464 112312 27470
rect 112260 27406 112312 27412
rect 112168 27328 112220 27334
rect 112168 27270 112220 27276
rect 112180 27062 112208 27270
rect 112168 27056 112220 27062
rect 112168 26998 112220 27004
rect 110972 26988 111024 26994
rect 110972 26930 111024 26936
rect 111248 26988 111300 26994
rect 111248 26930 111300 26936
rect 111340 26988 111392 26994
rect 111340 26930 111392 26936
rect 112076 26988 112128 26994
rect 112076 26930 112128 26936
rect 111260 26586 111288 26930
rect 112364 26926 112392 28086
rect 112640 28082 112668 28358
rect 113376 28218 113404 29242
rect 113468 29238 113496 30790
rect 113836 30734 113864 31282
rect 114192 31136 114244 31142
rect 114296 31124 114324 31282
rect 114388 31210 114416 31470
rect 114468 31476 114520 31482
rect 114468 31418 114520 31424
rect 114652 31340 114704 31346
rect 114652 31282 114704 31288
rect 114376 31204 114428 31210
rect 114376 31146 114428 31152
rect 114244 31096 114324 31124
rect 114560 31136 114612 31142
rect 114192 31078 114244 31084
rect 114560 31078 114612 31084
rect 114098 30832 114154 30841
rect 114098 30767 114154 30776
rect 114284 30796 114336 30802
rect 113824 30728 113876 30734
rect 113822 30696 113824 30705
rect 113876 30696 113878 30705
rect 113548 30660 113600 30666
rect 113822 30631 113878 30640
rect 113548 30602 113600 30608
rect 113560 30394 113588 30602
rect 114008 30592 114060 30598
rect 114008 30534 114060 30540
rect 113650 30492 113958 30501
rect 113650 30490 113656 30492
rect 113712 30490 113736 30492
rect 113792 30490 113816 30492
rect 113872 30490 113896 30492
rect 113952 30490 113958 30492
rect 113712 30438 113714 30490
rect 113894 30438 113896 30490
rect 113650 30436 113656 30438
rect 113712 30436 113736 30438
rect 113792 30436 113816 30438
rect 113872 30436 113896 30438
rect 113952 30436 113958 30438
rect 113650 30427 113958 30436
rect 113548 30388 113600 30394
rect 113548 30330 113600 30336
rect 114020 30274 114048 30534
rect 113744 30258 114048 30274
rect 113732 30252 114048 30258
rect 113784 30246 114048 30252
rect 113732 30194 113784 30200
rect 114112 29714 114140 30767
rect 114468 30796 114520 30802
rect 114336 30756 114468 30784
rect 114284 30738 114336 30744
rect 114468 30738 114520 30744
rect 114572 30326 114600 31078
rect 114664 30938 114692 31282
rect 114848 31142 114876 33458
rect 114940 32230 114968 33895
rect 115124 33658 115152 34478
rect 115308 33969 115336 34886
rect 115294 33960 115350 33969
rect 115294 33895 115350 33904
rect 115112 33652 115164 33658
rect 115112 33594 115164 33600
rect 115204 33652 115256 33658
rect 115204 33594 115256 33600
rect 115216 33114 115244 33594
rect 115400 33318 115428 36246
rect 115756 36168 115808 36174
rect 115860 36156 115888 36722
rect 116136 36242 116164 36722
rect 116124 36236 116176 36242
rect 116124 36178 116176 36184
rect 115808 36128 115888 36156
rect 115756 36110 115808 36116
rect 115480 36100 115532 36106
rect 115480 36042 115532 36048
rect 115492 35698 115520 36042
rect 115480 35692 115532 35698
rect 115480 35634 115532 35640
rect 115940 35624 115992 35630
rect 115940 35566 115992 35572
rect 116032 35624 116084 35630
rect 116032 35566 116084 35572
rect 115572 35556 115624 35562
rect 115572 35498 115624 35504
rect 115480 35080 115532 35086
rect 115480 35022 115532 35028
rect 115492 34678 115520 35022
rect 115480 34672 115532 34678
rect 115480 34614 115532 34620
rect 115584 34542 115612 35498
rect 115662 34640 115718 34649
rect 115662 34575 115664 34584
rect 115716 34575 115718 34584
rect 115664 34546 115716 34552
rect 115572 34536 115624 34542
rect 115572 34478 115624 34484
rect 115584 33862 115612 34478
rect 115572 33856 115624 33862
rect 115572 33798 115624 33804
rect 115584 33658 115612 33798
rect 115572 33652 115624 33658
rect 115572 33594 115624 33600
rect 115756 33584 115808 33590
rect 115756 33526 115808 33532
rect 115846 33552 115902 33561
rect 115664 33516 115716 33522
rect 115664 33458 115716 33464
rect 115480 33380 115532 33386
rect 115480 33322 115532 33328
rect 115388 33312 115440 33318
rect 115388 33254 115440 33260
rect 115204 33108 115256 33114
rect 115204 33050 115256 33056
rect 115020 32904 115072 32910
rect 115020 32846 115072 32852
rect 115294 32872 115350 32881
rect 114928 32224 114980 32230
rect 114928 32166 114980 32172
rect 114928 31816 114980 31822
rect 114928 31758 114980 31764
rect 114836 31136 114888 31142
rect 114836 31078 114888 31084
rect 114652 30932 114704 30938
rect 114652 30874 114704 30880
rect 114652 30728 114704 30734
rect 114650 30696 114652 30705
rect 114704 30696 114706 30705
rect 114650 30631 114706 30640
rect 114560 30320 114612 30326
rect 114560 30262 114612 30268
rect 114192 30184 114244 30190
rect 114192 30126 114244 30132
rect 114204 29850 114232 30126
rect 114192 29844 114244 29850
rect 114192 29786 114244 29792
rect 114100 29708 114152 29714
rect 114100 29650 114152 29656
rect 113650 29404 113958 29413
rect 113650 29402 113656 29404
rect 113712 29402 113736 29404
rect 113792 29402 113816 29404
rect 113872 29402 113896 29404
rect 113952 29402 113958 29404
rect 113712 29350 113714 29402
rect 113894 29350 113896 29402
rect 113650 29348 113656 29350
rect 113712 29348 113736 29350
rect 113792 29348 113816 29350
rect 113872 29348 113896 29350
rect 113952 29348 113958 29350
rect 113650 29339 113958 29348
rect 113456 29232 113508 29238
rect 113456 29174 113508 29180
rect 113732 29164 113784 29170
rect 113732 29106 113784 29112
rect 113744 28762 113772 29106
rect 114008 29096 114060 29102
rect 114112 29084 114140 29650
rect 114204 29170 114232 29786
rect 114744 29504 114796 29510
rect 114744 29446 114796 29452
rect 114192 29164 114244 29170
rect 114192 29106 114244 29112
rect 114060 29056 114140 29084
rect 114008 29038 114060 29044
rect 113456 28756 113508 28762
rect 113456 28698 113508 28704
rect 113732 28756 113784 28762
rect 113732 28698 113784 28704
rect 114100 28756 114152 28762
rect 114100 28698 114152 28704
rect 113468 28490 113496 28698
rect 113548 28552 113600 28558
rect 113548 28494 113600 28500
rect 113456 28484 113508 28490
rect 113456 28426 113508 28432
rect 113560 28422 113588 28494
rect 113548 28416 113600 28422
rect 113548 28358 113600 28364
rect 113560 28218 113588 28358
rect 113650 28316 113958 28325
rect 113650 28314 113656 28316
rect 113712 28314 113736 28316
rect 113792 28314 113816 28316
rect 113872 28314 113896 28316
rect 113952 28314 113958 28316
rect 113712 28262 113714 28314
rect 113894 28262 113896 28314
rect 113650 28260 113656 28262
rect 113712 28260 113736 28262
rect 113792 28260 113816 28262
rect 113872 28260 113896 28262
rect 113952 28260 113958 28262
rect 113650 28251 113958 28260
rect 113364 28212 113416 28218
rect 113364 28154 113416 28160
rect 113548 28212 113600 28218
rect 113548 28154 113600 28160
rect 114008 28144 114060 28150
rect 114008 28086 114060 28092
rect 112628 28076 112680 28082
rect 112628 28018 112680 28024
rect 113272 28076 113324 28082
rect 113272 28018 113324 28024
rect 112914 27772 113222 27781
rect 112914 27770 112920 27772
rect 112976 27770 113000 27772
rect 113056 27770 113080 27772
rect 113136 27770 113160 27772
rect 113216 27770 113222 27772
rect 112976 27718 112978 27770
rect 113158 27718 113160 27770
rect 112914 27716 112920 27718
rect 112976 27716 113000 27718
rect 113056 27716 113080 27718
rect 113136 27716 113160 27718
rect 113216 27716 113222 27718
rect 112914 27707 113222 27716
rect 113284 27538 113312 28018
rect 113548 27600 113600 27606
rect 113548 27542 113600 27548
rect 113272 27532 113324 27538
rect 113272 27474 113324 27480
rect 112536 27396 112588 27402
rect 112536 27338 112588 27344
rect 112720 27396 112772 27402
rect 112720 27338 112772 27344
rect 112548 27062 112576 27338
rect 112536 27056 112588 27062
rect 112536 26998 112588 27004
rect 112352 26920 112404 26926
rect 112352 26862 112404 26868
rect 111248 26580 111300 26586
rect 111248 26522 111300 26528
rect 112548 26382 112576 26998
rect 112732 26450 112760 27338
rect 113560 26994 113588 27542
rect 113650 27228 113958 27237
rect 113650 27226 113656 27228
rect 113712 27226 113736 27228
rect 113792 27226 113816 27228
rect 113872 27226 113896 27228
rect 113952 27226 113958 27228
rect 113712 27174 113714 27226
rect 113894 27174 113896 27226
rect 113650 27172 113656 27174
rect 113712 27172 113736 27174
rect 113792 27172 113816 27174
rect 113872 27172 113896 27174
rect 113952 27172 113958 27174
rect 113650 27163 113958 27172
rect 114020 27130 114048 28086
rect 114112 28014 114140 28698
rect 114756 28642 114784 29446
rect 114388 28626 114784 28642
rect 114848 28626 114876 31078
rect 114940 30802 114968 31758
rect 114928 30796 114980 30802
rect 114928 30738 114980 30744
rect 114928 30388 114980 30394
rect 114928 30330 114980 30336
rect 114940 29646 114968 30330
rect 115032 30122 115060 32846
rect 115294 32807 115296 32816
rect 115348 32807 115350 32816
rect 115296 32778 115348 32784
rect 115492 32774 115520 33322
rect 115480 32768 115532 32774
rect 115480 32710 115532 32716
rect 115676 32570 115704 33458
rect 115768 32978 115796 33526
rect 115846 33487 115902 33496
rect 115756 32972 115808 32978
rect 115756 32914 115808 32920
rect 115860 32910 115888 33487
rect 115952 32910 115980 35566
rect 116044 34542 116072 35566
rect 116320 35170 116348 37198
rect 116412 36854 116440 37266
rect 116492 37120 116544 37126
rect 116492 37062 116544 37068
rect 116400 36848 116452 36854
rect 116400 36790 116452 36796
rect 116504 36786 116532 37062
rect 116492 36780 116544 36786
rect 116492 36722 116544 36728
rect 116952 36780 117004 36786
rect 116952 36722 117004 36728
rect 116504 36106 116532 36722
rect 116964 36378 116992 36722
rect 117136 36712 117188 36718
rect 117136 36654 117188 36660
rect 116952 36372 117004 36378
rect 116952 36314 117004 36320
rect 117148 36174 117176 36654
rect 117412 36236 117464 36242
rect 117412 36178 117464 36184
rect 116860 36168 116912 36174
rect 116860 36110 116912 36116
rect 116952 36168 117004 36174
rect 116952 36110 117004 36116
rect 117136 36168 117188 36174
rect 117136 36110 117188 36116
rect 116492 36100 116544 36106
rect 116492 36042 116544 36048
rect 116584 35692 116636 35698
rect 116872 35680 116900 36110
rect 116964 35834 116992 36110
rect 116952 35828 117004 35834
rect 116952 35770 117004 35776
rect 117044 35692 117096 35698
rect 116872 35652 117044 35680
rect 116584 35634 116636 35640
rect 117044 35634 117096 35640
rect 116596 35290 116624 35634
rect 116584 35284 116636 35290
rect 116584 35226 116636 35232
rect 116124 35148 116176 35154
rect 116320 35142 116440 35170
rect 116124 35090 116176 35096
rect 116136 34746 116164 35090
rect 116308 35080 116360 35086
rect 116308 35022 116360 35028
rect 116124 34740 116176 34746
rect 116124 34682 116176 34688
rect 116032 34536 116084 34542
rect 116032 34478 116084 34484
rect 116320 34066 116348 35022
rect 116308 34060 116360 34066
rect 116308 34002 116360 34008
rect 116032 33992 116084 33998
rect 116124 33992 116176 33998
rect 116032 33934 116084 33940
rect 116122 33960 116124 33969
rect 116176 33960 116178 33969
rect 116044 33454 116072 33934
rect 116122 33895 116178 33904
rect 116308 33652 116360 33658
rect 116308 33594 116360 33600
rect 116216 33584 116268 33590
rect 116214 33552 116216 33561
rect 116268 33552 116270 33561
rect 116214 33487 116270 33496
rect 116032 33448 116084 33454
rect 116032 33390 116084 33396
rect 116124 33448 116176 33454
rect 116124 33390 116176 33396
rect 116044 33114 116072 33390
rect 116032 33108 116084 33114
rect 116032 33050 116084 33056
rect 115848 32904 115900 32910
rect 115848 32846 115900 32852
rect 115940 32904 115992 32910
rect 115940 32846 115992 32852
rect 115848 32768 115900 32774
rect 115848 32710 115900 32716
rect 115664 32564 115716 32570
rect 115664 32506 115716 32512
rect 115388 32428 115440 32434
rect 115388 32370 115440 32376
rect 115204 32360 115256 32366
rect 115204 32302 115256 32308
rect 115112 32224 115164 32230
rect 115112 32166 115164 32172
rect 115124 31414 115152 32166
rect 115216 31958 115244 32302
rect 115400 32026 115428 32370
rect 115860 32366 115888 32710
rect 115952 32416 115980 32846
rect 116136 32570 116164 33390
rect 116216 32904 116268 32910
rect 116216 32846 116268 32852
rect 116228 32570 116256 32846
rect 116124 32564 116176 32570
rect 116124 32506 116176 32512
rect 116216 32564 116268 32570
rect 116216 32506 116268 32512
rect 116320 32434 116348 33594
rect 116412 32910 116440 35142
rect 116492 35012 116544 35018
rect 116492 34954 116544 34960
rect 116504 34202 116532 34954
rect 117056 34406 117084 35634
rect 117148 35018 117176 36110
rect 117320 36032 117372 36038
rect 117320 35974 117372 35980
rect 117332 35290 117360 35974
rect 117424 35834 117452 36178
rect 117412 35828 117464 35834
rect 117412 35770 117464 35776
rect 118240 35692 118292 35698
rect 118240 35634 118292 35640
rect 117872 35624 117924 35630
rect 117872 35566 117924 35572
rect 117320 35284 117372 35290
rect 117320 35226 117372 35232
rect 117596 35148 117648 35154
rect 117596 35090 117648 35096
rect 117136 35012 117188 35018
rect 117136 34954 117188 34960
rect 117228 34944 117280 34950
rect 117228 34886 117280 34892
rect 117240 34610 117268 34886
rect 117228 34604 117280 34610
rect 117228 34546 117280 34552
rect 117504 34604 117556 34610
rect 117504 34546 117556 34552
rect 117412 34468 117464 34474
rect 117412 34410 117464 34416
rect 117044 34400 117096 34406
rect 117044 34342 117096 34348
rect 116492 34196 116544 34202
rect 116492 34138 116544 34144
rect 116504 33998 116532 34138
rect 117056 34134 117084 34342
rect 117424 34202 117452 34410
rect 117412 34196 117464 34202
rect 117412 34138 117464 34144
rect 117044 34128 117096 34134
rect 117044 34070 117096 34076
rect 116492 33992 116544 33998
rect 116492 33934 116544 33940
rect 116400 32904 116452 32910
rect 116504 32881 116532 33934
rect 117516 33658 117544 34546
rect 117608 33930 117636 35090
rect 117884 34950 117912 35566
rect 118252 35494 118280 35634
rect 118240 35488 118292 35494
rect 118240 35430 118292 35436
rect 118252 35290 118280 35430
rect 118240 35284 118292 35290
rect 118240 35226 118292 35232
rect 117964 35012 118016 35018
rect 117964 34954 118016 34960
rect 118148 35012 118200 35018
rect 118148 34954 118200 34960
rect 118332 35012 118384 35018
rect 118332 34954 118384 34960
rect 117872 34944 117924 34950
rect 117872 34886 117924 34892
rect 117688 34604 117740 34610
rect 117688 34546 117740 34552
rect 117700 34202 117728 34546
rect 117780 34536 117832 34542
rect 117780 34478 117832 34484
rect 117688 34196 117740 34202
rect 117688 34138 117740 34144
rect 117792 34066 117820 34478
rect 117780 34060 117832 34066
rect 117780 34002 117832 34008
rect 117976 33998 118004 34954
rect 118160 34474 118188 34954
rect 118344 34542 118372 34954
rect 118332 34536 118384 34542
rect 118332 34478 118384 34484
rect 118148 34468 118200 34474
rect 118148 34410 118200 34416
rect 117964 33992 118016 33998
rect 117964 33934 118016 33940
rect 117596 33924 117648 33930
rect 117596 33866 117648 33872
rect 117504 33652 117556 33658
rect 117504 33594 117556 33600
rect 117136 33448 117188 33454
rect 117136 33390 117188 33396
rect 116676 33380 116728 33386
rect 116676 33322 116728 33328
rect 116688 33114 116716 33322
rect 116952 33312 117004 33318
rect 116952 33254 117004 33260
rect 116676 33108 116728 33114
rect 116676 33050 116728 33056
rect 116400 32846 116452 32852
rect 116490 32872 116546 32881
rect 116308 32428 116360 32434
rect 115952 32388 116072 32416
rect 115480 32360 115532 32366
rect 115480 32302 115532 32308
rect 115848 32360 115900 32366
rect 115848 32302 115900 32308
rect 116044 32314 116072 32388
rect 116308 32370 116360 32376
rect 116216 32360 116268 32366
rect 115492 32026 115520 32302
rect 115940 32292 115992 32298
rect 116044 32286 116164 32314
rect 116216 32302 116268 32308
rect 115940 32234 115992 32240
rect 115388 32020 115440 32026
rect 115388 31962 115440 31968
rect 115480 32020 115532 32026
rect 115480 31962 115532 31968
rect 115204 31952 115256 31958
rect 115204 31894 115256 31900
rect 115754 31920 115810 31929
rect 115952 31890 115980 32234
rect 116032 32020 116084 32026
rect 116032 31962 116084 31968
rect 115754 31855 115810 31864
rect 115940 31884 115992 31890
rect 115768 31822 115796 31855
rect 115940 31826 115992 31832
rect 115756 31816 115808 31822
rect 115756 31758 115808 31764
rect 115952 31686 115980 31826
rect 115848 31680 115900 31686
rect 115848 31622 115900 31628
rect 115940 31680 115992 31686
rect 115940 31622 115992 31628
rect 115860 31498 115888 31622
rect 115860 31470 115980 31498
rect 115112 31408 115164 31414
rect 115112 31350 115164 31356
rect 115952 31346 115980 31470
rect 115940 31340 115992 31346
rect 115940 31282 115992 31288
rect 115112 30864 115164 30870
rect 115110 30832 115112 30841
rect 115164 30832 115166 30841
rect 115952 30818 115980 31282
rect 116044 30938 116072 31962
rect 116136 31793 116164 32286
rect 116228 32230 116256 32302
rect 116216 32224 116268 32230
rect 116216 32166 116268 32172
rect 116308 32224 116360 32230
rect 116308 32166 116360 32172
rect 116122 31784 116178 31793
rect 116320 31754 116348 32166
rect 116412 31890 116440 32846
rect 116490 32807 116546 32816
rect 116400 31884 116452 31890
rect 116400 31826 116452 31832
rect 116504 31754 116532 32807
rect 116766 32464 116822 32473
rect 116964 32434 116992 33254
rect 117148 33046 117176 33390
rect 117608 33114 117636 33866
rect 117688 33448 117740 33454
rect 117688 33390 117740 33396
rect 117700 33114 117728 33390
rect 117976 33386 118004 33934
rect 117964 33380 118016 33386
rect 117964 33322 118016 33328
rect 117780 33312 117832 33318
rect 117780 33254 117832 33260
rect 117596 33108 117648 33114
rect 117596 33050 117648 33056
rect 117688 33108 117740 33114
rect 117688 33050 117740 33056
rect 117136 33040 117188 33046
rect 117136 32982 117188 32988
rect 117688 32904 117740 32910
rect 117688 32846 117740 32852
rect 117136 32768 117188 32774
rect 117136 32710 117188 32716
rect 117228 32768 117280 32774
rect 117228 32710 117280 32716
rect 116766 32399 116768 32408
rect 116820 32399 116822 32408
rect 116860 32428 116912 32434
rect 116768 32370 116820 32376
rect 116860 32370 116912 32376
rect 116952 32428 117004 32434
rect 116952 32370 117004 32376
rect 116584 32360 116636 32366
rect 116582 32328 116584 32337
rect 116636 32328 116638 32337
rect 116582 32263 116638 32272
rect 116122 31719 116178 31728
rect 116216 31748 116268 31754
rect 116136 31482 116164 31719
rect 116320 31726 116532 31754
rect 116216 31690 116268 31696
rect 116124 31476 116176 31482
rect 116124 31418 116176 31424
rect 116032 30932 116084 30938
rect 116032 30874 116084 30880
rect 115110 30767 115166 30776
rect 115480 30796 115532 30802
rect 115952 30790 116072 30818
rect 115480 30738 115532 30744
rect 115020 30116 115072 30122
rect 115020 30058 115072 30064
rect 115388 30048 115440 30054
rect 115388 29990 115440 29996
rect 115400 29646 115428 29990
rect 114928 29640 114980 29646
rect 114928 29582 114980 29588
rect 115296 29640 115348 29646
rect 115296 29582 115348 29588
rect 115388 29640 115440 29646
rect 115388 29582 115440 29588
rect 115112 29504 115164 29510
rect 115112 29446 115164 29452
rect 115124 29170 115152 29446
rect 114928 29164 114980 29170
rect 114928 29106 114980 29112
rect 115112 29164 115164 29170
rect 115112 29106 115164 29112
rect 114940 28762 114968 29106
rect 115112 29028 115164 29034
rect 115112 28970 115164 28976
rect 114928 28756 114980 28762
rect 114928 28698 114980 28704
rect 114388 28620 114796 28626
rect 114388 28614 114744 28620
rect 114388 28558 114416 28614
rect 114376 28552 114428 28558
rect 114376 28494 114428 28500
rect 114468 28552 114520 28558
rect 114468 28494 114520 28500
rect 114376 28212 114428 28218
rect 114376 28154 114428 28160
rect 114100 28008 114152 28014
rect 114100 27950 114152 27956
rect 114112 27538 114140 27950
rect 114388 27946 114416 28154
rect 114480 28082 114508 28494
rect 114572 28082 114600 28614
rect 114744 28562 114796 28568
rect 114836 28620 114888 28626
rect 114836 28562 114888 28568
rect 115020 28620 115072 28626
rect 115020 28562 115072 28568
rect 115032 28506 115060 28562
rect 115124 28558 115152 28970
rect 115308 28558 115336 29582
rect 115492 29170 115520 30738
rect 116044 30734 116072 30790
rect 116032 30728 116084 30734
rect 116032 30670 116084 30676
rect 115940 30660 115992 30666
rect 115940 30602 115992 30608
rect 115952 30138 115980 30602
rect 116044 30190 116072 30670
rect 115768 30110 115980 30138
rect 116032 30184 116084 30190
rect 116032 30126 116084 30132
rect 115768 30054 115796 30110
rect 115756 30048 115808 30054
rect 115756 29990 115808 29996
rect 115848 30048 115900 30054
rect 115848 29990 115900 29996
rect 115860 29646 115888 29990
rect 115848 29640 115900 29646
rect 115848 29582 115900 29588
rect 115940 29504 115992 29510
rect 115940 29446 115992 29452
rect 115952 29170 115980 29446
rect 115480 29164 115532 29170
rect 115480 29106 115532 29112
rect 115940 29164 115992 29170
rect 115940 29106 115992 29112
rect 115492 28966 115520 29106
rect 115480 28960 115532 28966
rect 115480 28902 115532 28908
rect 115492 28626 115520 28902
rect 115940 28688 115992 28694
rect 115940 28630 115992 28636
rect 115480 28620 115532 28626
rect 115480 28562 115532 28568
rect 114848 28478 115060 28506
rect 115112 28552 115164 28558
rect 115112 28494 115164 28500
rect 115296 28552 115348 28558
rect 115296 28494 115348 28500
rect 114744 28144 114796 28150
rect 114744 28086 114796 28092
rect 114468 28076 114520 28082
rect 114468 28018 114520 28024
rect 114560 28076 114612 28082
rect 114560 28018 114612 28024
rect 114376 27940 114428 27946
rect 114376 27882 114428 27888
rect 114480 27674 114508 28018
rect 114468 27668 114520 27674
rect 114468 27610 114520 27616
rect 114100 27532 114152 27538
rect 114100 27474 114152 27480
rect 114652 27464 114704 27470
rect 114652 27406 114704 27412
rect 114100 27328 114152 27334
rect 114100 27270 114152 27276
rect 114008 27124 114060 27130
rect 114008 27066 114060 27072
rect 113548 26988 113600 26994
rect 113548 26930 113600 26936
rect 112914 26684 113222 26693
rect 112914 26682 112920 26684
rect 112976 26682 113000 26684
rect 113056 26682 113080 26684
rect 113136 26682 113160 26684
rect 113216 26682 113222 26684
rect 112976 26630 112978 26682
rect 113158 26630 113160 26682
rect 112914 26628 112920 26630
rect 112976 26628 113000 26630
rect 113056 26628 113080 26630
rect 113136 26628 113160 26630
rect 113216 26628 113222 26630
rect 112914 26619 113222 26628
rect 114112 26586 114140 27270
rect 114664 26926 114692 27406
rect 114756 26994 114784 28086
rect 114848 28082 114876 28478
rect 114928 28416 114980 28422
rect 114928 28358 114980 28364
rect 115572 28416 115624 28422
rect 115572 28358 115624 28364
rect 114836 28076 114888 28082
rect 114836 28018 114888 28024
rect 114848 27130 114876 28018
rect 114940 27470 114968 28358
rect 115584 28082 115612 28358
rect 115572 28076 115624 28082
rect 115572 28018 115624 28024
rect 115020 27872 115072 27878
rect 115020 27814 115072 27820
rect 115032 27470 115060 27814
rect 115296 27532 115348 27538
rect 115296 27474 115348 27480
rect 114928 27464 114980 27470
rect 114928 27406 114980 27412
rect 115020 27464 115072 27470
rect 115020 27406 115072 27412
rect 115308 27130 115336 27474
rect 115952 27470 115980 28630
rect 116044 28218 116072 30126
rect 116124 30048 116176 30054
rect 116228 30036 116256 31690
rect 116504 31346 116532 31726
rect 116596 31482 116624 32263
rect 116872 31958 116900 32370
rect 117148 32026 117176 32710
rect 117136 32020 117188 32026
rect 117136 31962 117188 31968
rect 116860 31952 116912 31958
rect 116860 31894 116912 31900
rect 116952 31816 117004 31822
rect 116952 31758 117004 31764
rect 117134 31784 117190 31793
rect 116676 31680 116728 31686
rect 116676 31622 116728 31628
rect 116584 31476 116636 31482
rect 116584 31418 116636 31424
rect 116688 31346 116716 31622
rect 116964 31414 116992 31758
rect 117134 31719 117190 31728
rect 116768 31408 116820 31414
rect 116768 31350 116820 31356
rect 116952 31408 117004 31414
rect 116952 31350 117004 31356
rect 116400 31340 116452 31346
rect 116400 31282 116452 31288
rect 116492 31340 116544 31346
rect 116492 31282 116544 31288
rect 116676 31340 116728 31346
rect 116676 31282 116728 31288
rect 116308 31136 116360 31142
rect 116308 31078 116360 31084
rect 116320 30326 116348 31078
rect 116412 30870 116440 31282
rect 116584 31272 116636 31278
rect 116584 31214 116636 31220
rect 116596 30938 116624 31214
rect 116584 30932 116636 30938
rect 116584 30874 116636 30880
rect 116400 30864 116452 30870
rect 116400 30806 116452 30812
rect 116400 30728 116452 30734
rect 116400 30670 116452 30676
rect 116308 30320 116360 30326
rect 116308 30262 116360 30268
rect 116412 30258 116440 30670
rect 116492 30592 116544 30598
rect 116492 30534 116544 30540
rect 116584 30592 116636 30598
rect 116584 30534 116636 30540
rect 116504 30258 116532 30534
rect 116596 30258 116624 30534
rect 116400 30252 116452 30258
rect 116400 30194 116452 30200
rect 116492 30252 116544 30258
rect 116492 30194 116544 30200
rect 116584 30252 116636 30258
rect 116584 30194 116636 30200
rect 116176 30008 116256 30036
rect 116124 29990 116176 29996
rect 116136 28694 116164 29990
rect 116216 29300 116268 29306
rect 116216 29242 116268 29248
rect 116124 28688 116176 28694
rect 116124 28630 116176 28636
rect 116228 28558 116256 29242
rect 116412 29152 116440 30194
rect 116504 29714 116532 30194
rect 116584 30048 116636 30054
rect 116584 29990 116636 29996
rect 116492 29708 116544 29714
rect 116492 29650 116544 29656
rect 116596 29646 116624 29990
rect 116584 29640 116636 29646
rect 116584 29582 116636 29588
rect 116780 29578 116808 31350
rect 117148 31226 117176 31719
rect 117240 31686 117268 32710
rect 117700 32570 117728 32846
rect 117596 32564 117648 32570
rect 117596 32506 117648 32512
rect 117688 32564 117740 32570
rect 117688 32506 117740 32512
rect 117318 32464 117374 32473
rect 117318 32399 117320 32408
rect 117372 32399 117374 32408
rect 117504 32428 117556 32434
rect 117320 32370 117372 32376
rect 117504 32370 117556 32376
rect 117332 31890 117360 32370
rect 117516 32337 117544 32370
rect 117502 32328 117558 32337
rect 117412 32292 117464 32298
rect 117502 32263 117558 32272
rect 117412 32234 117464 32240
rect 117320 31884 117372 31890
rect 117320 31826 117372 31832
rect 117424 31754 117452 32234
rect 117608 31958 117636 32506
rect 117792 32434 117820 33254
rect 118148 32972 118200 32978
rect 118148 32914 118200 32920
rect 118160 32570 118188 32914
rect 118148 32564 118200 32570
rect 118148 32506 118200 32512
rect 117780 32428 117832 32434
rect 117780 32370 117832 32376
rect 118514 32056 118570 32065
rect 118514 31991 118570 32000
rect 117596 31952 117648 31958
rect 117596 31894 117648 31900
rect 117608 31822 117636 31894
rect 118528 31822 118556 31991
rect 117596 31816 117648 31822
rect 117596 31758 117648 31764
rect 118516 31816 118568 31822
rect 118516 31758 118568 31764
rect 117424 31726 117544 31754
rect 117228 31680 117280 31686
rect 117228 31622 117280 31628
rect 117412 31340 117464 31346
rect 117412 31282 117464 31288
rect 117056 31198 117268 31226
rect 116860 30864 116912 30870
rect 116860 30806 116912 30812
rect 116872 30326 116900 30806
rect 116952 30728 117004 30734
rect 116952 30670 117004 30676
rect 116860 30320 116912 30326
rect 116860 30262 116912 30268
rect 116872 30122 116900 30262
rect 116964 30258 116992 30670
rect 116952 30252 117004 30258
rect 116952 30194 117004 30200
rect 116860 30116 116912 30122
rect 116860 30058 116912 30064
rect 116768 29572 116820 29578
rect 116768 29514 116820 29520
rect 116780 29170 116808 29514
rect 116860 29504 116912 29510
rect 116860 29446 116912 29452
rect 116872 29238 116900 29446
rect 116952 29300 117004 29306
rect 116952 29242 117004 29248
rect 116860 29232 116912 29238
rect 116860 29174 116912 29180
rect 116492 29164 116544 29170
rect 116412 29124 116492 29152
rect 116492 29106 116544 29112
rect 116768 29164 116820 29170
rect 116768 29106 116820 29112
rect 116964 28966 116992 29242
rect 116676 28960 116728 28966
rect 116676 28902 116728 28908
rect 116860 28960 116912 28966
rect 116860 28902 116912 28908
rect 116952 28960 117004 28966
rect 116952 28902 117004 28908
rect 116216 28552 116268 28558
rect 116216 28494 116268 28500
rect 116032 28212 116084 28218
rect 116032 28154 116084 28160
rect 116584 28212 116636 28218
rect 116584 28154 116636 28160
rect 116596 28082 116624 28154
rect 116688 28082 116716 28902
rect 116872 28082 116900 28902
rect 117056 28490 117084 31198
rect 117136 31136 117188 31142
rect 117136 31078 117188 31084
rect 117148 30938 117176 31078
rect 117240 30954 117268 31198
rect 117240 30938 117360 30954
rect 117136 30932 117188 30938
rect 117240 30932 117372 30938
rect 117240 30926 117320 30932
rect 117136 30874 117188 30880
rect 117320 30874 117372 30880
rect 117148 30682 117176 30874
rect 117148 30654 117268 30682
rect 117136 30592 117188 30598
rect 117136 30534 117188 30540
rect 117148 30394 117176 30534
rect 117136 30388 117188 30394
rect 117136 30330 117188 30336
rect 117240 30258 117268 30654
rect 117228 30252 117280 30258
rect 117228 30194 117280 30200
rect 117424 30138 117452 31282
rect 117332 30110 117452 30138
rect 117332 29510 117360 30110
rect 117412 30048 117464 30054
rect 117412 29990 117464 29996
rect 117320 29504 117372 29510
rect 117320 29446 117372 29452
rect 117424 29306 117452 29990
rect 117516 29782 117544 31726
rect 117964 31748 118016 31754
rect 117964 31690 118016 31696
rect 117976 31482 118004 31690
rect 118332 31680 118384 31686
rect 118332 31622 118384 31628
rect 117780 31476 117832 31482
rect 117780 31418 117832 31424
rect 117964 31476 118016 31482
rect 117964 31418 118016 31424
rect 117596 30592 117648 30598
rect 117596 30534 117648 30540
rect 117608 30326 117636 30534
rect 117596 30320 117648 30326
rect 117596 30262 117648 30268
rect 117504 29776 117556 29782
rect 117504 29718 117556 29724
rect 117608 29646 117636 30262
rect 117792 30258 117820 31418
rect 117964 31204 118016 31210
rect 117964 31146 118016 31152
rect 117976 30734 118004 31146
rect 118344 30734 118372 31622
rect 118514 31376 118570 31385
rect 118514 31311 118516 31320
rect 118568 31311 118570 31320
rect 118516 31282 118568 31288
rect 117964 30728 118016 30734
rect 117964 30670 118016 30676
rect 118332 30728 118384 30734
rect 118332 30670 118384 30676
rect 118514 30696 118570 30705
rect 117976 30410 118004 30670
rect 118514 30631 118570 30640
rect 117872 30388 117924 30394
rect 117976 30382 118188 30410
rect 117872 30330 117924 30336
rect 117780 30252 117832 30258
rect 117780 30194 117832 30200
rect 117792 29850 117820 30194
rect 117884 29850 117912 30330
rect 118056 30252 118108 30258
rect 118056 30194 118108 30200
rect 118068 30138 118096 30194
rect 117976 30110 118096 30138
rect 117780 29844 117832 29850
rect 117780 29786 117832 29792
rect 117872 29844 117924 29850
rect 117872 29786 117924 29792
rect 117596 29640 117648 29646
rect 117596 29582 117648 29588
rect 117976 29578 118004 30110
rect 118056 29640 118108 29646
rect 118056 29582 118108 29588
rect 117780 29572 117832 29578
rect 117780 29514 117832 29520
rect 117964 29572 118016 29578
rect 117964 29514 118016 29520
rect 117504 29504 117556 29510
rect 117504 29446 117556 29452
rect 117596 29504 117648 29510
rect 117596 29446 117648 29452
rect 117412 29300 117464 29306
rect 117412 29242 117464 29248
rect 117516 29186 117544 29446
rect 117608 29238 117636 29446
rect 117320 29164 117372 29170
rect 117320 29106 117372 29112
rect 117424 29158 117544 29186
rect 117596 29232 117648 29238
rect 117596 29174 117648 29180
rect 117332 28665 117360 29106
rect 117424 29102 117452 29158
rect 117412 29096 117464 29102
rect 117412 29038 117464 29044
rect 117596 29096 117648 29102
rect 117596 29038 117648 29044
rect 117318 28656 117374 28665
rect 117318 28591 117374 28600
rect 117136 28552 117188 28558
rect 117136 28494 117188 28500
rect 117044 28484 117096 28490
rect 117044 28426 117096 28432
rect 116952 28416 117004 28422
rect 116952 28358 117004 28364
rect 116964 28082 116992 28358
rect 116124 28076 116176 28082
rect 116124 28018 116176 28024
rect 116584 28076 116636 28082
rect 116584 28018 116636 28024
rect 116676 28076 116728 28082
rect 116676 28018 116728 28024
rect 116860 28076 116912 28082
rect 116860 28018 116912 28024
rect 116952 28076 117004 28082
rect 116952 28018 117004 28024
rect 116136 27674 116164 28018
rect 116492 27872 116544 27878
rect 116492 27814 116544 27820
rect 116124 27668 116176 27674
rect 116124 27610 116176 27616
rect 115940 27464 115992 27470
rect 115940 27406 115992 27412
rect 116124 27464 116176 27470
rect 116124 27406 116176 27412
rect 115388 27396 115440 27402
rect 115388 27338 115440 27344
rect 115400 27130 115428 27338
rect 115664 27328 115716 27334
rect 115664 27270 115716 27276
rect 114836 27124 114888 27130
rect 114836 27066 114888 27072
rect 115296 27124 115348 27130
rect 115296 27066 115348 27072
rect 115388 27124 115440 27130
rect 115388 27066 115440 27072
rect 114744 26988 114796 26994
rect 114744 26930 114796 26936
rect 114652 26920 114704 26926
rect 114652 26862 114704 26868
rect 114100 26580 114152 26586
rect 114100 26522 114152 26528
rect 112720 26444 112772 26450
rect 112720 26386 112772 26392
rect 109868 26376 109920 26382
rect 109868 26318 109920 26324
rect 112536 26376 112588 26382
rect 112536 26318 112588 26324
rect 114756 26246 114784 26930
rect 115308 26738 115336 27066
rect 115676 26994 115704 27270
rect 115952 27010 115980 27406
rect 116136 27062 116164 27406
rect 116504 27402 116532 27814
rect 116596 27470 116624 28018
rect 116688 27962 116716 28018
rect 116688 27934 116808 27962
rect 116780 27538 116808 27934
rect 116768 27532 116820 27538
rect 116768 27474 116820 27480
rect 116872 27470 116900 28018
rect 117056 27674 117084 28426
rect 117148 28150 117176 28494
rect 117608 28422 117636 29038
rect 117688 29028 117740 29034
rect 117688 28970 117740 28976
rect 117596 28416 117648 28422
rect 117596 28358 117648 28364
rect 117136 28144 117188 28150
rect 117136 28086 117188 28092
rect 117412 28008 117464 28014
rect 117412 27950 117464 27956
rect 117044 27668 117096 27674
rect 117044 27610 117096 27616
rect 117424 27606 117452 27950
rect 117412 27600 117464 27606
rect 117412 27542 117464 27548
rect 117608 27538 117636 28358
rect 117700 28082 117728 28970
rect 117792 28558 117820 29514
rect 117780 28552 117832 28558
rect 117780 28494 117832 28500
rect 117976 28490 118004 29514
rect 118068 28762 118096 29582
rect 118160 29510 118188 30382
rect 118528 30326 118556 30631
rect 118516 30320 118568 30326
rect 118516 30262 118568 30268
rect 118332 29776 118384 29782
rect 118332 29718 118384 29724
rect 118148 29504 118200 29510
rect 118148 29446 118200 29452
rect 118238 29336 118294 29345
rect 118238 29271 118294 29280
rect 118148 29028 118200 29034
rect 118148 28970 118200 28976
rect 118056 28756 118108 28762
rect 118056 28698 118108 28704
rect 117964 28484 118016 28490
rect 117964 28426 118016 28432
rect 117780 28416 117832 28422
rect 117780 28358 117832 28364
rect 117792 28218 117820 28358
rect 117780 28212 117832 28218
rect 117780 28154 117832 28160
rect 117688 28076 117740 28082
rect 117688 28018 117740 28024
rect 117596 27532 117648 27538
rect 117596 27474 117648 27480
rect 118160 27470 118188 28970
rect 118252 28558 118280 29271
rect 118240 28552 118292 28558
rect 118240 28494 118292 28500
rect 118252 28218 118280 28494
rect 118240 28212 118292 28218
rect 118240 28154 118292 28160
rect 118240 28076 118292 28082
rect 118240 28018 118292 28024
rect 118252 27985 118280 28018
rect 118238 27976 118294 27985
rect 118238 27911 118294 27920
rect 118252 27674 118280 27911
rect 118240 27668 118292 27674
rect 118240 27610 118292 27616
rect 118344 27606 118372 29718
rect 118528 29646 118556 30262
rect 118606 30016 118662 30025
rect 118606 29951 118662 29960
rect 118516 29640 118568 29646
rect 118516 29582 118568 29588
rect 118516 29028 118568 29034
rect 118516 28970 118568 28976
rect 118528 28665 118556 28970
rect 118514 28656 118570 28665
rect 118514 28591 118570 28600
rect 118620 28558 118648 29951
rect 118608 28552 118660 28558
rect 118608 28494 118660 28500
rect 118332 27600 118384 27606
rect 118332 27542 118384 27548
rect 116584 27464 116636 27470
rect 116584 27406 116636 27412
rect 116860 27464 116912 27470
rect 116860 27406 116912 27412
rect 118148 27464 118200 27470
rect 118148 27406 118200 27412
rect 118516 27464 118568 27470
rect 118516 27406 118568 27412
rect 116492 27396 116544 27402
rect 116492 27338 116544 27344
rect 118528 27305 118556 27406
rect 118514 27296 118570 27305
rect 118514 27231 118570 27240
rect 118528 27130 118556 27231
rect 118516 27124 118568 27130
rect 118516 27066 118568 27072
rect 115860 26994 115980 27010
rect 116124 27056 116176 27062
rect 116124 26998 116176 27004
rect 115664 26988 115716 26994
rect 115664 26930 115716 26936
rect 115848 26988 115980 26994
rect 115900 26982 115980 26988
rect 115848 26930 115900 26936
rect 115848 26784 115900 26790
rect 115308 26710 115428 26738
rect 115848 26726 115900 26732
rect 115296 26580 115348 26586
rect 115296 26522 115348 26528
rect 115020 26308 115072 26314
rect 115020 26250 115072 26256
rect 114744 26240 114796 26246
rect 114744 26182 114796 26188
rect 113650 26140 113958 26149
rect 113650 26138 113656 26140
rect 113712 26138 113736 26140
rect 113792 26138 113816 26140
rect 113872 26138 113896 26140
rect 113952 26138 113958 26140
rect 113712 26086 113714 26138
rect 113894 26086 113896 26138
rect 113650 26084 113656 26086
rect 113712 26084 113736 26086
rect 113792 26084 113816 26086
rect 113872 26084 113896 26086
rect 113952 26084 113958 26086
rect 113650 26075 113958 26084
rect 114756 25974 114784 26182
rect 114744 25968 114796 25974
rect 114744 25910 114796 25916
rect 115032 25770 115060 26250
rect 115308 25906 115336 26522
rect 115400 26314 115428 26710
rect 115860 26586 115888 26726
rect 115848 26580 115900 26586
rect 115848 26522 115900 26528
rect 115388 26308 115440 26314
rect 115388 26250 115440 26256
rect 115400 26042 115428 26250
rect 115388 26036 115440 26042
rect 115388 25978 115440 25984
rect 115296 25900 115348 25906
rect 115296 25842 115348 25848
rect 115020 25764 115072 25770
rect 115020 25706 115072 25712
rect 112914 25596 113222 25605
rect 112914 25594 112920 25596
rect 112976 25594 113000 25596
rect 113056 25594 113080 25596
rect 113136 25594 113160 25596
rect 113216 25594 113222 25596
rect 112976 25542 112978 25594
rect 113158 25542 113160 25594
rect 112914 25540 112920 25542
rect 112976 25540 113000 25542
rect 113056 25540 113080 25542
rect 113136 25540 113160 25542
rect 113216 25540 113222 25542
rect 112914 25531 113222 25540
rect 113650 25052 113958 25061
rect 113650 25050 113656 25052
rect 113712 25050 113736 25052
rect 113792 25050 113816 25052
rect 113872 25050 113896 25052
rect 113952 25050 113958 25052
rect 113712 24998 113714 25050
rect 113894 24998 113896 25050
rect 113650 24996 113656 24998
rect 113712 24996 113736 24998
rect 113792 24996 113816 24998
rect 113872 24996 113896 24998
rect 113952 24996 113958 24998
rect 113650 24987 113958 24996
rect 112914 24508 113222 24517
rect 112914 24506 112920 24508
rect 112976 24506 113000 24508
rect 113056 24506 113080 24508
rect 113136 24506 113160 24508
rect 113216 24506 113222 24508
rect 112976 24454 112978 24506
rect 113158 24454 113160 24506
rect 112914 24452 112920 24454
rect 112976 24452 113000 24454
rect 113056 24452 113080 24454
rect 113136 24452 113160 24454
rect 113216 24452 113222 24454
rect 112914 24443 113222 24452
rect 113650 23964 113958 23973
rect 113650 23962 113656 23964
rect 113712 23962 113736 23964
rect 113792 23962 113816 23964
rect 113872 23962 113896 23964
rect 113952 23962 113958 23964
rect 113712 23910 113714 23962
rect 113894 23910 113896 23962
rect 113650 23908 113656 23910
rect 113712 23908 113736 23910
rect 113792 23908 113816 23910
rect 113872 23908 113896 23910
rect 113952 23908 113958 23910
rect 113650 23899 113958 23908
rect 112914 23420 113222 23429
rect 112914 23418 112920 23420
rect 112976 23418 113000 23420
rect 113056 23418 113080 23420
rect 113136 23418 113160 23420
rect 113216 23418 113222 23420
rect 112976 23366 112978 23418
rect 113158 23366 113160 23418
rect 112914 23364 112920 23366
rect 112976 23364 113000 23366
rect 113056 23364 113080 23366
rect 113136 23364 113160 23366
rect 113216 23364 113222 23366
rect 112914 23355 113222 23364
rect 113650 22876 113958 22885
rect 113650 22874 113656 22876
rect 113712 22874 113736 22876
rect 113792 22874 113816 22876
rect 113872 22874 113896 22876
rect 113952 22874 113958 22876
rect 113712 22822 113714 22874
rect 113894 22822 113896 22874
rect 113650 22820 113656 22822
rect 113712 22820 113736 22822
rect 113792 22820 113816 22822
rect 113872 22820 113896 22822
rect 113952 22820 113958 22822
rect 113650 22811 113958 22820
rect 112914 22332 113222 22341
rect 112914 22330 112920 22332
rect 112976 22330 113000 22332
rect 113056 22330 113080 22332
rect 113136 22330 113160 22332
rect 113216 22330 113222 22332
rect 112976 22278 112978 22330
rect 113158 22278 113160 22330
rect 112914 22276 112920 22278
rect 112976 22276 113000 22278
rect 113056 22276 113080 22278
rect 113136 22276 113160 22278
rect 113216 22276 113222 22278
rect 112914 22267 113222 22276
rect 113650 21788 113958 21797
rect 113650 21786 113656 21788
rect 113712 21786 113736 21788
rect 113792 21786 113816 21788
rect 113872 21786 113896 21788
rect 113952 21786 113958 21788
rect 113712 21734 113714 21786
rect 113894 21734 113896 21786
rect 113650 21732 113656 21734
rect 113712 21732 113736 21734
rect 113792 21732 113816 21734
rect 113872 21732 113896 21734
rect 113952 21732 113958 21734
rect 113650 21723 113958 21732
rect 112914 21244 113222 21253
rect 112914 21242 112920 21244
rect 112976 21242 113000 21244
rect 113056 21242 113080 21244
rect 113136 21242 113160 21244
rect 113216 21242 113222 21244
rect 112976 21190 112978 21242
rect 113158 21190 113160 21242
rect 112914 21188 112920 21190
rect 112976 21188 113000 21190
rect 113056 21188 113080 21190
rect 113136 21188 113160 21190
rect 113216 21188 113222 21190
rect 112914 21179 113222 21188
rect 113650 20700 113958 20709
rect 113650 20698 113656 20700
rect 113712 20698 113736 20700
rect 113792 20698 113816 20700
rect 113872 20698 113896 20700
rect 113952 20698 113958 20700
rect 113712 20646 113714 20698
rect 113894 20646 113896 20698
rect 113650 20644 113656 20646
rect 113712 20644 113736 20646
rect 113792 20644 113816 20646
rect 113872 20644 113896 20646
rect 113952 20644 113958 20646
rect 113650 20635 113958 20644
rect 112914 20156 113222 20165
rect 112914 20154 112920 20156
rect 112976 20154 113000 20156
rect 113056 20154 113080 20156
rect 113136 20154 113160 20156
rect 113216 20154 113222 20156
rect 112976 20102 112978 20154
rect 113158 20102 113160 20154
rect 112914 20100 112920 20102
rect 112976 20100 113000 20102
rect 113056 20100 113080 20102
rect 113136 20100 113160 20102
rect 113216 20100 113222 20102
rect 112914 20091 113222 20100
rect 113650 19612 113958 19621
rect 113650 19610 113656 19612
rect 113712 19610 113736 19612
rect 113792 19610 113816 19612
rect 113872 19610 113896 19612
rect 113952 19610 113958 19612
rect 113712 19558 113714 19610
rect 113894 19558 113896 19610
rect 113650 19556 113656 19558
rect 113712 19556 113736 19558
rect 113792 19556 113816 19558
rect 113872 19556 113896 19558
rect 113952 19556 113958 19558
rect 113650 19547 113958 19556
rect 112914 19068 113222 19077
rect 112914 19066 112920 19068
rect 112976 19066 113000 19068
rect 113056 19066 113080 19068
rect 113136 19066 113160 19068
rect 113216 19066 113222 19068
rect 112976 19014 112978 19066
rect 113158 19014 113160 19066
rect 112914 19012 112920 19014
rect 112976 19012 113000 19014
rect 113056 19012 113080 19014
rect 113136 19012 113160 19014
rect 113216 19012 113222 19014
rect 112914 19003 113222 19012
rect 113650 18524 113958 18533
rect 113650 18522 113656 18524
rect 113712 18522 113736 18524
rect 113792 18522 113816 18524
rect 113872 18522 113896 18524
rect 113952 18522 113958 18524
rect 113712 18470 113714 18522
rect 113894 18470 113896 18522
rect 113650 18468 113656 18470
rect 113712 18468 113736 18470
rect 113792 18468 113816 18470
rect 113872 18468 113896 18470
rect 113952 18468 113958 18470
rect 113650 18459 113958 18468
rect 112914 17980 113222 17989
rect 112914 17978 112920 17980
rect 112976 17978 113000 17980
rect 113056 17978 113080 17980
rect 113136 17978 113160 17980
rect 113216 17978 113222 17980
rect 112976 17926 112978 17978
rect 113158 17926 113160 17978
rect 112914 17924 112920 17926
rect 112976 17924 113000 17926
rect 113056 17924 113080 17926
rect 113136 17924 113160 17926
rect 113216 17924 113222 17926
rect 112914 17915 113222 17924
rect 113650 17436 113958 17445
rect 113650 17434 113656 17436
rect 113712 17434 113736 17436
rect 113792 17434 113816 17436
rect 113872 17434 113896 17436
rect 113952 17434 113958 17436
rect 113712 17382 113714 17434
rect 113894 17382 113896 17434
rect 113650 17380 113656 17382
rect 113712 17380 113736 17382
rect 113792 17380 113816 17382
rect 113872 17380 113896 17382
rect 113952 17380 113958 17382
rect 113650 17371 113958 17380
rect 112914 16892 113222 16901
rect 112914 16890 112920 16892
rect 112976 16890 113000 16892
rect 113056 16890 113080 16892
rect 113136 16890 113160 16892
rect 113216 16890 113222 16892
rect 112976 16838 112978 16890
rect 113158 16838 113160 16890
rect 112914 16836 112920 16838
rect 112976 16836 113000 16838
rect 113056 16836 113080 16838
rect 113136 16836 113160 16838
rect 113216 16836 113222 16838
rect 112914 16827 113222 16836
rect 113650 16348 113958 16357
rect 113650 16346 113656 16348
rect 113712 16346 113736 16348
rect 113792 16346 113816 16348
rect 113872 16346 113896 16348
rect 113952 16346 113958 16348
rect 113712 16294 113714 16346
rect 113894 16294 113896 16346
rect 113650 16292 113656 16294
rect 113712 16292 113736 16294
rect 113792 16292 113816 16294
rect 113872 16292 113896 16294
rect 113952 16292 113958 16294
rect 113650 16283 113958 16292
rect 112914 15804 113222 15813
rect 112914 15802 112920 15804
rect 112976 15802 113000 15804
rect 113056 15802 113080 15804
rect 113136 15802 113160 15804
rect 113216 15802 113222 15804
rect 112976 15750 112978 15802
rect 113158 15750 113160 15802
rect 112914 15748 112920 15750
rect 112976 15748 113000 15750
rect 113056 15748 113080 15750
rect 113136 15748 113160 15750
rect 113216 15748 113222 15750
rect 112914 15739 113222 15748
rect 113650 15260 113958 15269
rect 113650 15258 113656 15260
rect 113712 15258 113736 15260
rect 113792 15258 113816 15260
rect 113872 15258 113896 15260
rect 113952 15258 113958 15260
rect 113712 15206 113714 15258
rect 113894 15206 113896 15258
rect 113650 15204 113656 15206
rect 113712 15204 113736 15206
rect 113792 15204 113816 15206
rect 113872 15204 113896 15206
rect 113952 15204 113958 15206
rect 113650 15195 113958 15204
rect 112914 14716 113222 14725
rect 112914 14714 112920 14716
rect 112976 14714 113000 14716
rect 113056 14714 113080 14716
rect 113136 14714 113160 14716
rect 113216 14714 113222 14716
rect 112976 14662 112978 14714
rect 113158 14662 113160 14714
rect 112914 14660 112920 14662
rect 112976 14660 113000 14662
rect 113056 14660 113080 14662
rect 113136 14660 113160 14662
rect 113216 14660 113222 14662
rect 112914 14651 113222 14660
rect 113650 14172 113958 14181
rect 113650 14170 113656 14172
rect 113712 14170 113736 14172
rect 113792 14170 113816 14172
rect 113872 14170 113896 14172
rect 113952 14170 113958 14172
rect 113712 14118 113714 14170
rect 113894 14118 113896 14170
rect 113650 14116 113656 14118
rect 113712 14116 113736 14118
rect 113792 14116 113816 14118
rect 113872 14116 113896 14118
rect 113952 14116 113958 14118
rect 113650 14107 113958 14116
rect 112914 13628 113222 13637
rect 112914 13626 112920 13628
rect 112976 13626 113000 13628
rect 113056 13626 113080 13628
rect 113136 13626 113160 13628
rect 113216 13626 113222 13628
rect 112976 13574 112978 13626
rect 113158 13574 113160 13626
rect 112914 13572 112920 13574
rect 112976 13572 113000 13574
rect 113056 13572 113080 13574
rect 113136 13572 113160 13574
rect 113216 13572 113222 13574
rect 112914 13563 113222 13572
rect 113650 13084 113958 13093
rect 113650 13082 113656 13084
rect 113712 13082 113736 13084
rect 113792 13082 113816 13084
rect 113872 13082 113896 13084
rect 113952 13082 113958 13084
rect 113712 13030 113714 13082
rect 113894 13030 113896 13082
rect 113650 13028 113656 13030
rect 113712 13028 113736 13030
rect 113792 13028 113816 13030
rect 113872 13028 113896 13030
rect 113952 13028 113958 13030
rect 113650 13019 113958 13028
rect 112914 12540 113222 12549
rect 112914 12538 112920 12540
rect 112976 12538 113000 12540
rect 113056 12538 113080 12540
rect 113136 12538 113160 12540
rect 113216 12538 113222 12540
rect 112976 12486 112978 12538
rect 113158 12486 113160 12538
rect 112914 12484 112920 12486
rect 112976 12484 113000 12486
rect 113056 12484 113080 12486
rect 113136 12484 113160 12486
rect 113216 12484 113222 12486
rect 112914 12475 113222 12484
rect 113650 11996 113958 12005
rect 113650 11994 113656 11996
rect 113712 11994 113736 11996
rect 113792 11994 113816 11996
rect 113872 11994 113896 11996
rect 113952 11994 113958 11996
rect 113712 11942 113714 11994
rect 113894 11942 113896 11994
rect 113650 11940 113656 11942
rect 113712 11940 113736 11942
rect 113792 11940 113816 11942
rect 113872 11940 113896 11942
rect 113952 11940 113958 11942
rect 113650 11931 113958 11940
rect 112914 11452 113222 11461
rect 112914 11450 112920 11452
rect 112976 11450 113000 11452
rect 113056 11450 113080 11452
rect 113136 11450 113160 11452
rect 113216 11450 113222 11452
rect 112976 11398 112978 11450
rect 113158 11398 113160 11450
rect 112914 11396 112920 11398
rect 112976 11396 113000 11398
rect 113056 11396 113080 11398
rect 113136 11396 113160 11398
rect 113216 11396 113222 11398
rect 112914 11387 113222 11396
rect 113650 10908 113958 10917
rect 113650 10906 113656 10908
rect 113712 10906 113736 10908
rect 113792 10906 113816 10908
rect 113872 10906 113896 10908
rect 113952 10906 113958 10908
rect 113712 10854 113714 10906
rect 113894 10854 113896 10906
rect 113650 10852 113656 10854
rect 113712 10852 113736 10854
rect 113792 10852 113816 10854
rect 113872 10852 113896 10854
rect 113952 10852 113958 10854
rect 113650 10843 113958 10852
rect 112914 10364 113222 10373
rect 112914 10362 112920 10364
rect 112976 10362 113000 10364
rect 113056 10362 113080 10364
rect 113136 10362 113160 10364
rect 113216 10362 113222 10364
rect 112976 10310 112978 10362
rect 113158 10310 113160 10362
rect 112914 10308 112920 10310
rect 112976 10308 113000 10310
rect 113056 10308 113080 10310
rect 113136 10308 113160 10310
rect 113216 10308 113222 10310
rect 112914 10299 113222 10308
rect 109500 10056 109552 10062
rect 108762 10024 108818 10033
rect 108304 9988 108356 9994
rect 109500 9998 109552 10004
rect 108762 9959 108818 9968
rect 108304 9930 108356 9936
rect 106464 9920 106516 9926
rect 93032 9862 93084 9868
rect 93398 9888 93454 9897
rect 92754 9823 92810 9832
rect 15856 9654 15884 9823
rect 26974 9752 27030 9761
rect 26974 9687 27030 9696
rect 27802 9752 27858 9761
rect 27802 9687 27858 9696
rect 29550 9752 29606 9761
rect 29550 9687 29606 9696
rect 30194 9752 30250 9761
rect 30194 9687 30250 9696
rect 51630 9752 51686 9761
rect 51630 9687 51686 9696
rect 52458 9752 52514 9761
rect 52458 9687 52514 9696
rect 53562 9752 53618 9761
rect 53562 9687 53618 9696
rect 55034 9752 55090 9761
rect 55034 9687 55090 9696
rect 56138 9752 56194 9761
rect 56138 9687 56194 9696
rect 57426 9752 57482 9761
rect 57426 9687 57482 9696
rect 58254 9752 58310 9761
rect 58254 9687 58310 9696
rect 59542 9752 59598 9761
rect 59542 9687 59598 9696
rect 60830 9752 60886 9761
rect 60830 9687 60886 9696
rect 67730 9752 67786 9761
rect 67730 9687 67786 9696
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 15856 7546 15884 9590
rect 25870 8256 25926 8265
rect 25870 8191 25926 8200
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 25884 2650 25912 8191
rect 26988 7546 27016 9687
rect 27816 7546 27844 9687
rect 29564 7546 29592 9687
rect 30208 7546 30236 9687
rect 31666 8256 31722 8265
rect 31666 8191 31722 8200
rect 32954 8256 33010 8265
rect 32954 8191 33010 8200
rect 33782 8256 33838 8265
rect 33782 8191 33838 8200
rect 34794 8256 34850 8265
rect 34794 8191 34850 8200
rect 36174 8256 36230 8265
rect 36174 8191 36230 8200
rect 37462 8256 37518 8265
rect 37462 8191 37518 8200
rect 38290 8256 38346 8265
rect 38290 8191 38346 8200
rect 40866 8256 40922 8265
rect 40866 8191 40922 8200
rect 41970 8256 42026 8265
rect 41970 8191 42026 8200
rect 43258 8256 43314 8265
rect 43258 8191 43314 8200
rect 44546 8256 44602 8265
rect 44546 8191 44602 8200
rect 46662 8256 46718 8265
rect 46662 8191 46718 8200
rect 47766 8256 47822 8265
rect 47766 8191 47822 8200
rect 49054 8256 49110 8265
rect 49054 8191 49110 8200
rect 50342 8256 50398 8265
rect 50342 8191 50398 8200
rect 26976 7540 27028 7546
rect 26976 7482 27028 7488
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 30196 7540 30248 7546
rect 30196 7482 30248 7488
rect 31680 2650 31708 8191
rect 32968 2650 32996 8191
rect 33796 2650 33824 8191
rect 34808 2650 34836 8191
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 36188 2650 36216 8191
rect 37476 2650 37504 8191
rect 38304 2650 38332 8191
rect 40038 2680 40094 2689
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 32956 2644 33008 2650
rect 32956 2586 33008 2592
rect 33784 2644 33836 2650
rect 33784 2586 33836 2592
rect 34796 2644 34848 2650
rect 34796 2586 34848 2592
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 38292 2644 38344 2650
rect 40880 2650 40908 8191
rect 41984 2650 42012 8191
rect 43272 2650 43300 8191
rect 44560 2650 44588 8191
rect 45834 7168 45890 7177
rect 45834 7103 45890 7112
rect 45848 2650 45876 7103
rect 46676 2650 46704 8191
rect 47780 2650 47808 8191
rect 49068 2650 49096 8191
rect 50356 2650 50384 8191
rect 51644 2650 51672 9687
rect 52472 2650 52500 9687
rect 53576 2650 53604 9687
rect 55048 2650 55076 9687
rect 56152 2650 56180 9687
rect 57440 2650 57468 9687
rect 58268 2650 58296 9687
rect 59556 2650 59584 9687
rect 60844 2650 60872 9687
rect 61934 8256 61990 8265
rect 61934 8191 61990 8200
rect 63222 8256 63278 8265
rect 63222 8191 63278 8200
rect 64050 8256 64106 8265
rect 64050 8191 64106 8200
rect 65338 8256 65394 8265
rect 65338 8191 65394 8200
rect 66718 8256 66774 8265
rect 66718 8191 66774 8200
rect 61948 2650 61976 8191
rect 63236 2650 63264 8191
rect 64064 2650 64092 8191
rect 65352 2650 65380 8191
rect 66314 7644 66622 7653
rect 66314 7642 66320 7644
rect 66376 7642 66400 7644
rect 66456 7642 66480 7644
rect 66536 7642 66560 7644
rect 66616 7642 66622 7644
rect 66376 7590 66378 7642
rect 66558 7590 66560 7642
rect 66314 7588 66320 7590
rect 66376 7588 66400 7590
rect 66456 7588 66480 7590
rect 66536 7588 66560 7590
rect 66616 7588 66622 7590
rect 66314 7579 66622 7588
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 66314 6556 66622 6565
rect 66314 6554 66320 6556
rect 66376 6554 66400 6556
rect 66456 6554 66480 6556
rect 66536 6554 66560 6556
rect 66616 6554 66622 6556
rect 66376 6502 66378 6554
rect 66558 6502 66560 6554
rect 66314 6500 66320 6502
rect 66376 6500 66400 6502
rect 66456 6500 66480 6502
rect 66536 6500 66560 6502
rect 66616 6500 66622 6502
rect 66314 6491 66622 6500
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 66314 5468 66622 5477
rect 66314 5466 66320 5468
rect 66376 5466 66400 5468
rect 66456 5466 66480 5468
rect 66536 5466 66560 5468
rect 66616 5466 66622 5468
rect 66376 5414 66378 5466
rect 66558 5414 66560 5466
rect 66314 5412 66320 5414
rect 66376 5412 66400 5414
rect 66456 5412 66480 5414
rect 66536 5412 66560 5414
rect 66616 5412 66622 5414
rect 66314 5403 66622 5412
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 66314 4380 66622 4389
rect 66314 4378 66320 4380
rect 66376 4378 66400 4380
rect 66456 4378 66480 4380
rect 66536 4378 66560 4380
rect 66616 4378 66622 4380
rect 66376 4326 66378 4378
rect 66558 4326 66560 4378
rect 66314 4324 66320 4326
rect 66376 4324 66400 4326
rect 66456 4324 66480 4326
rect 66536 4324 66560 4326
rect 66616 4324 66622 4326
rect 66314 4315 66622 4324
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 66314 3292 66622 3301
rect 66314 3290 66320 3292
rect 66376 3290 66400 3292
rect 66456 3290 66480 3292
rect 66536 3290 66560 3292
rect 66616 3290 66622 3292
rect 66376 3238 66378 3290
rect 66558 3238 66560 3290
rect 66314 3236 66320 3238
rect 66376 3236 66400 3238
rect 66456 3236 66480 3238
rect 66536 3236 66560 3238
rect 66616 3236 66622 3238
rect 66314 3227 66622 3236
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 66732 2650 66760 8191
rect 67744 2650 67772 9687
rect 92860 7546 92888 9846
rect 93044 9761 93072 9862
rect 106464 9862 106516 9868
rect 93398 9823 93454 9832
rect 93030 9752 93086 9761
rect 93030 9687 93086 9696
rect 93044 7546 93072 9687
rect 93214 8256 93270 8265
rect 93214 8191 93270 8200
rect 93228 7546 93256 8191
rect 93412 7546 93440 9823
rect 113650 9820 113958 9829
rect 113650 9818 113656 9820
rect 113712 9818 113736 9820
rect 113792 9818 113816 9820
rect 113872 9818 113896 9820
rect 113952 9818 113958 9820
rect 113712 9766 113714 9818
rect 113894 9766 113896 9818
rect 113650 9764 113656 9766
rect 113712 9764 113736 9766
rect 113792 9764 113816 9766
rect 113872 9764 113896 9766
rect 113952 9764 113958 9766
rect 113650 9755 113958 9764
rect 112914 9276 113222 9285
rect 112914 9274 112920 9276
rect 112976 9274 113000 9276
rect 113056 9274 113080 9276
rect 113136 9274 113160 9276
rect 113216 9274 113222 9276
rect 112976 9222 112978 9274
rect 113158 9222 113160 9274
rect 112914 9220 112920 9222
rect 112976 9220 113000 9222
rect 113056 9220 113080 9222
rect 113136 9220 113160 9222
rect 113216 9220 113222 9222
rect 112914 9211 113222 9220
rect 113650 8732 113958 8741
rect 113650 8730 113656 8732
rect 113712 8730 113736 8732
rect 113792 8730 113816 8732
rect 113872 8730 113896 8732
rect 113952 8730 113958 8732
rect 113712 8678 113714 8730
rect 113894 8678 113896 8730
rect 113650 8676 113656 8678
rect 113712 8676 113736 8678
rect 113792 8676 113816 8678
rect 113872 8676 113896 8678
rect 113952 8676 113958 8678
rect 113650 8667 113958 8676
rect 112914 8188 113222 8197
rect 112914 8186 112920 8188
rect 112976 8186 113000 8188
rect 113056 8186 113080 8188
rect 113136 8186 113160 8188
rect 113216 8186 113222 8188
rect 112976 8134 112978 8186
rect 113158 8134 113160 8186
rect 112914 8132 112920 8134
rect 112976 8132 113000 8134
rect 113056 8132 113080 8134
rect 113136 8132 113160 8134
rect 113216 8132 113222 8134
rect 112914 8123 113222 8132
rect 97034 7644 97342 7653
rect 97034 7642 97040 7644
rect 97096 7642 97120 7644
rect 97176 7642 97200 7644
rect 97256 7642 97280 7644
rect 97336 7642 97342 7644
rect 97096 7590 97098 7642
rect 97278 7590 97280 7642
rect 97034 7588 97040 7590
rect 97096 7588 97120 7590
rect 97176 7588 97200 7590
rect 97256 7588 97280 7590
rect 97336 7588 97342 7590
rect 97034 7579 97342 7588
rect 113650 7644 113958 7653
rect 113650 7642 113656 7644
rect 113712 7642 113736 7644
rect 113792 7642 113816 7644
rect 113872 7642 113896 7644
rect 113952 7642 113958 7644
rect 113712 7590 113714 7642
rect 113894 7590 113896 7642
rect 113650 7588 113656 7590
rect 113712 7588 113736 7590
rect 113792 7588 113816 7590
rect 113872 7588 113896 7590
rect 113952 7588 113958 7590
rect 113650 7579 113958 7588
rect 92848 7540 92900 7546
rect 92848 7482 92900 7488
rect 93032 7540 93084 7546
rect 93032 7482 93084 7488
rect 93216 7540 93268 7546
rect 93216 7482 93268 7488
rect 93400 7540 93452 7546
rect 93400 7482 93452 7488
rect 96374 7100 96682 7109
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7035 96682 7044
rect 112914 7100 113222 7109
rect 112914 7098 112920 7100
rect 112976 7098 113000 7100
rect 113056 7098 113080 7100
rect 113136 7098 113160 7100
rect 113216 7098 113222 7100
rect 112976 7046 112978 7098
rect 113158 7046 113160 7098
rect 112914 7044 112920 7046
rect 112976 7044 113000 7046
rect 113056 7044 113080 7046
rect 113136 7044 113160 7046
rect 113216 7044 113222 7046
rect 112914 7035 113222 7044
rect 97034 6556 97342 6565
rect 97034 6554 97040 6556
rect 97096 6554 97120 6556
rect 97176 6554 97200 6556
rect 97256 6554 97280 6556
rect 97336 6554 97342 6556
rect 97096 6502 97098 6554
rect 97278 6502 97280 6554
rect 97034 6500 97040 6502
rect 97096 6500 97120 6502
rect 97176 6500 97200 6502
rect 97256 6500 97280 6502
rect 97336 6500 97342 6502
rect 97034 6491 97342 6500
rect 96374 6012 96682 6021
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5947 96682 5956
rect 97034 5468 97342 5477
rect 97034 5466 97040 5468
rect 97096 5466 97120 5468
rect 97176 5466 97200 5468
rect 97256 5466 97280 5468
rect 97336 5466 97342 5468
rect 97096 5414 97098 5466
rect 97278 5414 97280 5466
rect 97034 5412 97040 5414
rect 97096 5412 97120 5414
rect 97176 5412 97200 5414
rect 97256 5412 97280 5414
rect 97336 5412 97342 5414
rect 97034 5403 97342 5412
rect 96374 4924 96682 4933
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4859 96682 4868
rect 97034 4380 97342 4389
rect 97034 4378 97040 4380
rect 97096 4378 97120 4380
rect 97176 4378 97200 4380
rect 97256 4378 97280 4380
rect 97336 4378 97342 4380
rect 97096 4326 97098 4378
rect 97278 4326 97280 4378
rect 97034 4324 97040 4326
rect 97096 4324 97120 4326
rect 97176 4324 97200 4326
rect 97256 4324 97280 4326
rect 97336 4324 97342 4326
rect 97034 4315 97342 4324
rect 96374 3836 96682 3845
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3771 96682 3780
rect 97034 3292 97342 3301
rect 97034 3290 97040 3292
rect 97096 3290 97120 3292
rect 97176 3290 97200 3292
rect 97256 3290 97280 3292
rect 97336 3290 97342 3292
rect 97096 3238 97098 3290
rect 97278 3238 97280 3290
rect 97034 3236 97040 3238
rect 97096 3236 97120 3238
rect 97176 3236 97200 3238
rect 97256 3236 97280 3238
rect 97336 3236 97342 3238
rect 97034 3227 97342 3236
rect 96374 2748 96682 2757
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2683 96682 2692
rect 40038 2615 40040 2624
rect 38292 2586 38344 2592
rect 40092 2615 40094 2624
rect 40868 2644 40920 2650
rect 40040 2586 40092 2592
rect 40868 2586 40920 2592
rect 41972 2644 42024 2650
rect 41972 2586 42024 2592
rect 43260 2644 43312 2650
rect 43260 2586 43312 2592
rect 44548 2644 44600 2650
rect 44548 2586 44600 2592
rect 45836 2644 45888 2650
rect 45836 2586 45888 2592
rect 46664 2644 46716 2650
rect 46664 2586 46716 2592
rect 47768 2644 47820 2650
rect 47768 2586 47820 2592
rect 49056 2644 49108 2650
rect 49056 2586 49108 2592
rect 50344 2644 50396 2650
rect 50344 2586 50396 2592
rect 51632 2644 51684 2650
rect 51632 2586 51684 2592
rect 52460 2644 52512 2650
rect 52460 2586 52512 2592
rect 53564 2644 53616 2650
rect 53564 2586 53616 2592
rect 55036 2644 55088 2650
rect 55036 2586 55088 2592
rect 56140 2644 56192 2650
rect 56140 2586 56192 2592
rect 57428 2644 57480 2650
rect 57428 2586 57480 2592
rect 58256 2644 58308 2650
rect 58256 2586 58308 2592
rect 59544 2644 59596 2650
rect 59544 2586 59596 2592
rect 60832 2644 60884 2650
rect 60832 2586 60884 2592
rect 61936 2644 61988 2650
rect 61936 2586 61988 2592
rect 63224 2644 63276 2650
rect 63224 2586 63276 2592
rect 64052 2644 64104 2650
rect 64052 2586 64104 2592
rect 65340 2644 65392 2650
rect 65340 2586 65392 2592
rect 66720 2644 66772 2650
rect 66720 2586 66772 2592
rect 67732 2644 67784 2650
rect 67732 2586 67784 2592
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 39948 2304 40000 2310
rect 39948 2246 40000 2252
rect 40592 2304 40644 2310
rect 40592 2246 40644 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 44456 2304 44508 2310
rect 44456 2246 44508 2252
rect 45744 2304 45796 2310
rect 45744 2246 45796 2252
rect 46388 2304 46440 2310
rect 46388 2246 46440 2252
rect 47676 2304 47728 2310
rect 47676 2246 47728 2252
rect 48964 2304 49016 2310
rect 48964 2246 49016 2252
rect 50252 2304 50304 2310
rect 50252 2246 50304 2252
rect 51540 2304 51592 2310
rect 51540 2246 51592 2252
rect 52184 2304 52236 2310
rect 52184 2246 52236 2252
rect 53472 2304 53524 2310
rect 53472 2246 53524 2252
rect 54760 2304 54812 2310
rect 54760 2246 54812 2252
rect 56048 2304 56100 2310
rect 56048 2246 56100 2252
rect 57336 2304 57388 2310
rect 57336 2246 57388 2252
rect 57980 2304 58032 2310
rect 57980 2246 58032 2252
rect 59268 2304 59320 2310
rect 59268 2246 59320 2252
rect 60556 2304 60608 2310
rect 60556 2246 60608 2252
rect 61844 2304 61896 2310
rect 61844 2246 61896 2252
rect 63132 2304 63184 2310
rect 63132 2246 63184 2252
rect 63776 2304 63828 2310
rect 63776 2246 63828 2252
rect 65064 2304 65116 2310
rect 65064 2246 65116 2252
rect 66720 2304 66772 2310
rect 66720 2246 66772 2252
rect 67640 2304 67692 2310
rect 67640 2246 67692 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 25792 800 25820 2246
rect 31588 800 31616 2246
rect 32876 800 32904 2246
rect 33520 800 33548 2246
rect 34808 800 34836 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36096 800 36124 2246
rect 37384 800 37412 2246
rect 38028 800 38056 2246
rect 39960 800 39988 2246
rect 40604 800 40632 2246
rect 41892 800 41920 2246
rect 43180 800 43208 2246
rect 44468 800 44496 2246
rect 45756 800 45784 2246
rect 46400 800 46428 2246
rect 47688 800 47716 2246
rect 48976 800 49004 2246
rect 50264 800 50292 2246
rect 51552 800 51580 2246
rect 52196 800 52224 2246
rect 53484 800 53512 2246
rect 54772 800 54800 2246
rect 56060 800 56088 2246
rect 57348 800 57376 2246
rect 57992 800 58020 2246
rect 59280 800 59308 2246
rect 60568 800 60596 2246
rect 61856 800 61884 2246
rect 63144 800 63172 2246
rect 63788 800 63816 2246
rect 65076 800 65104 2246
rect 66314 2204 66622 2213
rect 66314 2202 66320 2204
rect 66376 2202 66400 2204
rect 66456 2202 66480 2204
rect 66536 2202 66560 2204
rect 66616 2202 66622 2204
rect 66376 2150 66378 2202
rect 66558 2150 66560 2202
rect 66314 2148 66320 2150
rect 66376 2148 66400 2150
rect 66456 2148 66480 2150
rect 66536 2148 66560 2150
rect 66616 2148 66622 2150
rect 66314 2139 66622 2148
rect 66364 870 66484 898
rect 66364 800 66392 870
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 25778 0 25834 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 44454 0 44510 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 47674 0 47730 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 51538 0 51594 800
rect 52182 0 52238 800
rect 53470 0 53526 800
rect 54758 0 54814 800
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 57978 0 58034 800
rect 59266 0 59322 800
rect 60554 0 60610 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 63774 0 63830 800
rect 65062 0 65118 800
rect 66350 0 66406 800
rect 66456 762 66484 870
rect 66732 762 66760 2246
rect 67652 800 67680 2246
rect 97034 2204 97342 2213
rect 97034 2202 97040 2204
rect 97096 2202 97120 2204
rect 97176 2202 97200 2204
rect 97256 2202 97280 2204
rect 97336 2202 97342 2204
rect 97096 2150 97098 2202
rect 97278 2150 97280 2202
rect 97034 2148 97040 2150
rect 97096 2148 97120 2150
rect 97176 2148 97200 2150
rect 97256 2148 97280 2150
rect 97336 2148 97342 2150
rect 97034 2139 97342 2148
rect 66456 734 66760 762
rect 67638 0 67694 800
<< via2 >>
rect 4220 97402 4276 97404
rect 4300 97402 4356 97404
rect 4380 97402 4436 97404
rect 4460 97402 4516 97404
rect 4220 97350 4266 97402
rect 4266 97350 4276 97402
rect 4300 97350 4330 97402
rect 4330 97350 4342 97402
rect 4342 97350 4356 97402
rect 4380 97350 4394 97402
rect 4394 97350 4406 97402
rect 4406 97350 4436 97402
rect 4460 97350 4470 97402
rect 4470 97350 4516 97402
rect 4220 97348 4276 97350
rect 4300 97348 4356 97350
rect 4380 97348 4436 97350
rect 4460 97348 4516 97350
rect 34940 97402 34996 97404
rect 35020 97402 35076 97404
rect 35100 97402 35156 97404
rect 35180 97402 35236 97404
rect 34940 97350 34986 97402
rect 34986 97350 34996 97402
rect 35020 97350 35050 97402
rect 35050 97350 35062 97402
rect 35062 97350 35076 97402
rect 35100 97350 35114 97402
rect 35114 97350 35126 97402
rect 35126 97350 35156 97402
rect 35180 97350 35190 97402
rect 35190 97350 35236 97402
rect 34940 97348 34996 97350
rect 35020 97348 35076 97350
rect 35100 97348 35156 97350
rect 35180 97348 35236 97350
rect 65660 97402 65716 97404
rect 65740 97402 65796 97404
rect 65820 97402 65876 97404
rect 65900 97402 65956 97404
rect 65660 97350 65706 97402
rect 65706 97350 65716 97402
rect 65740 97350 65770 97402
rect 65770 97350 65782 97402
rect 65782 97350 65796 97402
rect 65820 97350 65834 97402
rect 65834 97350 65846 97402
rect 65846 97350 65876 97402
rect 65900 97350 65910 97402
rect 65910 97350 65956 97402
rect 65660 97348 65716 97350
rect 65740 97348 65796 97350
rect 65820 97348 65876 97350
rect 65900 97348 65956 97350
rect 4880 96858 4936 96860
rect 4960 96858 5016 96860
rect 5040 96858 5096 96860
rect 5120 96858 5176 96860
rect 4880 96806 4926 96858
rect 4926 96806 4936 96858
rect 4960 96806 4990 96858
rect 4990 96806 5002 96858
rect 5002 96806 5016 96858
rect 5040 96806 5054 96858
rect 5054 96806 5066 96858
rect 5066 96806 5096 96858
rect 5120 96806 5130 96858
rect 5130 96806 5176 96858
rect 4880 96804 4936 96806
rect 4960 96804 5016 96806
rect 5040 96804 5096 96806
rect 5120 96804 5176 96806
rect 35600 96858 35656 96860
rect 35680 96858 35736 96860
rect 35760 96858 35816 96860
rect 35840 96858 35896 96860
rect 35600 96806 35646 96858
rect 35646 96806 35656 96858
rect 35680 96806 35710 96858
rect 35710 96806 35722 96858
rect 35722 96806 35736 96858
rect 35760 96806 35774 96858
rect 35774 96806 35786 96858
rect 35786 96806 35816 96858
rect 35840 96806 35850 96858
rect 35850 96806 35896 96858
rect 35600 96804 35656 96806
rect 35680 96804 35736 96806
rect 35760 96804 35816 96806
rect 35840 96804 35896 96806
rect 4220 96314 4276 96316
rect 4300 96314 4356 96316
rect 4380 96314 4436 96316
rect 4460 96314 4516 96316
rect 4220 96262 4266 96314
rect 4266 96262 4276 96314
rect 4300 96262 4330 96314
rect 4330 96262 4342 96314
rect 4342 96262 4356 96314
rect 4380 96262 4394 96314
rect 4394 96262 4406 96314
rect 4406 96262 4436 96314
rect 4460 96262 4470 96314
rect 4470 96262 4516 96314
rect 4220 96260 4276 96262
rect 4300 96260 4356 96262
rect 4380 96260 4436 96262
rect 4460 96260 4516 96262
rect 34940 96314 34996 96316
rect 35020 96314 35076 96316
rect 35100 96314 35156 96316
rect 35180 96314 35236 96316
rect 34940 96262 34986 96314
rect 34986 96262 34996 96314
rect 35020 96262 35050 96314
rect 35050 96262 35062 96314
rect 35062 96262 35076 96314
rect 35100 96262 35114 96314
rect 35114 96262 35126 96314
rect 35126 96262 35156 96314
rect 35180 96262 35190 96314
rect 35190 96262 35236 96314
rect 34940 96260 34996 96262
rect 35020 96260 35076 96262
rect 35100 96260 35156 96262
rect 35180 96260 35236 96262
rect 4880 95770 4936 95772
rect 4960 95770 5016 95772
rect 5040 95770 5096 95772
rect 5120 95770 5176 95772
rect 4880 95718 4926 95770
rect 4926 95718 4936 95770
rect 4960 95718 4990 95770
rect 4990 95718 5002 95770
rect 5002 95718 5016 95770
rect 5040 95718 5054 95770
rect 5054 95718 5066 95770
rect 5066 95718 5096 95770
rect 5120 95718 5130 95770
rect 5130 95718 5176 95770
rect 4880 95716 4936 95718
rect 4960 95716 5016 95718
rect 5040 95716 5096 95718
rect 5120 95716 5176 95718
rect 35600 95770 35656 95772
rect 35680 95770 35736 95772
rect 35760 95770 35816 95772
rect 35840 95770 35896 95772
rect 35600 95718 35646 95770
rect 35646 95718 35656 95770
rect 35680 95718 35710 95770
rect 35710 95718 35722 95770
rect 35722 95718 35736 95770
rect 35760 95718 35774 95770
rect 35774 95718 35786 95770
rect 35786 95718 35816 95770
rect 35840 95718 35850 95770
rect 35850 95718 35896 95770
rect 35600 95716 35656 95718
rect 35680 95716 35736 95718
rect 35760 95716 35816 95718
rect 35840 95716 35896 95718
rect 4220 95226 4276 95228
rect 4300 95226 4356 95228
rect 4380 95226 4436 95228
rect 4460 95226 4516 95228
rect 4220 95174 4266 95226
rect 4266 95174 4276 95226
rect 4300 95174 4330 95226
rect 4330 95174 4342 95226
rect 4342 95174 4356 95226
rect 4380 95174 4394 95226
rect 4394 95174 4406 95226
rect 4406 95174 4436 95226
rect 4460 95174 4470 95226
rect 4470 95174 4516 95226
rect 4220 95172 4276 95174
rect 4300 95172 4356 95174
rect 4380 95172 4436 95174
rect 4460 95172 4516 95174
rect 34940 95226 34996 95228
rect 35020 95226 35076 95228
rect 35100 95226 35156 95228
rect 35180 95226 35236 95228
rect 34940 95174 34986 95226
rect 34986 95174 34996 95226
rect 35020 95174 35050 95226
rect 35050 95174 35062 95226
rect 35062 95174 35076 95226
rect 35100 95174 35114 95226
rect 35114 95174 35126 95226
rect 35126 95174 35156 95226
rect 35180 95174 35190 95226
rect 35190 95174 35236 95226
rect 34940 95172 34996 95174
rect 35020 95172 35076 95174
rect 35100 95172 35156 95174
rect 35180 95172 35236 95174
rect 4880 94682 4936 94684
rect 4960 94682 5016 94684
rect 5040 94682 5096 94684
rect 5120 94682 5176 94684
rect 4880 94630 4926 94682
rect 4926 94630 4936 94682
rect 4960 94630 4990 94682
rect 4990 94630 5002 94682
rect 5002 94630 5016 94682
rect 5040 94630 5054 94682
rect 5054 94630 5066 94682
rect 5066 94630 5096 94682
rect 5120 94630 5130 94682
rect 5130 94630 5176 94682
rect 4880 94628 4936 94630
rect 4960 94628 5016 94630
rect 5040 94628 5096 94630
rect 5120 94628 5176 94630
rect 35600 94682 35656 94684
rect 35680 94682 35736 94684
rect 35760 94682 35816 94684
rect 35840 94682 35896 94684
rect 35600 94630 35646 94682
rect 35646 94630 35656 94682
rect 35680 94630 35710 94682
rect 35710 94630 35722 94682
rect 35722 94630 35736 94682
rect 35760 94630 35774 94682
rect 35774 94630 35786 94682
rect 35786 94630 35816 94682
rect 35840 94630 35850 94682
rect 35850 94630 35896 94682
rect 35600 94628 35656 94630
rect 35680 94628 35736 94630
rect 35760 94628 35816 94630
rect 35840 94628 35896 94630
rect 4220 94138 4276 94140
rect 4300 94138 4356 94140
rect 4380 94138 4436 94140
rect 4460 94138 4516 94140
rect 4220 94086 4266 94138
rect 4266 94086 4276 94138
rect 4300 94086 4330 94138
rect 4330 94086 4342 94138
rect 4342 94086 4356 94138
rect 4380 94086 4394 94138
rect 4394 94086 4406 94138
rect 4406 94086 4436 94138
rect 4460 94086 4470 94138
rect 4470 94086 4516 94138
rect 4220 94084 4276 94086
rect 4300 94084 4356 94086
rect 4380 94084 4436 94086
rect 4460 94084 4516 94086
rect 34940 94138 34996 94140
rect 35020 94138 35076 94140
rect 35100 94138 35156 94140
rect 35180 94138 35236 94140
rect 34940 94086 34986 94138
rect 34986 94086 34996 94138
rect 35020 94086 35050 94138
rect 35050 94086 35062 94138
rect 35062 94086 35076 94138
rect 35100 94086 35114 94138
rect 35114 94086 35126 94138
rect 35126 94086 35156 94138
rect 35180 94086 35190 94138
rect 35190 94086 35236 94138
rect 34940 94084 34996 94086
rect 35020 94084 35076 94086
rect 35100 94084 35156 94086
rect 35180 94084 35236 94086
rect 4880 93594 4936 93596
rect 4960 93594 5016 93596
rect 5040 93594 5096 93596
rect 5120 93594 5176 93596
rect 4880 93542 4926 93594
rect 4926 93542 4936 93594
rect 4960 93542 4990 93594
rect 4990 93542 5002 93594
rect 5002 93542 5016 93594
rect 5040 93542 5054 93594
rect 5054 93542 5066 93594
rect 5066 93542 5096 93594
rect 5120 93542 5130 93594
rect 5130 93542 5176 93594
rect 4880 93540 4936 93542
rect 4960 93540 5016 93542
rect 5040 93540 5096 93542
rect 5120 93540 5176 93542
rect 35600 93594 35656 93596
rect 35680 93594 35736 93596
rect 35760 93594 35816 93596
rect 35840 93594 35896 93596
rect 35600 93542 35646 93594
rect 35646 93542 35656 93594
rect 35680 93542 35710 93594
rect 35710 93542 35722 93594
rect 35722 93542 35736 93594
rect 35760 93542 35774 93594
rect 35774 93542 35786 93594
rect 35786 93542 35816 93594
rect 35840 93542 35850 93594
rect 35850 93542 35896 93594
rect 35600 93540 35656 93542
rect 35680 93540 35736 93542
rect 35760 93540 35816 93542
rect 35840 93540 35896 93542
rect 4220 93050 4276 93052
rect 4300 93050 4356 93052
rect 4380 93050 4436 93052
rect 4460 93050 4516 93052
rect 4220 92998 4266 93050
rect 4266 92998 4276 93050
rect 4300 92998 4330 93050
rect 4330 92998 4342 93050
rect 4342 92998 4356 93050
rect 4380 92998 4394 93050
rect 4394 92998 4406 93050
rect 4406 92998 4436 93050
rect 4460 92998 4470 93050
rect 4470 92998 4516 93050
rect 4220 92996 4276 92998
rect 4300 92996 4356 92998
rect 4380 92996 4436 92998
rect 4460 92996 4516 92998
rect 34940 93050 34996 93052
rect 35020 93050 35076 93052
rect 35100 93050 35156 93052
rect 35180 93050 35236 93052
rect 34940 92998 34986 93050
rect 34986 92998 34996 93050
rect 35020 92998 35050 93050
rect 35050 92998 35062 93050
rect 35062 92998 35076 93050
rect 35100 92998 35114 93050
rect 35114 92998 35126 93050
rect 35126 92998 35156 93050
rect 35180 92998 35190 93050
rect 35190 92998 35236 93050
rect 34940 92996 34996 92998
rect 35020 92996 35076 92998
rect 35100 92996 35156 92998
rect 35180 92996 35236 92998
rect 49330 93220 49386 93256
rect 49330 93200 49332 93220
rect 49332 93200 49384 93220
rect 49384 93200 49386 93220
rect 44178 92520 44234 92576
rect 4880 92506 4936 92508
rect 4960 92506 5016 92508
rect 5040 92506 5096 92508
rect 5120 92506 5176 92508
rect 4880 92454 4926 92506
rect 4926 92454 4936 92506
rect 4960 92454 4990 92506
rect 4990 92454 5002 92506
rect 5002 92454 5016 92506
rect 5040 92454 5054 92506
rect 5054 92454 5066 92506
rect 5066 92454 5096 92506
rect 5120 92454 5130 92506
rect 5130 92454 5176 92506
rect 4880 92452 4936 92454
rect 4960 92452 5016 92454
rect 5040 92452 5096 92454
rect 5120 92452 5176 92454
rect 35600 92506 35656 92508
rect 35680 92506 35736 92508
rect 35760 92506 35816 92508
rect 35840 92506 35896 92508
rect 35600 92454 35646 92506
rect 35646 92454 35656 92506
rect 35680 92454 35710 92506
rect 35710 92454 35722 92506
rect 35722 92454 35736 92506
rect 35760 92454 35774 92506
rect 35774 92454 35786 92506
rect 35786 92454 35816 92506
rect 35840 92454 35850 92506
rect 35850 92454 35896 92506
rect 35600 92452 35656 92454
rect 35680 92452 35736 92454
rect 35760 92452 35816 92454
rect 35840 92452 35896 92454
rect 47122 92676 47178 92712
rect 47122 92656 47124 92676
rect 47124 92656 47176 92676
rect 47176 92656 47178 92676
rect 50618 92812 50674 92848
rect 50618 92792 50620 92812
rect 50620 92792 50672 92812
rect 50672 92792 50674 92812
rect 52550 92676 52606 92712
rect 52550 92656 52552 92676
rect 52552 92656 52604 92676
rect 52604 92656 52606 92676
rect 54022 92520 54078 92576
rect 50250 92132 50306 92168
rect 50250 92112 50252 92132
rect 50252 92112 50304 92132
rect 50304 92112 50306 92132
rect 52918 92112 52974 92168
rect 53194 92012 53196 92032
rect 53196 92012 53248 92032
rect 53248 92012 53250 92032
rect 4220 91962 4276 91964
rect 4300 91962 4356 91964
rect 4380 91962 4436 91964
rect 4460 91962 4516 91964
rect 4220 91910 4266 91962
rect 4266 91910 4276 91962
rect 4300 91910 4330 91962
rect 4330 91910 4342 91962
rect 4342 91910 4356 91962
rect 4380 91910 4394 91962
rect 4394 91910 4406 91962
rect 4406 91910 4436 91962
rect 4460 91910 4470 91962
rect 4470 91910 4516 91962
rect 4220 91908 4276 91910
rect 4300 91908 4356 91910
rect 4380 91908 4436 91910
rect 4460 91908 4516 91910
rect 4880 91418 4936 91420
rect 4960 91418 5016 91420
rect 5040 91418 5096 91420
rect 5120 91418 5176 91420
rect 4880 91366 4926 91418
rect 4926 91366 4936 91418
rect 4960 91366 4990 91418
rect 4990 91366 5002 91418
rect 5002 91366 5016 91418
rect 5040 91366 5054 91418
rect 5054 91366 5066 91418
rect 5066 91366 5096 91418
rect 5120 91366 5130 91418
rect 5130 91366 5176 91418
rect 4880 91364 4936 91366
rect 4960 91364 5016 91366
rect 5040 91364 5096 91366
rect 5120 91364 5176 91366
rect 4220 90874 4276 90876
rect 4300 90874 4356 90876
rect 4380 90874 4436 90876
rect 4460 90874 4516 90876
rect 4220 90822 4266 90874
rect 4266 90822 4276 90874
rect 4300 90822 4330 90874
rect 4330 90822 4342 90874
rect 4342 90822 4356 90874
rect 4380 90822 4394 90874
rect 4394 90822 4406 90874
rect 4406 90822 4436 90874
rect 4460 90822 4470 90874
rect 4470 90822 4516 90874
rect 4220 90820 4276 90822
rect 4300 90820 4356 90822
rect 4380 90820 4436 90822
rect 4460 90820 4516 90822
rect 4880 90330 4936 90332
rect 4960 90330 5016 90332
rect 5040 90330 5096 90332
rect 5120 90330 5176 90332
rect 4880 90278 4926 90330
rect 4926 90278 4936 90330
rect 4960 90278 4990 90330
rect 4990 90278 5002 90330
rect 5002 90278 5016 90330
rect 5040 90278 5054 90330
rect 5054 90278 5066 90330
rect 5066 90278 5096 90330
rect 5120 90278 5130 90330
rect 5130 90278 5176 90330
rect 4880 90276 4936 90278
rect 4960 90276 5016 90278
rect 5040 90276 5096 90278
rect 5120 90276 5176 90278
rect 4220 89786 4276 89788
rect 4300 89786 4356 89788
rect 4380 89786 4436 89788
rect 4460 89786 4516 89788
rect 4220 89734 4266 89786
rect 4266 89734 4276 89786
rect 4300 89734 4330 89786
rect 4330 89734 4342 89786
rect 4342 89734 4356 89786
rect 4380 89734 4394 89786
rect 4394 89734 4406 89786
rect 4406 89734 4436 89786
rect 4460 89734 4470 89786
rect 4470 89734 4516 89786
rect 4220 89732 4276 89734
rect 4300 89732 4356 89734
rect 4380 89732 4436 89734
rect 4460 89732 4516 89734
rect 4880 89242 4936 89244
rect 4960 89242 5016 89244
rect 5040 89242 5096 89244
rect 5120 89242 5176 89244
rect 4880 89190 4926 89242
rect 4926 89190 4936 89242
rect 4960 89190 4990 89242
rect 4990 89190 5002 89242
rect 5002 89190 5016 89242
rect 5040 89190 5054 89242
rect 5054 89190 5066 89242
rect 5066 89190 5096 89242
rect 5120 89190 5130 89242
rect 5130 89190 5176 89242
rect 4880 89188 4936 89190
rect 4960 89188 5016 89190
rect 5040 89188 5096 89190
rect 5120 89188 5176 89190
rect 4220 88698 4276 88700
rect 4300 88698 4356 88700
rect 4380 88698 4436 88700
rect 4460 88698 4516 88700
rect 4220 88646 4266 88698
rect 4266 88646 4276 88698
rect 4300 88646 4330 88698
rect 4330 88646 4342 88698
rect 4342 88646 4356 88698
rect 4380 88646 4394 88698
rect 4394 88646 4406 88698
rect 4406 88646 4436 88698
rect 4460 88646 4470 88698
rect 4470 88646 4516 88698
rect 4220 88644 4276 88646
rect 4300 88644 4356 88646
rect 4380 88644 4436 88646
rect 4460 88644 4516 88646
rect 4880 88154 4936 88156
rect 4960 88154 5016 88156
rect 5040 88154 5096 88156
rect 5120 88154 5176 88156
rect 4880 88102 4926 88154
rect 4926 88102 4936 88154
rect 4960 88102 4990 88154
rect 4990 88102 5002 88154
rect 5002 88102 5016 88154
rect 5040 88102 5054 88154
rect 5054 88102 5066 88154
rect 5066 88102 5096 88154
rect 5120 88102 5130 88154
rect 5130 88102 5176 88154
rect 4880 88100 4936 88102
rect 4960 88100 5016 88102
rect 5040 88100 5096 88102
rect 5120 88100 5176 88102
rect 4220 87610 4276 87612
rect 4300 87610 4356 87612
rect 4380 87610 4436 87612
rect 4460 87610 4516 87612
rect 4220 87558 4266 87610
rect 4266 87558 4276 87610
rect 4300 87558 4330 87610
rect 4330 87558 4342 87610
rect 4342 87558 4356 87610
rect 4380 87558 4394 87610
rect 4394 87558 4406 87610
rect 4406 87558 4436 87610
rect 4460 87558 4470 87610
rect 4470 87558 4516 87610
rect 4220 87556 4276 87558
rect 4300 87556 4356 87558
rect 4380 87556 4436 87558
rect 4460 87556 4516 87558
rect 4880 87066 4936 87068
rect 4960 87066 5016 87068
rect 5040 87066 5096 87068
rect 5120 87066 5176 87068
rect 4880 87014 4926 87066
rect 4926 87014 4936 87066
rect 4960 87014 4990 87066
rect 4990 87014 5002 87066
rect 5002 87014 5016 87066
rect 5040 87014 5054 87066
rect 5054 87014 5066 87066
rect 5066 87014 5096 87066
rect 5120 87014 5130 87066
rect 5130 87014 5176 87066
rect 4880 87012 4936 87014
rect 4960 87012 5016 87014
rect 5040 87012 5096 87014
rect 5120 87012 5176 87014
rect 4220 86522 4276 86524
rect 4300 86522 4356 86524
rect 4380 86522 4436 86524
rect 4460 86522 4516 86524
rect 4220 86470 4266 86522
rect 4266 86470 4276 86522
rect 4300 86470 4330 86522
rect 4330 86470 4342 86522
rect 4342 86470 4356 86522
rect 4380 86470 4394 86522
rect 4394 86470 4406 86522
rect 4406 86470 4436 86522
rect 4460 86470 4470 86522
rect 4470 86470 4516 86522
rect 4220 86468 4276 86470
rect 4300 86468 4356 86470
rect 4380 86468 4436 86470
rect 4460 86468 4516 86470
rect 4880 85978 4936 85980
rect 4960 85978 5016 85980
rect 5040 85978 5096 85980
rect 5120 85978 5176 85980
rect 4880 85926 4926 85978
rect 4926 85926 4936 85978
rect 4960 85926 4990 85978
rect 4990 85926 5002 85978
rect 5002 85926 5016 85978
rect 5040 85926 5054 85978
rect 5054 85926 5066 85978
rect 5066 85926 5096 85978
rect 5120 85926 5130 85978
rect 5130 85926 5176 85978
rect 4880 85924 4936 85926
rect 4960 85924 5016 85926
rect 5040 85924 5096 85926
rect 5120 85924 5176 85926
rect 4220 85434 4276 85436
rect 4300 85434 4356 85436
rect 4380 85434 4436 85436
rect 4460 85434 4516 85436
rect 4220 85382 4266 85434
rect 4266 85382 4276 85434
rect 4300 85382 4330 85434
rect 4330 85382 4342 85434
rect 4342 85382 4356 85434
rect 4380 85382 4394 85434
rect 4394 85382 4406 85434
rect 4406 85382 4436 85434
rect 4460 85382 4470 85434
rect 4470 85382 4516 85434
rect 4220 85380 4276 85382
rect 4300 85380 4356 85382
rect 4380 85380 4436 85382
rect 4460 85380 4516 85382
rect 4880 84890 4936 84892
rect 4960 84890 5016 84892
rect 5040 84890 5096 84892
rect 5120 84890 5176 84892
rect 4880 84838 4926 84890
rect 4926 84838 4936 84890
rect 4960 84838 4990 84890
rect 4990 84838 5002 84890
rect 5002 84838 5016 84890
rect 5040 84838 5054 84890
rect 5054 84838 5066 84890
rect 5066 84838 5096 84890
rect 5120 84838 5130 84890
rect 5130 84838 5176 84890
rect 4880 84836 4936 84838
rect 4960 84836 5016 84838
rect 5040 84836 5096 84838
rect 5120 84836 5176 84838
rect 4220 84346 4276 84348
rect 4300 84346 4356 84348
rect 4380 84346 4436 84348
rect 4460 84346 4516 84348
rect 4220 84294 4266 84346
rect 4266 84294 4276 84346
rect 4300 84294 4330 84346
rect 4330 84294 4342 84346
rect 4342 84294 4356 84346
rect 4380 84294 4394 84346
rect 4394 84294 4406 84346
rect 4406 84294 4436 84346
rect 4460 84294 4470 84346
rect 4470 84294 4516 84346
rect 4220 84292 4276 84294
rect 4300 84292 4356 84294
rect 4380 84292 4436 84294
rect 4460 84292 4516 84294
rect 4880 83802 4936 83804
rect 4960 83802 5016 83804
rect 5040 83802 5096 83804
rect 5120 83802 5176 83804
rect 4880 83750 4926 83802
rect 4926 83750 4936 83802
rect 4960 83750 4990 83802
rect 4990 83750 5002 83802
rect 5002 83750 5016 83802
rect 5040 83750 5054 83802
rect 5054 83750 5066 83802
rect 5066 83750 5096 83802
rect 5120 83750 5130 83802
rect 5130 83750 5176 83802
rect 4880 83748 4936 83750
rect 4960 83748 5016 83750
rect 5040 83748 5096 83750
rect 5120 83748 5176 83750
rect 4220 83258 4276 83260
rect 4300 83258 4356 83260
rect 4380 83258 4436 83260
rect 4460 83258 4516 83260
rect 4220 83206 4266 83258
rect 4266 83206 4276 83258
rect 4300 83206 4330 83258
rect 4330 83206 4342 83258
rect 4342 83206 4356 83258
rect 4380 83206 4394 83258
rect 4394 83206 4406 83258
rect 4406 83206 4436 83258
rect 4460 83206 4470 83258
rect 4470 83206 4516 83258
rect 4220 83204 4276 83206
rect 4300 83204 4356 83206
rect 4380 83204 4436 83206
rect 4460 83204 4516 83206
rect 4880 82714 4936 82716
rect 4960 82714 5016 82716
rect 5040 82714 5096 82716
rect 5120 82714 5176 82716
rect 4880 82662 4926 82714
rect 4926 82662 4936 82714
rect 4960 82662 4990 82714
rect 4990 82662 5002 82714
rect 5002 82662 5016 82714
rect 5040 82662 5054 82714
rect 5054 82662 5066 82714
rect 5066 82662 5096 82714
rect 5120 82662 5130 82714
rect 5130 82662 5176 82714
rect 4880 82660 4936 82662
rect 4960 82660 5016 82662
rect 5040 82660 5096 82662
rect 5120 82660 5176 82662
rect 4220 82170 4276 82172
rect 4300 82170 4356 82172
rect 4380 82170 4436 82172
rect 4460 82170 4516 82172
rect 4220 82118 4266 82170
rect 4266 82118 4276 82170
rect 4300 82118 4330 82170
rect 4330 82118 4342 82170
rect 4342 82118 4356 82170
rect 4380 82118 4394 82170
rect 4394 82118 4406 82170
rect 4406 82118 4436 82170
rect 4460 82118 4470 82170
rect 4470 82118 4516 82170
rect 4220 82116 4276 82118
rect 4300 82116 4356 82118
rect 4380 82116 4436 82118
rect 4460 82116 4516 82118
rect 4880 81626 4936 81628
rect 4960 81626 5016 81628
rect 5040 81626 5096 81628
rect 5120 81626 5176 81628
rect 4880 81574 4926 81626
rect 4926 81574 4936 81626
rect 4960 81574 4990 81626
rect 4990 81574 5002 81626
rect 5002 81574 5016 81626
rect 5040 81574 5054 81626
rect 5054 81574 5066 81626
rect 5066 81574 5096 81626
rect 5120 81574 5130 81626
rect 5130 81574 5176 81626
rect 4880 81572 4936 81574
rect 4960 81572 5016 81574
rect 5040 81572 5096 81574
rect 5120 81572 5176 81574
rect 4220 81082 4276 81084
rect 4300 81082 4356 81084
rect 4380 81082 4436 81084
rect 4460 81082 4516 81084
rect 4220 81030 4266 81082
rect 4266 81030 4276 81082
rect 4300 81030 4330 81082
rect 4330 81030 4342 81082
rect 4342 81030 4356 81082
rect 4380 81030 4394 81082
rect 4394 81030 4406 81082
rect 4406 81030 4436 81082
rect 4460 81030 4470 81082
rect 4470 81030 4516 81082
rect 4220 81028 4276 81030
rect 4300 81028 4356 81030
rect 4380 81028 4436 81030
rect 4460 81028 4516 81030
rect 4880 80538 4936 80540
rect 4960 80538 5016 80540
rect 5040 80538 5096 80540
rect 5120 80538 5176 80540
rect 4880 80486 4926 80538
rect 4926 80486 4936 80538
rect 4960 80486 4990 80538
rect 4990 80486 5002 80538
rect 5002 80486 5016 80538
rect 5040 80486 5054 80538
rect 5054 80486 5066 80538
rect 5066 80486 5096 80538
rect 5120 80486 5130 80538
rect 5130 80486 5176 80538
rect 4880 80484 4936 80486
rect 4960 80484 5016 80486
rect 5040 80484 5096 80486
rect 5120 80484 5176 80486
rect 4220 79994 4276 79996
rect 4300 79994 4356 79996
rect 4380 79994 4436 79996
rect 4460 79994 4516 79996
rect 4220 79942 4266 79994
rect 4266 79942 4276 79994
rect 4300 79942 4330 79994
rect 4330 79942 4342 79994
rect 4342 79942 4356 79994
rect 4380 79942 4394 79994
rect 4394 79942 4406 79994
rect 4406 79942 4436 79994
rect 4460 79942 4470 79994
rect 4470 79942 4516 79994
rect 4220 79940 4276 79942
rect 4300 79940 4356 79942
rect 4380 79940 4436 79942
rect 4460 79940 4516 79942
rect 4880 79450 4936 79452
rect 4960 79450 5016 79452
rect 5040 79450 5096 79452
rect 5120 79450 5176 79452
rect 4880 79398 4926 79450
rect 4926 79398 4936 79450
rect 4960 79398 4990 79450
rect 4990 79398 5002 79450
rect 5002 79398 5016 79450
rect 5040 79398 5054 79450
rect 5054 79398 5066 79450
rect 5066 79398 5096 79450
rect 5120 79398 5130 79450
rect 5130 79398 5176 79450
rect 4880 79396 4936 79398
rect 4960 79396 5016 79398
rect 5040 79396 5096 79398
rect 5120 79396 5176 79398
rect 4220 78906 4276 78908
rect 4300 78906 4356 78908
rect 4380 78906 4436 78908
rect 4460 78906 4516 78908
rect 4220 78854 4266 78906
rect 4266 78854 4276 78906
rect 4300 78854 4330 78906
rect 4330 78854 4342 78906
rect 4342 78854 4356 78906
rect 4380 78854 4394 78906
rect 4394 78854 4406 78906
rect 4406 78854 4436 78906
rect 4460 78854 4470 78906
rect 4470 78854 4516 78906
rect 4220 78852 4276 78854
rect 4300 78852 4356 78854
rect 4380 78852 4436 78854
rect 4460 78852 4516 78854
rect 4880 78362 4936 78364
rect 4960 78362 5016 78364
rect 5040 78362 5096 78364
rect 5120 78362 5176 78364
rect 4880 78310 4926 78362
rect 4926 78310 4936 78362
rect 4960 78310 4990 78362
rect 4990 78310 5002 78362
rect 5002 78310 5016 78362
rect 5040 78310 5054 78362
rect 5054 78310 5066 78362
rect 5066 78310 5096 78362
rect 5120 78310 5130 78362
rect 5130 78310 5176 78362
rect 4880 78308 4936 78310
rect 4960 78308 5016 78310
rect 5040 78308 5096 78310
rect 5120 78308 5176 78310
rect 4220 77818 4276 77820
rect 4300 77818 4356 77820
rect 4380 77818 4436 77820
rect 4460 77818 4516 77820
rect 4220 77766 4266 77818
rect 4266 77766 4276 77818
rect 4300 77766 4330 77818
rect 4330 77766 4342 77818
rect 4342 77766 4356 77818
rect 4380 77766 4394 77818
rect 4394 77766 4406 77818
rect 4406 77766 4436 77818
rect 4460 77766 4470 77818
rect 4470 77766 4516 77818
rect 4220 77764 4276 77766
rect 4300 77764 4356 77766
rect 4380 77764 4436 77766
rect 4460 77764 4516 77766
rect 4880 77274 4936 77276
rect 4960 77274 5016 77276
rect 5040 77274 5096 77276
rect 5120 77274 5176 77276
rect 4880 77222 4926 77274
rect 4926 77222 4936 77274
rect 4960 77222 4990 77274
rect 4990 77222 5002 77274
rect 5002 77222 5016 77274
rect 5040 77222 5054 77274
rect 5054 77222 5066 77274
rect 5066 77222 5096 77274
rect 5120 77222 5130 77274
rect 5130 77222 5176 77274
rect 4880 77220 4936 77222
rect 4960 77220 5016 77222
rect 5040 77220 5096 77222
rect 5120 77220 5176 77222
rect 4220 76730 4276 76732
rect 4300 76730 4356 76732
rect 4380 76730 4436 76732
rect 4460 76730 4516 76732
rect 4220 76678 4266 76730
rect 4266 76678 4276 76730
rect 4300 76678 4330 76730
rect 4330 76678 4342 76730
rect 4342 76678 4356 76730
rect 4380 76678 4394 76730
rect 4394 76678 4406 76730
rect 4406 76678 4436 76730
rect 4460 76678 4470 76730
rect 4470 76678 4516 76730
rect 4220 76676 4276 76678
rect 4300 76676 4356 76678
rect 4380 76676 4436 76678
rect 4460 76676 4516 76678
rect 4880 76186 4936 76188
rect 4960 76186 5016 76188
rect 5040 76186 5096 76188
rect 5120 76186 5176 76188
rect 4880 76134 4926 76186
rect 4926 76134 4936 76186
rect 4960 76134 4990 76186
rect 4990 76134 5002 76186
rect 5002 76134 5016 76186
rect 5040 76134 5054 76186
rect 5054 76134 5066 76186
rect 5066 76134 5096 76186
rect 5120 76134 5130 76186
rect 5130 76134 5176 76186
rect 4880 76132 4936 76134
rect 4960 76132 5016 76134
rect 5040 76132 5096 76134
rect 5120 76132 5176 76134
rect 4220 75642 4276 75644
rect 4300 75642 4356 75644
rect 4380 75642 4436 75644
rect 4460 75642 4516 75644
rect 4220 75590 4266 75642
rect 4266 75590 4276 75642
rect 4300 75590 4330 75642
rect 4330 75590 4342 75642
rect 4342 75590 4356 75642
rect 4380 75590 4394 75642
rect 4394 75590 4406 75642
rect 4406 75590 4436 75642
rect 4460 75590 4470 75642
rect 4470 75590 4516 75642
rect 4220 75588 4276 75590
rect 4300 75588 4356 75590
rect 4380 75588 4436 75590
rect 4460 75588 4516 75590
rect 4880 75098 4936 75100
rect 4960 75098 5016 75100
rect 5040 75098 5096 75100
rect 5120 75098 5176 75100
rect 4880 75046 4926 75098
rect 4926 75046 4936 75098
rect 4960 75046 4990 75098
rect 4990 75046 5002 75098
rect 5002 75046 5016 75098
rect 5040 75046 5054 75098
rect 5054 75046 5066 75098
rect 5066 75046 5096 75098
rect 5120 75046 5130 75098
rect 5130 75046 5176 75098
rect 4880 75044 4936 75046
rect 4960 75044 5016 75046
rect 5040 75044 5096 75046
rect 5120 75044 5176 75046
rect 4220 74554 4276 74556
rect 4300 74554 4356 74556
rect 4380 74554 4436 74556
rect 4460 74554 4516 74556
rect 4220 74502 4266 74554
rect 4266 74502 4276 74554
rect 4300 74502 4330 74554
rect 4330 74502 4342 74554
rect 4342 74502 4356 74554
rect 4380 74502 4394 74554
rect 4394 74502 4406 74554
rect 4406 74502 4436 74554
rect 4460 74502 4470 74554
rect 4470 74502 4516 74554
rect 4220 74500 4276 74502
rect 4300 74500 4356 74502
rect 4380 74500 4436 74502
rect 4460 74500 4516 74502
rect 4880 74010 4936 74012
rect 4960 74010 5016 74012
rect 5040 74010 5096 74012
rect 5120 74010 5176 74012
rect 4880 73958 4926 74010
rect 4926 73958 4936 74010
rect 4960 73958 4990 74010
rect 4990 73958 5002 74010
rect 5002 73958 5016 74010
rect 5040 73958 5054 74010
rect 5054 73958 5066 74010
rect 5066 73958 5096 74010
rect 5120 73958 5130 74010
rect 5130 73958 5176 74010
rect 4880 73956 4936 73958
rect 4960 73956 5016 73958
rect 5040 73956 5096 73958
rect 5120 73956 5176 73958
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 4880 72922 4936 72924
rect 4960 72922 5016 72924
rect 5040 72922 5096 72924
rect 5120 72922 5176 72924
rect 4880 72870 4926 72922
rect 4926 72870 4936 72922
rect 4960 72870 4990 72922
rect 4990 72870 5002 72922
rect 5002 72870 5016 72922
rect 5040 72870 5054 72922
rect 5054 72870 5066 72922
rect 5066 72870 5096 72922
rect 5120 72870 5130 72922
rect 5130 72870 5176 72922
rect 4880 72868 4936 72870
rect 4960 72868 5016 72870
rect 5040 72868 5096 72870
rect 5120 72868 5176 72870
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 4880 71834 4936 71836
rect 4960 71834 5016 71836
rect 5040 71834 5096 71836
rect 5120 71834 5176 71836
rect 4880 71782 4926 71834
rect 4926 71782 4936 71834
rect 4960 71782 4990 71834
rect 4990 71782 5002 71834
rect 5002 71782 5016 71834
rect 5040 71782 5054 71834
rect 5054 71782 5066 71834
rect 5066 71782 5096 71834
rect 5120 71782 5130 71834
rect 5130 71782 5176 71834
rect 4880 71780 4936 71782
rect 4960 71780 5016 71782
rect 5040 71780 5096 71782
rect 5120 71780 5176 71782
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 4880 70746 4936 70748
rect 4960 70746 5016 70748
rect 5040 70746 5096 70748
rect 5120 70746 5176 70748
rect 4880 70694 4926 70746
rect 4926 70694 4936 70746
rect 4960 70694 4990 70746
rect 4990 70694 5002 70746
rect 5002 70694 5016 70746
rect 5040 70694 5054 70746
rect 5054 70694 5066 70746
rect 5066 70694 5096 70746
rect 5120 70694 5130 70746
rect 5130 70694 5176 70746
rect 4880 70692 4936 70694
rect 4960 70692 5016 70694
rect 5040 70692 5096 70694
rect 5120 70692 5176 70694
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 4880 69658 4936 69660
rect 4960 69658 5016 69660
rect 5040 69658 5096 69660
rect 5120 69658 5176 69660
rect 4880 69606 4926 69658
rect 4926 69606 4936 69658
rect 4960 69606 4990 69658
rect 4990 69606 5002 69658
rect 5002 69606 5016 69658
rect 5040 69606 5054 69658
rect 5054 69606 5066 69658
rect 5066 69606 5096 69658
rect 5120 69606 5130 69658
rect 5130 69606 5176 69658
rect 4880 69604 4936 69606
rect 4960 69604 5016 69606
rect 5040 69604 5096 69606
rect 5120 69604 5176 69606
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 4880 68570 4936 68572
rect 4960 68570 5016 68572
rect 5040 68570 5096 68572
rect 5120 68570 5176 68572
rect 4880 68518 4926 68570
rect 4926 68518 4936 68570
rect 4960 68518 4990 68570
rect 4990 68518 5002 68570
rect 5002 68518 5016 68570
rect 5040 68518 5054 68570
rect 5054 68518 5066 68570
rect 5066 68518 5096 68570
rect 5120 68518 5130 68570
rect 5130 68518 5176 68570
rect 4880 68516 4936 68518
rect 4960 68516 5016 68518
rect 5040 68516 5096 68518
rect 5120 68516 5176 68518
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4880 67482 4936 67484
rect 4960 67482 5016 67484
rect 5040 67482 5096 67484
rect 5120 67482 5176 67484
rect 4880 67430 4926 67482
rect 4926 67430 4936 67482
rect 4960 67430 4990 67482
rect 4990 67430 5002 67482
rect 5002 67430 5016 67482
rect 5040 67430 5054 67482
rect 5054 67430 5066 67482
rect 5066 67430 5096 67482
rect 5120 67430 5130 67482
rect 5130 67430 5176 67482
rect 4880 67428 4936 67430
rect 4960 67428 5016 67430
rect 5040 67428 5096 67430
rect 5120 67428 5176 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 4880 66394 4936 66396
rect 4960 66394 5016 66396
rect 5040 66394 5096 66396
rect 5120 66394 5176 66396
rect 4880 66342 4926 66394
rect 4926 66342 4936 66394
rect 4960 66342 4990 66394
rect 4990 66342 5002 66394
rect 5002 66342 5016 66394
rect 5040 66342 5054 66394
rect 5054 66342 5066 66394
rect 5066 66342 5096 66394
rect 5120 66342 5130 66394
rect 5130 66342 5176 66394
rect 4880 66340 4936 66342
rect 4960 66340 5016 66342
rect 5040 66340 5096 66342
rect 5120 66340 5176 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 4880 65306 4936 65308
rect 4960 65306 5016 65308
rect 5040 65306 5096 65308
rect 5120 65306 5176 65308
rect 4880 65254 4926 65306
rect 4926 65254 4936 65306
rect 4960 65254 4990 65306
rect 4990 65254 5002 65306
rect 5002 65254 5016 65306
rect 5040 65254 5054 65306
rect 5054 65254 5066 65306
rect 5066 65254 5096 65306
rect 5120 65254 5130 65306
rect 5130 65254 5176 65306
rect 4880 65252 4936 65254
rect 4960 65252 5016 65254
rect 5040 65252 5096 65254
rect 5120 65252 5176 65254
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4880 64218 4936 64220
rect 4960 64218 5016 64220
rect 5040 64218 5096 64220
rect 5120 64218 5176 64220
rect 4880 64166 4926 64218
rect 4926 64166 4936 64218
rect 4960 64166 4990 64218
rect 4990 64166 5002 64218
rect 5002 64166 5016 64218
rect 5040 64166 5054 64218
rect 5054 64166 5066 64218
rect 5066 64166 5096 64218
rect 5120 64166 5130 64218
rect 5130 64166 5176 64218
rect 4880 64164 4936 64166
rect 4960 64164 5016 64166
rect 5040 64164 5096 64166
rect 5120 64164 5176 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4880 63130 4936 63132
rect 4960 63130 5016 63132
rect 5040 63130 5096 63132
rect 5120 63130 5176 63132
rect 4880 63078 4926 63130
rect 4926 63078 4936 63130
rect 4960 63078 4990 63130
rect 4990 63078 5002 63130
rect 5002 63078 5016 63130
rect 5040 63078 5054 63130
rect 5054 63078 5066 63130
rect 5066 63078 5096 63130
rect 5120 63078 5130 63130
rect 5130 63078 5176 63130
rect 4880 63076 4936 63078
rect 4960 63076 5016 63078
rect 5040 63076 5096 63078
rect 5120 63076 5176 63078
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4880 62042 4936 62044
rect 4960 62042 5016 62044
rect 5040 62042 5096 62044
rect 5120 62042 5176 62044
rect 4880 61990 4926 62042
rect 4926 61990 4936 62042
rect 4960 61990 4990 62042
rect 4990 61990 5002 62042
rect 5002 61990 5016 62042
rect 5040 61990 5054 62042
rect 5054 61990 5066 62042
rect 5066 61990 5096 62042
rect 5120 61990 5130 62042
rect 5130 61990 5176 62042
rect 4880 61988 4936 61990
rect 4960 61988 5016 61990
rect 5040 61988 5096 61990
rect 5120 61988 5176 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4880 60954 4936 60956
rect 4960 60954 5016 60956
rect 5040 60954 5096 60956
rect 5120 60954 5176 60956
rect 4880 60902 4926 60954
rect 4926 60902 4936 60954
rect 4960 60902 4990 60954
rect 4990 60902 5002 60954
rect 5002 60902 5016 60954
rect 5040 60902 5054 60954
rect 5054 60902 5066 60954
rect 5066 60902 5096 60954
rect 5120 60902 5130 60954
rect 5130 60902 5176 60954
rect 4880 60900 4936 60902
rect 4960 60900 5016 60902
rect 5040 60900 5096 60902
rect 5120 60900 5176 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4880 59866 4936 59868
rect 4960 59866 5016 59868
rect 5040 59866 5096 59868
rect 5120 59866 5176 59868
rect 4880 59814 4926 59866
rect 4926 59814 4936 59866
rect 4960 59814 4990 59866
rect 4990 59814 5002 59866
rect 5002 59814 5016 59866
rect 5040 59814 5054 59866
rect 5054 59814 5066 59866
rect 5066 59814 5096 59866
rect 5120 59814 5130 59866
rect 5130 59814 5176 59866
rect 4880 59812 4936 59814
rect 4960 59812 5016 59814
rect 5040 59812 5096 59814
rect 5120 59812 5176 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4880 58778 4936 58780
rect 4960 58778 5016 58780
rect 5040 58778 5096 58780
rect 5120 58778 5176 58780
rect 4880 58726 4926 58778
rect 4926 58726 4936 58778
rect 4960 58726 4990 58778
rect 4990 58726 5002 58778
rect 5002 58726 5016 58778
rect 5040 58726 5054 58778
rect 5054 58726 5066 58778
rect 5066 58726 5096 58778
rect 5120 58726 5130 58778
rect 5130 58726 5176 58778
rect 4880 58724 4936 58726
rect 4960 58724 5016 58726
rect 5040 58724 5096 58726
rect 5120 58724 5176 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 1306 44240 1362 44296
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 1306 42880 1362 42936
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 1306 40840 1362 40896
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 1306 40160 1362 40216
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 1214 38120 1270 38176
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1306 37440 1362 37496
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 1306 35400 1362 35456
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1306 15680 1362 15736
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 34940 91962 34996 91964
rect 35020 91962 35076 91964
rect 35100 91962 35156 91964
rect 35180 91962 35236 91964
rect 34940 91910 34986 91962
rect 34986 91910 34996 91962
rect 35020 91910 35050 91962
rect 35050 91910 35062 91962
rect 35062 91910 35076 91962
rect 35100 91910 35114 91962
rect 35114 91910 35126 91962
rect 35126 91910 35156 91962
rect 35180 91910 35190 91962
rect 35190 91910 35236 91962
rect 34940 91908 34996 91910
rect 35020 91908 35076 91910
rect 35100 91908 35156 91910
rect 35180 91908 35236 91910
rect 53194 91976 53250 92012
rect 55586 93916 55588 93936
rect 55588 93916 55640 93936
rect 55640 93916 55642 93936
rect 55586 93880 55642 93916
rect 57978 92812 58034 92848
rect 57978 92792 57980 92812
rect 57980 92792 58032 92812
rect 58032 92792 58034 92812
rect 56598 92520 56654 92576
rect 58438 92792 58494 92848
rect 58714 92132 58770 92168
rect 58714 92112 58716 92132
rect 58716 92112 58768 92132
rect 58768 92112 58770 92132
rect 58162 89936 58218 89992
rect 59266 89800 59322 89856
rect 59818 92656 59874 92712
rect 59450 89936 59506 89992
rect 46846 89664 46902 89720
rect 59358 89664 59414 89720
rect 63498 92948 63554 92984
rect 63498 92928 63500 92948
rect 63500 92928 63552 92948
rect 63552 92928 63554 92948
rect 64878 93200 64934 93256
rect 63498 92520 63554 92576
rect 63774 92520 63830 92576
rect 62854 91024 62910 91080
rect 66320 96858 66376 96860
rect 66400 96858 66456 96860
rect 66480 96858 66536 96860
rect 66560 96858 66616 96860
rect 66320 96806 66366 96858
rect 66366 96806 66376 96858
rect 66400 96806 66430 96858
rect 66430 96806 66442 96858
rect 66442 96806 66456 96858
rect 66480 96806 66494 96858
rect 66494 96806 66506 96858
rect 66506 96806 66536 96858
rect 66560 96806 66570 96858
rect 66570 96806 66616 96858
rect 66320 96804 66376 96806
rect 66400 96804 66456 96806
rect 66480 96804 66536 96806
rect 66560 96804 66616 96806
rect 65660 96314 65716 96316
rect 65740 96314 65796 96316
rect 65820 96314 65876 96316
rect 65900 96314 65956 96316
rect 65660 96262 65706 96314
rect 65706 96262 65716 96314
rect 65740 96262 65770 96314
rect 65770 96262 65782 96314
rect 65782 96262 65796 96314
rect 65820 96262 65834 96314
rect 65834 96262 65846 96314
rect 65846 96262 65876 96314
rect 65900 96262 65910 96314
rect 65910 96262 65956 96314
rect 65660 96260 65716 96262
rect 65740 96260 65796 96262
rect 65820 96260 65876 96262
rect 65900 96260 65956 96262
rect 66320 95770 66376 95772
rect 66400 95770 66456 95772
rect 66480 95770 66536 95772
rect 66560 95770 66616 95772
rect 66320 95718 66366 95770
rect 66366 95718 66376 95770
rect 66400 95718 66430 95770
rect 66430 95718 66442 95770
rect 66442 95718 66456 95770
rect 66480 95718 66494 95770
rect 66494 95718 66506 95770
rect 66506 95718 66536 95770
rect 66560 95718 66570 95770
rect 66570 95718 66616 95770
rect 66320 95716 66376 95718
rect 66400 95716 66456 95718
rect 66480 95716 66536 95718
rect 66560 95716 66616 95718
rect 65660 95226 65716 95228
rect 65740 95226 65796 95228
rect 65820 95226 65876 95228
rect 65900 95226 65956 95228
rect 65660 95174 65706 95226
rect 65706 95174 65716 95226
rect 65740 95174 65770 95226
rect 65770 95174 65782 95226
rect 65782 95174 65796 95226
rect 65820 95174 65834 95226
rect 65834 95174 65846 95226
rect 65846 95174 65876 95226
rect 65900 95174 65910 95226
rect 65910 95174 65956 95226
rect 65660 95172 65716 95174
rect 65740 95172 65796 95174
rect 65820 95172 65876 95174
rect 65900 95172 65956 95174
rect 66320 94682 66376 94684
rect 66400 94682 66456 94684
rect 66480 94682 66536 94684
rect 66560 94682 66616 94684
rect 66320 94630 66366 94682
rect 66366 94630 66376 94682
rect 66400 94630 66430 94682
rect 66430 94630 66442 94682
rect 66442 94630 66456 94682
rect 66480 94630 66494 94682
rect 66494 94630 66506 94682
rect 66506 94630 66536 94682
rect 66560 94630 66570 94682
rect 66570 94630 66616 94682
rect 66320 94628 66376 94630
rect 66400 94628 66456 94630
rect 66480 94628 66536 94630
rect 66560 94628 66616 94630
rect 65660 94138 65716 94140
rect 65740 94138 65796 94140
rect 65820 94138 65876 94140
rect 65900 94138 65956 94140
rect 65660 94086 65706 94138
rect 65706 94086 65716 94138
rect 65740 94086 65770 94138
rect 65770 94086 65782 94138
rect 65782 94086 65796 94138
rect 65820 94086 65834 94138
rect 65834 94086 65846 94138
rect 65846 94086 65876 94138
rect 65900 94086 65910 94138
rect 65910 94086 65956 94138
rect 65660 94084 65716 94086
rect 65740 94084 65796 94086
rect 65820 94084 65876 94086
rect 65900 94084 65956 94086
rect 65890 93780 65892 93800
rect 65892 93780 65944 93800
rect 65944 93780 65946 93800
rect 65890 93744 65946 93780
rect 66320 93594 66376 93596
rect 66400 93594 66456 93596
rect 66480 93594 66536 93596
rect 66560 93594 66616 93596
rect 66320 93542 66366 93594
rect 66366 93542 66376 93594
rect 66400 93542 66430 93594
rect 66430 93542 66442 93594
rect 66442 93542 66456 93594
rect 66480 93542 66494 93594
rect 66494 93542 66506 93594
rect 66506 93542 66536 93594
rect 66560 93542 66570 93594
rect 66570 93542 66616 93594
rect 66320 93540 66376 93542
rect 66400 93540 66456 93542
rect 66480 93540 66536 93542
rect 66560 93540 66616 93542
rect 67270 93764 67326 93800
rect 67270 93744 67272 93764
rect 67272 93744 67324 93764
rect 67324 93744 67326 93764
rect 65660 93050 65716 93052
rect 65740 93050 65796 93052
rect 65820 93050 65876 93052
rect 65900 93050 65956 93052
rect 65660 92998 65706 93050
rect 65706 92998 65716 93050
rect 65740 92998 65770 93050
rect 65770 92998 65782 93050
rect 65782 92998 65796 93050
rect 65820 92998 65834 93050
rect 65834 92998 65846 93050
rect 65846 92998 65876 93050
rect 65900 92998 65910 93050
rect 65910 92998 65956 93050
rect 65660 92996 65716 92998
rect 65740 92996 65796 92998
rect 65820 92996 65876 92998
rect 65900 92996 65956 92998
rect 66320 92506 66376 92508
rect 66400 92506 66456 92508
rect 66480 92506 66536 92508
rect 66560 92506 66616 92508
rect 66320 92454 66366 92506
rect 66366 92454 66376 92506
rect 66400 92454 66430 92506
rect 66430 92454 66442 92506
rect 66442 92454 66456 92506
rect 66480 92454 66494 92506
rect 66494 92454 66506 92506
rect 66506 92454 66536 92506
rect 66560 92454 66570 92506
rect 66570 92454 66616 92506
rect 66320 92452 66376 92454
rect 66400 92452 66456 92454
rect 66480 92452 66536 92454
rect 66560 92452 66616 92454
rect 65660 91962 65716 91964
rect 65740 91962 65796 91964
rect 65820 91962 65876 91964
rect 65900 91962 65956 91964
rect 65660 91910 65706 91962
rect 65706 91910 65716 91962
rect 65740 91910 65770 91962
rect 65770 91910 65782 91962
rect 65782 91910 65796 91962
rect 65820 91910 65834 91962
rect 65834 91910 65846 91962
rect 65846 91910 65876 91962
rect 65900 91910 65910 91962
rect 65910 91910 65956 91962
rect 65660 91908 65716 91910
rect 65740 91908 65796 91910
rect 65820 91908 65876 91910
rect 65900 91908 65956 91910
rect 96380 97402 96436 97404
rect 96460 97402 96516 97404
rect 96540 97402 96596 97404
rect 96620 97402 96676 97404
rect 96380 97350 96426 97402
rect 96426 97350 96436 97402
rect 96460 97350 96490 97402
rect 96490 97350 96502 97402
rect 96502 97350 96516 97402
rect 96540 97350 96554 97402
rect 96554 97350 96566 97402
rect 96566 97350 96596 97402
rect 96620 97350 96630 97402
rect 96630 97350 96676 97402
rect 96380 97348 96436 97350
rect 96460 97348 96516 97350
rect 96540 97348 96596 97350
rect 96620 97348 96676 97350
rect 69202 93200 69258 93256
rect 69202 92520 69258 92576
rect 70490 92520 70546 92576
rect 97040 96858 97096 96860
rect 97120 96858 97176 96860
rect 97200 96858 97256 96860
rect 97280 96858 97336 96860
rect 97040 96806 97086 96858
rect 97086 96806 97096 96858
rect 97120 96806 97150 96858
rect 97150 96806 97162 96858
rect 97162 96806 97176 96858
rect 97200 96806 97214 96858
rect 97214 96806 97226 96858
rect 97226 96806 97256 96858
rect 97280 96806 97290 96858
rect 97290 96806 97336 96858
rect 97040 96804 97096 96806
rect 97120 96804 97176 96806
rect 97200 96804 97256 96806
rect 97280 96804 97336 96806
rect 96380 96314 96436 96316
rect 96460 96314 96516 96316
rect 96540 96314 96596 96316
rect 96620 96314 96676 96316
rect 96380 96262 96426 96314
rect 96426 96262 96436 96314
rect 96460 96262 96490 96314
rect 96490 96262 96502 96314
rect 96502 96262 96516 96314
rect 96540 96262 96554 96314
rect 96554 96262 96566 96314
rect 96566 96262 96596 96314
rect 96620 96262 96630 96314
rect 96630 96262 96676 96314
rect 96380 96260 96436 96262
rect 96460 96260 96516 96262
rect 96540 96260 96596 96262
rect 96620 96260 96676 96262
rect 97040 95770 97096 95772
rect 97120 95770 97176 95772
rect 97200 95770 97256 95772
rect 97280 95770 97336 95772
rect 97040 95718 97086 95770
rect 97086 95718 97096 95770
rect 97120 95718 97150 95770
rect 97150 95718 97162 95770
rect 97162 95718 97176 95770
rect 97200 95718 97214 95770
rect 97214 95718 97226 95770
rect 97226 95718 97256 95770
rect 97280 95718 97290 95770
rect 97290 95718 97336 95770
rect 97040 95716 97096 95718
rect 97120 95716 97176 95718
rect 97200 95716 97256 95718
rect 97280 95716 97336 95718
rect 96380 95226 96436 95228
rect 96460 95226 96516 95228
rect 96540 95226 96596 95228
rect 96620 95226 96676 95228
rect 96380 95174 96426 95226
rect 96426 95174 96436 95226
rect 96460 95174 96490 95226
rect 96490 95174 96502 95226
rect 96502 95174 96516 95226
rect 96540 95174 96554 95226
rect 96554 95174 96566 95226
rect 96566 95174 96596 95226
rect 96620 95174 96630 95226
rect 96630 95174 96676 95226
rect 96380 95172 96436 95174
rect 96460 95172 96516 95174
rect 96540 95172 96596 95174
rect 96620 95172 96676 95174
rect 97040 94682 97096 94684
rect 97120 94682 97176 94684
rect 97200 94682 97256 94684
rect 97280 94682 97336 94684
rect 97040 94630 97086 94682
rect 97086 94630 97096 94682
rect 97120 94630 97150 94682
rect 97150 94630 97162 94682
rect 97162 94630 97176 94682
rect 97200 94630 97214 94682
rect 97214 94630 97226 94682
rect 97226 94630 97256 94682
rect 97280 94630 97290 94682
rect 97290 94630 97336 94682
rect 97040 94628 97096 94630
rect 97120 94628 97176 94630
rect 97200 94628 97256 94630
rect 97280 94628 97336 94630
rect 96380 94138 96436 94140
rect 96460 94138 96516 94140
rect 96540 94138 96596 94140
rect 96620 94138 96676 94140
rect 96380 94086 96426 94138
rect 96426 94086 96436 94138
rect 96460 94086 96490 94138
rect 96490 94086 96502 94138
rect 96502 94086 96516 94138
rect 96540 94086 96554 94138
rect 96554 94086 96566 94138
rect 96566 94086 96596 94138
rect 96620 94086 96630 94138
rect 96630 94086 96676 94138
rect 96380 94084 96436 94086
rect 96460 94084 96516 94086
rect 96540 94084 96596 94086
rect 96620 94084 96676 94086
rect 97040 93594 97096 93596
rect 97120 93594 97176 93596
rect 97200 93594 97256 93596
rect 97280 93594 97336 93596
rect 97040 93542 97086 93594
rect 97086 93542 97096 93594
rect 97120 93542 97150 93594
rect 97150 93542 97162 93594
rect 97162 93542 97176 93594
rect 97200 93542 97214 93594
rect 97214 93542 97226 93594
rect 97226 93542 97256 93594
rect 97280 93542 97290 93594
rect 97290 93542 97336 93594
rect 97040 93540 97096 93542
rect 97120 93540 97176 93542
rect 97200 93540 97256 93542
rect 97280 93540 97336 93542
rect 73250 91024 73306 91080
rect 96380 93050 96436 93052
rect 96460 93050 96516 93052
rect 96540 93050 96596 93052
rect 96620 93050 96676 93052
rect 96380 92998 96426 93050
rect 96426 92998 96436 93050
rect 96460 92998 96490 93050
rect 96490 92998 96502 93050
rect 96502 92998 96516 93050
rect 96540 92998 96554 93050
rect 96554 92998 96566 93050
rect 96566 92998 96596 93050
rect 96620 92998 96630 93050
rect 96630 92998 96676 93050
rect 96380 92996 96436 92998
rect 96460 92996 96516 92998
rect 96540 92996 96596 92998
rect 96620 92996 96676 92998
rect 74170 91024 74226 91080
rect 97040 92506 97096 92508
rect 97120 92506 97176 92508
rect 97200 92506 97256 92508
rect 97280 92506 97336 92508
rect 97040 92454 97086 92506
rect 97086 92454 97096 92506
rect 97120 92454 97150 92506
rect 97150 92454 97162 92506
rect 97162 92454 97176 92506
rect 97200 92454 97214 92506
rect 97214 92454 97226 92506
rect 97226 92454 97256 92506
rect 97280 92454 97290 92506
rect 97290 92454 97336 92506
rect 97040 92452 97096 92454
rect 97120 92452 97176 92454
rect 97200 92452 97256 92454
rect 97280 92452 97336 92454
rect 96380 91962 96436 91964
rect 96460 91962 96516 91964
rect 96540 91962 96596 91964
rect 96620 91962 96676 91964
rect 96380 91910 96426 91962
rect 96426 91910 96436 91962
rect 96460 91910 96490 91962
rect 96490 91910 96502 91962
rect 96502 91910 96516 91962
rect 96540 91910 96554 91962
rect 96554 91910 96566 91962
rect 96566 91910 96596 91962
rect 96620 91910 96630 91962
rect 96630 91910 96676 91962
rect 96380 91908 96436 91910
rect 96460 91908 96516 91910
rect 96540 91908 96596 91910
rect 96620 91908 96676 91910
rect 100022 91160 100078 91216
rect 65246 89664 65302 89720
rect 66810 89664 66866 89720
rect 67546 89664 67602 89720
rect 71870 89664 71926 89720
rect 73710 89664 73766 89720
rect 75918 89664 75974 89720
rect 89442 89664 89498 89720
rect 60554 89528 60610 89584
rect 106922 89528 106978 89584
rect 106186 86442 106242 86498
rect 113656 92506 113712 92508
rect 113736 92506 113792 92508
rect 113816 92506 113872 92508
rect 113896 92506 113952 92508
rect 113656 92454 113702 92506
rect 113702 92454 113712 92506
rect 113736 92454 113766 92506
rect 113766 92454 113778 92506
rect 113778 92454 113792 92506
rect 113816 92454 113830 92506
rect 113830 92454 113842 92506
rect 113842 92454 113872 92506
rect 113896 92454 113906 92506
rect 113906 92454 113952 92506
rect 113656 92452 113712 92454
rect 113736 92452 113792 92454
rect 113816 92452 113872 92454
rect 113896 92452 113952 92454
rect 112920 91962 112976 91964
rect 113000 91962 113056 91964
rect 113080 91962 113136 91964
rect 113160 91962 113216 91964
rect 112920 91910 112966 91962
rect 112966 91910 112976 91962
rect 113000 91910 113030 91962
rect 113030 91910 113042 91962
rect 113042 91910 113056 91962
rect 113080 91910 113094 91962
rect 113094 91910 113106 91962
rect 113106 91910 113136 91962
rect 113160 91910 113170 91962
rect 113170 91910 113216 91962
rect 112920 91908 112976 91910
rect 113000 91908 113056 91910
rect 113080 91908 113136 91910
rect 113160 91908 113216 91910
rect 113656 91418 113712 91420
rect 113736 91418 113792 91420
rect 113816 91418 113872 91420
rect 113896 91418 113952 91420
rect 113656 91366 113702 91418
rect 113702 91366 113712 91418
rect 113736 91366 113766 91418
rect 113766 91366 113778 91418
rect 113778 91366 113792 91418
rect 113816 91366 113830 91418
rect 113830 91366 113842 91418
rect 113842 91366 113872 91418
rect 113896 91366 113906 91418
rect 113906 91366 113952 91418
rect 113656 91364 113712 91366
rect 113736 91364 113792 91366
rect 113816 91364 113872 91366
rect 113896 91364 113952 91366
rect 112920 90874 112976 90876
rect 113000 90874 113056 90876
rect 113080 90874 113136 90876
rect 113160 90874 113216 90876
rect 112920 90822 112966 90874
rect 112966 90822 112976 90874
rect 113000 90822 113030 90874
rect 113030 90822 113042 90874
rect 113042 90822 113056 90874
rect 113080 90822 113094 90874
rect 113094 90822 113106 90874
rect 113106 90822 113136 90874
rect 113160 90822 113170 90874
rect 113170 90822 113216 90874
rect 112920 90820 112976 90822
rect 113000 90820 113056 90822
rect 113080 90820 113136 90822
rect 113160 90820 113216 90822
rect 113656 90330 113712 90332
rect 113736 90330 113792 90332
rect 113816 90330 113872 90332
rect 113896 90330 113952 90332
rect 113656 90278 113702 90330
rect 113702 90278 113712 90330
rect 113736 90278 113766 90330
rect 113766 90278 113778 90330
rect 113778 90278 113792 90330
rect 113816 90278 113830 90330
rect 113830 90278 113842 90330
rect 113842 90278 113872 90330
rect 113896 90278 113906 90330
rect 113906 90278 113952 90330
rect 113656 90276 113712 90278
rect 113736 90276 113792 90278
rect 113816 90276 113872 90278
rect 113896 90276 113952 90278
rect 112920 89786 112976 89788
rect 113000 89786 113056 89788
rect 113080 89786 113136 89788
rect 113160 89786 113216 89788
rect 112920 89734 112966 89786
rect 112966 89734 112976 89786
rect 113000 89734 113030 89786
rect 113030 89734 113042 89786
rect 113042 89734 113056 89786
rect 113080 89734 113094 89786
rect 113094 89734 113106 89786
rect 113106 89734 113136 89786
rect 113160 89734 113170 89786
rect 113170 89734 113216 89786
rect 112920 89732 112976 89734
rect 113000 89732 113056 89734
rect 113080 89732 113136 89734
rect 113160 89732 113216 89734
rect 113656 89242 113712 89244
rect 113736 89242 113792 89244
rect 113816 89242 113872 89244
rect 113896 89242 113952 89244
rect 113656 89190 113702 89242
rect 113702 89190 113712 89242
rect 113736 89190 113766 89242
rect 113766 89190 113778 89242
rect 113778 89190 113792 89242
rect 113816 89190 113830 89242
rect 113830 89190 113842 89242
rect 113842 89190 113872 89242
rect 113896 89190 113906 89242
rect 113906 89190 113952 89242
rect 113656 89188 113712 89190
rect 113736 89188 113792 89190
rect 113816 89188 113872 89190
rect 113896 89188 113952 89190
rect 112920 88698 112976 88700
rect 113000 88698 113056 88700
rect 113080 88698 113136 88700
rect 113160 88698 113216 88700
rect 112920 88646 112966 88698
rect 112966 88646 112976 88698
rect 113000 88646 113030 88698
rect 113030 88646 113042 88698
rect 113042 88646 113056 88698
rect 113080 88646 113094 88698
rect 113094 88646 113106 88698
rect 113106 88646 113136 88698
rect 113160 88646 113170 88698
rect 113170 88646 113216 88698
rect 112920 88644 112976 88646
rect 113000 88644 113056 88646
rect 113080 88644 113136 88646
rect 113160 88644 113216 88646
rect 113656 88154 113712 88156
rect 113736 88154 113792 88156
rect 113816 88154 113872 88156
rect 113896 88154 113952 88156
rect 113656 88102 113702 88154
rect 113702 88102 113712 88154
rect 113736 88102 113766 88154
rect 113766 88102 113778 88154
rect 113778 88102 113792 88154
rect 113816 88102 113830 88154
rect 113830 88102 113842 88154
rect 113842 88102 113872 88154
rect 113896 88102 113906 88154
rect 113906 88102 113952 88154
rect 113656 88100 113712 88102
rect 113736 88100 113792 88102
rect 113816 88100 113872 88102
rect 113896 88100 113952 88102
rect 112920 87610 112976 87612
rect 113000 87610 113056 87612
rect 113080 87610 113136 87612
rect 113160 87610 113216 87612
rect 112920 87558 112966 87610
rect 112966 87558 112976 87610
rect 113000 87558 113030 87610
rect 113030 87558 113042 87610
rect 113042 87558 113056 87610
rect 113080 87558 113094 87610
rect 113094 87558 113106 87610
rect 113106 87558 113136 87610
rect 113160 87558 113170 87610
rect 113170 87558 113216 87610
rect 112920 87556 112976 87558
rect 113000 87556 113056 87558
rect 113080 87556 113136 87558
rect 113160 87556 113216 87558
rect 113656 87066 113712 87068
rect 113736 87066 113792 87068
rect 113816 87066 113872 87068
rect 113896 87066 113952 87068
rect 113656 87014 113702 87066
rect 113702 87014 113712 87066
rect 113736 87014 113766 87066
rect 113766 87014 113778 87066
rect 113778 87014 113792 87066
rect 113816 87014 113830 87066
rect 113830 87014 113842 87066
rect 113842 87014 113872 87066
rect 113896 87014 113906 87066
rect 113906 87014 113952 87066
rect 113656 87012 113712 87014
rect 113736 87012 113792 87014
rect 113816 87012 113872 87014
rect 113896 87012 113952 87014
rect 112920 86522 112976 86524
rect 113000 86522 113056 86524
rect 113080 86522 113136 86524
rect 113160 86522 113216 86524
rect 112920 86470 112966 86522
rect 112966 86470 112976 86522
rect 113000 86470 113030 86522
rect 113030 86470 113042 86522
rect 113042 86470 113056 86522
rect 113080 86470 113094 86522
rect 113094 86470 113106 86522
rect 113106 86470 113136 86522
rect 113160 86470 113170 86522
rect 113170 86470 113216 86522
rect 112920 86468 112976 86470
rect 113000 86468 113056 86470
rect 113080 86468 113136 86470
rect 113160 86468 113216 86470
rect 113656 85978 113712 85980
rect 113736 85978 113792 85980
rect 113816 85978 113872 85980
rect 113896 85978 113952 85980
rect 113656 85926 113702 85978
rect 113702 85926 113712 85978
rect 113736 85926 113766 85978
rect 113766 85926 113778 85978
rect 113778 85926 113792 85978
rect 113816 85926 113830 85978
rect 113830 85926 113842 85978
rect 113842 85926 113872 85978
rect 113896 85926 113906 85978
rect 113906 85926 113952 85978
rect 113656 85924 113712 85926
rect 113736 85924 113792 85926
rect 113816 85924 113872 85926
rect 113896 85924 113952 85926
rect 112920 85434 112976 85436
rect 113000 85434 113056 85436
rect 113080 85434 113136 85436
rect 113160 85434 113216 85436
rect 112920 85382 112966 85434
rect 112966 85382 112976 85434
rect 113000 85382 113030 85434
rect 113030 85382 113042 85434
rect 113042 85382 113056 85434
rect 113080 85382 113094 85434
rect 113094 85382 113106 85434
rect 113106 85382 113136 85434
rect 113160 85382 113170 85434
rect 113170 85382 113216 85434
rect 112920 85380 112976 85382
rect 113000 85380 113056 85382
rect 113080 85380 113136 85382
rect 113160 85380 113216 85382
rect 113656 84890 113712 84892
rect 113736 84890 113792 84892
rect 113816 84890 113872 84892
rect 113896 84890 113952 84892
rect 113656 84838 113702 84890
rect 113702 84838 113712 84890
rect 113736 84838 113766 84890
rect 113766 84838 113778 84890
rect 113778 84838 113792 84890
rect 113816 84838 113830 84890
rect 113830 84838 113842 84890
rect 113842 84838 113872 84890
rect 113896 84838 113906 84890
rect 113906 84838 113952 84890
rect 113656 84836 113712 84838
rect 113736 84836 113792 84838
rect 113816 84836 113872 84838
rect 113896 84836 113952 84838
rect 112920 84346 112976 84348
rect 113000 84346 113056 84348
rect 113080 84346 113136 84348
rect 113160 84346 113216 84348
rect 112920 84294 112966 84346
rect 112966 84294 112976 84346
rect 113000 84294 113030 84346
rect 113030 84294 113042 84346
rect 113042 84294 113056 84346
rect 113080 84294 113094 84346
rect 113094 84294 113106 84346
rect 113106 84294 113136 84346
rect 113160 84294 113170 84346
rect 113170 84294 113216 84346
rect 112920 84292 112976 84294
rect 113000 84292 113056 84294
rect 113080 84292 113136 84294
rect 113160 84292 113216 84294
rect 113656 83802 113712 83804
rect 113736 83802 113792 83804
rect 113816 83802 113872 83804
rect 113896 83802 113952 83804
rect 113656 83750 113702 83802
rect 113702 83750 113712 83802
rect 113736 83750 113766 83802
rect 113766 83750 113778 83802
rect 113778 83750 113792 83802
rect 113816 83750 113830 83802
rect 113830 83750 113842 83802
rect 113842 83750 113872 83802
rect 113896 83750 113906 83802
rect 113906 83750 113952 83802
rect 113656 83748 113712 83750
rect 113736 83748 113792 83750
rect 113816 83748 113872 83750
rect 113896 83748 113952 83750
rect 112920 83258 112976 83260
rect 113000 83258 113056 83260
rect 113080 83258 113136 83260
rect 113160 83258 113216 83260
rect 112920 83206 112966 83258
rect 112966 83206 112976 83258
rect 113000 83206 113030 83258
rect 113030 83206 113042 83258
rect 113042 83206 113056 83258
rect 113080 83206 113094 83258
rect 113094 83206 113106 83258
rect 113106 83206 113136 83258
rect 113160 83206 113170 83258
rect 113170 83206 113216 83258
rect 112920 83204 112976 83206
rect 113000 83204 113056 83206
rect 113080 83204 113136 83206
rect 113160 83204 113216 83206
rect 113656 82714 113712 82716
rect 113736 82714 113792 82716
rect 113816 82714 113872 82716
rect 113896 82714 113952 82716
rect 113656 82662 113702 82714
rect 113702 82662 113712 82714
rect 113736 82662 113766 82714
rect 113766 82662 113778 82714
rect 113778 82662 113792 82714
rect 113816 82662 113830 82714
rect 113830 82662 113842 82714
rect 113842 82662 113872 82714
rect 113896 82662 113906 82714
rect 113906 82662 113952 82714
rect 113656 82660 113712 82662
rect 113736 82660 113792 82662
rect 113816 82660 113872 82662
rect 113896 82660 113952 82662
rect 112920 82170 112976 82172
rect 113000 82170 113056 82172
rect 113080 82170 113136 82172
rect 113160 82170 113216 82172
rect 112920 82118 112966 82170
rect 112966 82118 112976 82170
rect 113000 82118 113030 82170
rect 113030 82118 113042 82170
rect 113042 82118 113056 82170
rect 113080 82118 113094 82170
rect 113094 82118 113106 82170
rect 113106 82118 113136 82170
rect 113160 82118 113170 82170
rect 113170 82118 113216 82170
rect 112920 82116 112976 82118
rect 113000 82116 113056 82118
rect 113080 82116 113136 82118
rect 113160 82116 113216 82118
rect 113656 81626 113712 81628
rect 113736 81626 113792 81628
rect 113816 81626 113872 81628
rect 113896 81626 113952 81628
rect 113656 81574 113702 81626
rect 113702 81574 113712 81626
rect 113736 81574 113766 81626
rect 113766 81574 113778 81626
rect 113778 81574 113792 81626
rect 113816 81574 113830 81626
rect 113830 81574 113842 81626
rect 113842 81574 113872 81626
rect 113896 81574 113906 81626
rect 113906 81574 113952 81626
rect 113656 81572 113712 81574
rect 113736 81572 113792 81574
rect 113816 81572 113872 81574
rect 113896 81572 113952 81574
rect 112920 81082 112976 81084
rect 113000 81082 113056 81084
rect 113080 81082 113136 81084
rect 113160 81082 113216 81084
rect 112920 81030 112966 81082
rect 112966 81030 112976 81082
rect 113000 81030 113030 81082
rect 113030 81030 113042 81082
rect 113042 81030 113056 81082
rect 113080 81030 113094 81082
rect 113094 81030 113106 81082
rect 113106 81030 113136 81082
rect 113160 81030 113170 81082
rect 113170 81030 113216 81082
rect 112920 81028 112976 81030
rect 113000 81028 113056 81030
rect 113080 81028 113136 81030
rect 113160 81028 113216 81030
rect 113656 80538 113712 80540
rect 113736 80538 113792 80540
rect 113816 80538 113872 80540
rect 113896 80538 113952 80540
rect 113656 80486 113702 80538
rect 113702 80486 113712 80538
rect 113736 80486 113766 80538
rect 113766 80486 113778 80538
rect 113778 80486 113792 80538
rect 113816 80486 113830 80538
rect 113830 80486 113842 80538
rect 113842 80486 113872 80538
rect 113896 80486 113906 80538
rect 113906 80486 113952 80538
rect 113656 80484 113712 80486
rect 113736 80484 113792 80486
rect 113816 80484 113872 80486
rect 113896 80484 113952 80486
rect 112920 79994 112976 79996
rect 113000 79994 113056 79996
rect 113080 79994 113136 79996
rect 113160 79994 113216 79996
rect 112920 79942 112966 79994
rect 112966 79942 112976 79994
rect 113000 79942 113030 79994
rect 113030 79942 113042 79994
rect 113042 79942 113056 79994
rect 113080 79942 113094 79994
rect 113094 79942 113106 79994
rect 113106 79942 113136 79994
rect 113160 79942 113170 79994
rect 113170 79942 113216 79994
rect 112920 79940 112976 79942
rect 113000 79940 113056 79942
rect 113080 79940 113136 79942
rect 113160 79940 113216 79942
rect 113656 79450 113712 79452
rect 113736 79450 113792 79452
rect 113816 79450 113872 79452
rect 113896 79450 113952 79452
rect 113656 79398 113702 79450
rect 113702 79398 113712 79450
rect 113736 79398 113766 79450
rect 113766 79398 113778 79450
rect 113778 79398 113792 79450
rect 113816 79398 113830 79450
rect 113830 79398 113842 79450
rect 113842 79398 113872 79450
rect 113896 79398 113906 79450
rect 113906 79398 113952 79450
rect 113656 79396 113712 79398
rect 113736 79396 113792 79398
rect 113816 79396 113872 79398
rect 113896 79396 113952 79398
rect 112920 78906 112976 78908
rect 113000 78906 113056 78908
rect 113080 78906 113136 78908
rect 113160 78906 113216 78908
rect 112920 78854 112966 78906
rect 112966 78854 112976 78906
rect 113000 78854 113030 78906
rect 113030 78854 113042 78906
rect 113042 78854 113056 78906
rect 113080 78854 113094 78906
rect 113094 78854 113106 78906
rect 113106 78854 113136 78906
rect 113160 78854 113170 78906
rect 113170 78854 113216 78906
rect 112920 78852 112976 78854
rect 113000 78852 113056 78854
rect 113080 78852 113136 78854
rect 113160 78852 113216 78854
rect 113656 78362 113712 78364
rect 113736 78362 113792 78364
rect 113816 78362 113872 78364
rect 113896 78362 113952 78364
rect 113656 78310 113702 78362
rect 113702 78310 113712 78362
rect 113736 78310 113766 78362
rect 113766 78310 113778 78362
rect 113778 78310 113792 78362
rect 113816 78310 113830 78362
rect 113830 78310 113842 78362
rect 113842 78310 113872 78362
rect 113896 78310 113906 78362
rect 113906 78310 113952 78362
rect 113656 78308 113712 78310
rect 113736 78308 113792 78310
rect 113816 78308 113872 78310
rect 113896 78308 113952 78310
rect 112920 77818 112976 77820
rect 113000 77818 113056 77820
rect 113080 77818 113136 77820
rect 113160 77818 113216 77820
rect 112920 77766 112966 77818
rect 112966 77766 112976 77818
rect 113000 77766 113030 77818
rect 113030 77766 113042 77818
rect 113042 77766 113056 77818
rect 113080 77766 113094 77818
rect 113094 77766 113106 77818
rect 113106 77766 113136 77818
rect 113160 77766 113170 77818
rect 113170 77766 113216 77818
rect 112920 77764 112976 77766
rect 113000 77764 113056 77766
rect 113080 77764 113136 77766
rect 113160 77764 113216 77766
rect 113656 77274 113712 77276
rect 113736 77274 113792 77276
rect 113816 77274 113872 77276
rect 113896 77274 113952 77276
rect 113656 77222 113702 77274
rect 113702 77222 113712 77274
rect 113736 77222 113766 77274
rect 113766 77222 113778 77274
rect 113778 77222 113792 77274
rect 113816 77222 113830 77274
rect 113830 77222 113842 77274
rect 113842 77222 113872 77274
rect 113896 77222 113906 77274
rect 113906 77222 113952 77274
rect 113656 77220 113712 77222
rect 113736 77220 113792 77222
rect 113816 77220 113872 77222
rect 113896 77220 113952 77222
rect 112920 76730 112976 76732
rect 113000 76730 113056 76732
rect 113080 76730 113136 76732
rect 113160 76730 113216 76732
rect 112920 76678 112966 76730
rect 112966 76678 112976 76730
rect 113000 76678 113030 76730
rect 113030 76678 113042 76730
rect 113042 76678 113056 76730
rect 113080 76678 113094 76730
rect 113094 76678 113106 76730
rect 113106 76678 113136 76730
rect 113160 76678 113170 76730
rect 113170 76678 113216 76730
rect 112920 76676 112976 76678
rect 113000 76676 113056 76678
rect 113080 76676 113136 76678
rect 113160 76676 113216 76678
rect 113656 76186 113712 76188
rect 113736 76186 113792 76188
rect 113816 76186 113872 76188
rect 113896 76186 113952 76188
rect 113656 76134 113702 76186
rect 113702 76134 113712 76186
rect 113736 76134 113766 76186
rect 113766 76134 113778 76186
rect 113778 76134 113792 76186
rect 113816 76134 113830 76186
rect 113830 76134 113842 76186
rect 113842 76134 113872 76186
rect 113896 76134 113906 76186
rect 113906 76134 113952 76186
rect 113656 76132 113712 76134
rect 113736 76132 113792 76134
rect 113816 76132 113872 76134
rect 113896 76132 113952 76134
rect 112920 75642 112976 75644
rect 113000 75642 113056 75644
rect 113080 75642 113136 75644
rect 113160 75642 113216 75644
rect 112920 75590 112966 75642
rect 112966 75590 112976 75642
rect 113000 75590 113030 75642
rect 113030 75590 113042 75642
rect 113042 75590 113056 75642
rect 113080 75590 113094 75642
rect 113094 75590 113106 75642
rect 113106 75590 113136 75642
rect 113160 75590 113170 75642
rect 113170 75590 113216 75642
rect 112920 75588 112976 75590
rect 113000 75588 113056 75590
rect 113080 75588 113136 75590
rect 113160 75588 113216 75590
rect 113656 75098 113712 75100
rect 113736 75098 113792 75100
rect 113816 75098 113872 75100
rect 113896 75098 113952 75100
rect 113656 75046 113702 75098
rect 113702 75046 113712 75098
rect 113736 75046 113766 75098
rect 113766 75046 113778 75098
rect 113778 75046 113792 75098
rect 113816 75046 113830 75098
rect 113830 75046 113842 75098
rect 113842 75046 113872 75098
rect 113896 75046 113906 75098
rect 113906 75046 113952 75098
rect 113656 75044 113712 75046
rect 113736 75044 113792 75046
rect 113816 75044 113872 75046
rect 113896 75044 113952 75046
rect 112920 74554 112976 74556
rect 113000 74554 113056 74556
rect 113080 74554 113136 74556
rect 113160 74554 113216 74556
rect 112920 74502 112966 74554
rect 112966 74502 112976 74554
rect 113000 74502 113030 74554
rect 113030 74502 113042 74554
rect 113042 74502 113056 74554
rect 113080 74502 113094 74554
rect 113094 74502 113106 74554
rect 113106 74502 113136 74554
rect 113160 74502 113170 74554
rect 113170 74502 113216 74554
rect 112920 74500 112976 74502
rect 113000 74500 113056 74502
rect 113080 74500 113136 74502
rect 113160 74500 113216 74502
rect 113656 74010 113712 74012
rect 113736 74010 113792 74012
rect 113816 74010 113872 74012
rect 113896 74010 113952 74012
rect 113656 73958 113702 74010
rect 113702 73958 113712 74010
rect 113736 73958 113766 74010
rect 113766 73958 113778 74010
rect 113778 73958 113792 74010
rect 113816 73958 113830 74010
rect 113830 73958 113842 74010
rect 113842 73958 113872 74010
rect 113896 73958 113906 74010
rect 113906 73958 113952 74010
rect 113656 73956 113712 73958
rect 113736 73956 113792 73958
rect 113816 73956 113872 73958
rect 113896 73956 113952 73958
rect 112920 73466 112976 73468
rect 113000 73466 113056 73468
rect 113080 73466 113136 73468
rect 113160 73466 113216 73468
rect 112920 73414 112966 73466
rect 112966 73414 112976 73466
rect 113000 73414 113030 73466
rect 113030 73414 113042 73466
rect 113042 73414 113056 73466
rect 113080 73414 113094 73466
rect 113094 73414 113106 73466
rect 113106 73414 113136 73466
rect 113160 73414 113170 73466
rect 113170 73414 113216 73466
rect 112920 73412 112976 73414
rect 113000 73412 113056 73414
rect 113080 73412 113136 73414
rect 113160 73412 113216 73414
rect 113656 72922 113712 72924
rect 113736 72922 113792 72924
rect 113816 72922 113872 72924
rect 113896 72922 113952 72924
rect 113656 72870 113702 72922
rect 113702 72870 113712 72922
rect 113736 72870 113766 72922
rect 113766 72870 113778 72922
rect 113778 72870 113792 72922
rect 113816 72870 113830 72922
rect 113830 72870 113842 72922
rect 113842 72870 113872 72922
rect 113896 72870 113906 72922
rect 113906 72870 113952 72922
rect 113656 72868 113712 72870
rect 113736 72868 113792 72870
rect 113816 72868 113872 72870
rect 113896 72868 113952 72870
rect 112920 72378 112976 72380
rect 113000 72378 113056 72380
rect 113080 72378 113136 72380
rect 113160 72378 113216 72380
rect 112920 72326 112966 72378
rect 112966 72326 112976 72378
rect 113000 72326 113030 72378
rect 113030 72326 113042 72378
rect 113042 72326 113056 72378
rect 113080 72326 113094 72378
rect 113094 72326 113106 72378
rect 113106 72326 113136 72378
rect 113160 72326 113170 72378
rect 113170 72326 113216 72378
rect 112920 72324 112976 72326
rect 113000 72324 113056 72326
rect 113080 72324 113136 72326
rect 113160 72324 113216 72326
rect 113656 71834 113712 71836
rect 113736 71834 113792 71836
rect 113816 71834 113872 71836
rect 113896 71834 113952 71836
rect 113656 71782 113702 71834
rect 113702 71782 113712 71834
rect 113736 71782 113766 71834
rect 113766 71782 113778 71834
rect 113778 71782 113792 71834
rect 113816 71782 113830 71834
rect 113830 71782 113842 71834
rect 113842 71782 113872 71834
rect 113896 71782 113906 71834
rect 113906 71782 113952 71834
rect 113656 71780 113712 71782
rect 113736 71780 113792 71782
rect 113816 71780 113872 71782
rect 113896 71780 113952 71782
rect 112920 71290 112976 71292
rect 113000 71290 113056 71292
rect 113080 71290 113136 71292
rect 113160 71290 113216 71292
rect 112920 71238 112966 71290
rect 112966 71238 112976 71290
rect 113000 71238 113030 71290
rect 113030 71238 113042 71290
rect 113042 71238 113056 71290
rect 113080 71238 113094 71290
rect 113094 71238 113106 71290
rect 113106 71238 113136 71290
rect 113160 71238 113170 71290
rect 113170 71238 113216 71290
rect 112920 71236 112976 71238
rect 113000 71236 113056 71238
rect 113080 71236 113136 71238
rect 113160 71236 113216 71238
rect 113656 70746 113712 70748
rect 113736 70746 113792 70748
rect 113816 70746 113872 70748
rect 113896 70746 113952 70748
rect 113656 70694 113702 70746
rect 113702 70694 113712 70746
rect 113736 70694 113766 70746
rect 113766 70694 113778 70746
rect 113778 70694 113792 70746
rect 113816 70694 113830 70746
rect 113830 70694 113842 70746
rect 113842 70694 113872 70746
rect 113896 70694 113906 70746
rect 113906 70694 113952 70746
rect 113656 70692 113712 70694
rect 113736 70692 113792 70694
rect 113816 70692 113872 70694
rect 113896 70692 113952 70694
rect 112920 70202 112976 70204
rect 113000 70202 113056 70204
rect 113080 70202 113136 70204
rect 113160 70202 113216 70204
rect 112920 70150 112966 70202
rect 112966 70150 112976 70202
rect 113000 70150 113030 70202
rect 113030 70150 113042 70202
rect 113042 70150 113056 70202
rect 113080 70150 113094 70202
rect 113094 70150 113106 70202
rect 113106 70150 113136 70202
rect 113160 70150 113170 70202
rect 113170 70150 113216 70202
rect 112920 70148 112976 70150
rect 113000 70148 113056 70150
rect 113080 70148 113136 70150
rect 113160 70148 113216 70150
rect 113656 69658 113712 69660
rect 113736 69658 113792 69660
rect 113816 69658 113872 69660
rect 113896 69658 113952 69660
rect 113656 69606 113702 69658
rect 113702 69606 113712 69658
rect 113736 69606 113766 69658
rect 113766 69606 113778 69658
rect 113778 69606 113792 69658
rect 113816 69606 113830 69658
rect 113830 69606 113842 69658
rect 113842 69606 113872 69658
rect 113896 69606 113906 69658
rect 113906 69606 113952 69658
rect 113656 69604 113712 69606
rect 113736 69604 113792 69606
rect 113816 69604 113872 69606
rect 113896 69604 113952 69606
rect 112920 69114 112976 69116
rect 113000 69114 113056 69116
rect 113080 69114 113136 69116
rect 113160 69114 113216 69116
rect 112920 69062 112966 69114
rect 112966 69062 112976 69114
rect 113000 69062 113030 69114
rect 113030 69062 113042 69114
rect 113042 69062 113056 69114
rect 113080 69062 113094 69114
rect 113094 69062 113106 69114
rect 113106 69062 113136 69114
rect 113160 69062 113170 69114
rect 113170 69062 113216 69114
rect 112920 69060 112976 69062
rect 113000 69060 113056 69062
rect 113080 69060 113136 69062
rect 113160 69060 113216 69062
rect 113656 68570 113712 68572
rect 113736 68570 113792 68572
rect 113816 68570 113872 68572
rect 113896 68570 113952 68572
rect 113656 68518 113702 68570
rect 113702 68518 113712 68570
rect 113736 68518 113766 68570
rect 113766 68518 113778 68570
rect 113778 68518 113792 68570
rect 113816 68518 113830 68570
rect 113830 68518 113842 68570
rect 113842 68518 113872 68570
rect 113896 68518 113906 68570
rect 113906 68518 113952 68570
rect 113656 68516 113712 68518
rect 113736 68516 113792 68518
rect 113816 68516 113872 68518
rect 113896 68516 113952 68518
rect 112920 68026 112976 68028
rect 113000 68026 113056 68028
rect 113080 68026 113136 68028
rect 113160 68026 113216 68028
rect 112920 67974 112966 68026
rect 112966 67974 112976 68026
rect 113000 67974 113030 68026
rect 113030 67974 113042 68026
rect 113042 67974 113056 68026
rect 113080 67974 113094 68026
rect 113094 67974 113106 68026
rect 113106 67974 113136 68026
rect 113160 67974 113170 68026
rect 113170 67974 113216 68026
rect 112920 67972 112976 67974
rect 113000 67972 113056 67974
rect 113080 67972 113136 67974
rect 113160 67972 113216 67974
rect 113656 67482 113712 67484
rect 113736 67482 113792 67484
rect 113816 67482 113872 67484
rect 113896 67482 113952 67484
rect 113656 67430 113702 67482
rect 113702 67430 113712 67482
rect 113736 67430 113766 67482
rect 113766 67430 113778 67482
rect 113778 67430 113792 67482
rect 113816 67430 113830 67482
rect 113830 67430 113842 67482
rect 113842 67430 113872 67482
rect 113896 67430 113906 67482
rect 113906 67430 113952 67482
rect 113656 67428 113712 67430
rect 113736 67428 113792 67430
rect 113816 67428 113872 67430
rect 113896 67428 113952 67430
rect 112920 66938 112976 66940
rect 113000 66938 113056 66940
rect 113080 66938 113136 66940
rect 113160 66938 113216 66940
rect 112920 66886 112966 66938
rect 112966 66886 112976 66938
rect 113000 66886 113030 66938
rect 113030 66886 113042 66938
rect 113042 66886 113056 66938
rect 113080 66886 113094 66938
rect 113094 66886 113106 66938
rect 113106 66886 113136 66938
rect 113160 66886 113170 66938
rect 113170 66886 113216 66938
rect 112920 66884 112976 66886
rect 113000 66884 113056 66886
rect 113080 66884 113136 66886
rect 113160 66884 113216 66886
rect 113656 66394 113712 66396
rect 113736 66394 113792 66396
rect 113816 66394 113872 66396
rect 113896 66394 113952 66396
rect 113656 66342 113702 66394
rect 113702 66342 113712 66394
rect 113736 66342 113766 66394
rect 113766 66342 113778 66394
rect 113778 66342 113792 66394
rect 113816 66342 113830 66394
rect 113830 66342 113842 66394
rect 113842 66342 113872 66394
rect 113896 66342 113906 66394
rect 113906 66342 113952 66394
rect 113656 66340 113712 66342
rect 113736 66340 113792 66342
rect 113816 66340 113872 66342
rect 113896 66340 113952 66342
rect 112920 65850 112976 65852
rect 113000 65850 113056 65852
rect 113080 65850 113136 65852
rect 113160 65850 113216 65852
rect 112920 65798 112966 65850
rect 112966 65798 112976 65850
rect 113000 65798 113030 65850
rect 113030 65798 113042 65850
rect 113042 65798 113056 65850
rect 113080 65798 113094 65850
rect 113094 65798 113106 65850
rect 113106 65798 113136 65850
rect 113160 65798 113170 65850
rect 113170 65798 113216 65850
rect 112920 65796 112976 65798
rect 113000 65796 113056 65798
rect 113080 65796 113136 65798
rect 113160 65796 113216 65798
rect 113656 65306 113712 65308
rect 113736 65306 113792 65308
rect 113816 65306 113872 65308
rect 113896 65306 113952 65308
rect 113656 65254 113702 65306
rect 113702 65254 113712 65306
rect 113736 65254 113766 65306
rect 113766 65254 113778 65306
rect 113778 65254 113792 65306
rect 113816 65254 113830 65306
rect 113830 65254 113842 65306
rect 113842 65254 113872 65306
rect 113896 65254 113906 65306
rect 113906 65254 113952 65306
rect 113656 65252 113712 65254
rect 113736 65252 113792 65254
rect 113816 65252 113872 65254
rect 113896 65252 113952 65254
rect 112920 64762 112976 64764
rect 113000 64762 113056 64764
rect 113080 64762 113136 64764
rect 113160 64762 113216 64764
rect 112920 64710 112966 64762
rect 112966 64710 112976 64762
rect 113000 64710 113030 64762
rect 113030 64710 113042 64762
rect 113042 64710 113056 64762
rect 113080 64710 113094 64762
rect 113094 64710 113106 64762
rect 113106 64710 113136 64762
rect 113160 64710 113170 64762
rect 113170 64710 113216 64762
rect 112920 64708 112976 64710
rect 113000 64708 113056 64710
rect 113080 64708 113136 64710
rect 113160 64708 113216 64710
rect 113656 64218 113712 64220
rect 113736 64218 113792 64220
rect 113816 64218 113872 64220
rect 113896 64218 113952 64220
rect 113656 64166 113702 64218
rect 113702 64166 113712 64218
rect 113736 64166 113766 64218
rect 113766 64166 113778 64218
rect 113778 64166 113792 64218
rect 113816 64166 113830 64218
rect 113830 64166 113842 64218
rect 113842 64166 113872 64218
rect 113896 64166 113906 64218
rect 113906 64166 113952 64218
rect 113656 64164 113712 64166
rect 113736 64164 113792 64166
rect 113816 64164 113872 64166
rect 113896 64164 113952 64166
rect 112920 63674 112976 63676
rect 113000 63674 113056 63676
rect 113080 63674 113136 63676
rect 113160 63674 113216 63676
rect 112920 63622 112966 63674
rect 112966 63622 112976 63674
rect 113000 63622 113030 63674
rect 113030 63622 113042 63674
rect 113042 63622 113056 63674
rect 113080 63622 113094 63674
rect 113094 63622 113106 63674
rect 113106 63622 113136 63674
rect 113160 63622 113170 63674
rect 113170 63622 113216 63674
rect 112920 63620 112976 63622
rect 113000 63620 113056 63622
rect 113080 63620 113136 63622
rect 113160 63620 113216 63622
rect 113656 63130 113712 63132
rect 113736 63130 113792 63132
rect 113816 63130 113872 63132
rect 113896 63130 113952 63132
rect 113656 63078 113702 63130
rect 113702 63078 113712 63130
rect 113736 63078 113766 63130
rect 113766 63078 113778 63130
rect 113778 63078 113792 63130
rect 113816 63078 113830 63130
rect 113830 63078 113842 63130
rect 113842 63078 113872 63130
rect 113896 63078 113906 63130
rect 113906 63078 113952 63130
rect 113656 63076 113712 63078
rect 113736 63076 113792 63078
rect 113816 63076 113872 63078
rect 113896 63076 113952 63078
rect 112920 62586 112976 62588
rect 113000 62586 113056 62588
rect 113080 62586 113136 62588
rect 113160 62586 113216 62588
rect 112920 62534 112966 62586
rect 112966 62534 112976 62586
rect 113000 62534 113030 62586
rect 113030 62534 113042 62586
rect 113042 62534 113056 62586
rect 113080 62534 113094 62586
rect 113094 62534 113106 62586
rect 113106 62534 113136 62586
rect 113160 62534 113170 62586
rect 113170 62534 113216 62586
rect 112920 62532 112976 62534
rect 113000 62532 113056 62534
rect 113080 62532 113136 62534
rect 113160 62532 113216 62534
rect 113656 62042 113712 62044
rect 113736 62042 113792 62044
rect 113816 62042 113872 62044
rect 113896 62042 113952 62044
rect 113656 61990 113702 62042
rect 113702 61990 113712 62042
rect 113736 61990 113766 62042
rect 113766 61990 113778 62042
rect 113778 61990 113792 62042
rect 113816 61990 113830 62042
rect 113830 61990 113842 62042
rect 113842 61990 113872 62042
rect 113896 61990 113906 62042
rect 113906 61990 113952 62042
rect 113656 61988 113712 61990
rect 113736 61988 113792 61990
rect 113816 61988 113872 61990
rect 113896 61988 113952 61990
rect 112920 61498 112976 61500
rect 113000 61498 113056 61500
rect 113080 61498 113136 61500
rect 113160 61498 113216 61500
rect 112920 61446 112966 61498
rect 112966 61446 112976 61498
rect 113000 61446 113030 61498
rect 113030 61446 113042 61498
rect 113042 61446 113056 61498
rect 113080 61446 113094 61498
rect 113094 61446 113106 61498
rect 113106 61446 113136 61498
rect 113160 61446 113170 61498
rect 113170 61446 113216 61498
rect 112920 61444 112976 61446
rect 113000 61444 113056 61446
rect 113080 61444 113136 61446
rect 113160 61444 113216 61446
rect 113656 60954 113712 60956
rect 113736 60954 113792 60956
rect 113816 60954 113872 60956
rect 113896 60954 113952 60956
rect 113656 60902 113702 60954
rect 113702 60902 113712 60954
rect 113736 60902 113766 60954
rect 113766 60902 113778 60954
rect 113778 60902 113792 60954
rect 113816 60902 113830 60954
rect 113830 60902 113842 60954
rect 113842 60902 113872 60954
rect 113896 60902 113906 60954
rect 113906 60902 113952 60954
rect 113656 60900 113712 60902
rect 113736 60900 113792 60902
rect 113816 60900 113872 60902
rect 113896 60900 113952 60902
rect 112920 60410 112976 60412
rect 113000 60410 113056 60412
rect 113080 60410 113136 60412
rect 113160 60410 113216 60412
rect 112920 60358 112966 60410
rect 112966 60358 112976 60410
rect 113000 60358 113030 60410
rect 113030 60358 113042 60410
rect 113042 60358 113056 60410
rect 113080 60358 113094 60410
rect 113094 60358 113106 60410
rect 113106 60358 113136 60410
rect 113160 60358 113170 60410
rect 113170 60358 113216 60410
rect 112920 60356 112976 60358
rect 113000 60356 113056 60358
rect 113080 60356 113136 60358
rect 113160 60356 113216 60358
rect 113656 59866 113712 59868
rect 113736 59866 113792 59868
rect 113816 59866 113872 59868
rect 113896 59866 113952 59868
rect 113656 59814 113702 59866
rect 113702 59814 113712 59866
rect 113736 59814 113766 59866
rect 113766 59814 113778 59866
rect 113778 59814 113792 59866
rect 113816 59814 113830 59866
rect 113830 59814 113842 59866
rect 113842 59814 113872 59866
rect 113896 59814 113906 59866
rect 113906 59814 113952 59866
rect 113656 59812 113712 59814
rect 113736 59812 113792 59814
rect 113816 59812 113872 59814
rect 113896 59812 113952 59814
rect 112920 59322 112976 59324
rect 113000 59322 113056 59324
rect 113080 59322 113136 59324
rect 113160 59322 113216 59324
rect 112920 59270 112966 59322
rect 112966 59270 112976 59322
rect 113000 59270 113030 59322
rect 113030 59270 113042 59322
rect 113042 59270 113056 59322
rect 113080 59270 113094 59322
rect 113094 59270 113106 59322
rect 113106 59270 113136 59322
rect 113160 59270 113170 59322
rect 113170 59270 113216 59322
rect 112920 59268 112976 59270
rect 113000 59268 113056 59270
rect 113080 59268 113136 59270
rect 113160 59268 113216 59270
rect 113656 58778 113712 58780
rect 113736 58778 113792 58780
rect 113816 58778 113872 58780
rect 113896 58778 113952 58780
rect 113656 58726 113702 58778
rect 113702 58726 113712 58778
rect 113736 58726 113766 58778
rect 113766 58726 113778 58778
rect 113778 58726 113792 58778
rect 113816 58726 113830 58778
rect 113830 58726 113842 58778
rect 113842 58726 113872 58778
rect 113896 58726 113906 58778
rect 113906 58726 113952 58778
rect 113656 58724 113712 58726
rect 113736 58724 113792 58726
rect 113816 58724 113872 58726
rect 113896 58724 113952 58726
rect 112920 58234 112976 58236
rect 113000 58234 113056 58236
rect 113080 58234 113136 58236
rect 113160 58234 113216 58236
rect 112920 58182 112966 58234
rect 112966 58182 112976 58234
rect 113000 58182 113030 58234
rect 113030 58182 113042 58234
rect 113042 58182 113056 58234
rect 113080 58182 113094 58234
rect 113094 58182 113106 58234
rect 113106 58182 113136 58234
rect 113160 58182 113170 58234
rect 113170 58182 113216 58234
rect 112920 58180 112976 58182
rect 113000 58180 113056 58182
rect 113080 58180 113136 58182
rect 113160 58180 113216 58182
rect 113656 57690 113712 57692
rect 113736 57690 113792 57692
rect 113816 57690 113872 57692
rect 113896 57690 113952 57692
rect 113656 57638 113702 57690
rect 113702 57638 113712 57690
rect 113736 57638 113766 57690
rect 113766 57638 113778 57690
rect 113778 57638 113792 57690
rect 113816 57638 113830 57690
rect 113830 57638 113842 57690
rect 113842 57638 113872 57690
rect 113896 57638 113906 57690
rect 113906 57638 113952 57690
rect 113656 57636 113712 57638
rect 113736 57636 113792 57638
rect 113816 57636 113872 57638
rect 113896 57636 113952 57638
rect 112920 57146 112976 57148
rect 113000 57146 113056 57148
rect 113080 57146 113136 57148
rect 113160 57146 113216 57148
rect 112920 57094 112966 57146
rect 112966 57094 112976 57146
rect 113000 57094 113030 57146
rect 113030 57094 113042 57146
rect 113042 57094 113056 57146
rect 113080 57094 113094 57146
rect 113094 57094 113106 57146
rect 113106 57094 113136 57146
rect 113160 57094 113170 57146
rect 113170 57094 113216 57146
rect 112920 57092 112976 57094
rect 113000 57092 113056 57094
rect 113080 57092 113136 57094
rect 113160 57092 113216 57094
rect 113656 56602 113712 56604
rect 113736 56602 113792 56604
rect 113816 56602 113872 56604
rect 113896 56602 113952 56604
rect 113656 56550 113702 56602
rect 113702 56550 113712 56602
rect 113736 56550 113766 56602
rect 113766 56550 113778 56602
rect 113778 56550 113792 56602
rect 113816 56550 113830 56602
rect 113830 56550 113842 56602
rect 113842 56550 113872 56602
rect 113896 56550 113906 56602
rect 113906 56550 113952 56602
rect 113656 56548 113712 56550
rect 113736 56548 113792 56550
rect 113816 56548 113872 56550
rect 113896 56548 113952 56550
rect 112920 56058 112976 56060
rect 113000 56058 113056 56060
rect 113080 56058 113136 56060
rect 113160 56058 113216 56060
rect 112920 56006 112966 56058
rect 112966 56006 112976 56058
rect 113000 56006 113030 56058
rect 113030 56006 113042 56058
rect 113042 56006 113056 56058
rect 113080 56006 113094 56058
rect 113094 56006 113106 56058
rect 113106 56006 113136 56058
rect 113160 56006 113170 56058
rect 113170 56006 113216 56058
rect 112920 56004 112976 56006
rect 113000 56004 113056 56006
rect 113080 56004 113136 56006
rect 113160 56004 113216 56006
rect 113656 55514 113712 55516
rect 113736 55514 113792 55516
rect 113816 55514 113872 55516
rect 113896 55514 113952 55516
rect 113656 55462 113702 55514
rect 113702 55462 113712 55514
rect 113736 55462 113766 55514
rect 113766 55462 113778 55514
rect 113778 55462 113792 55514
rect 113816 55462 113830 55514
rect 113830 55462 113842 55514
rect 113842 55462 113872 55514
rect 113896 55462 113906 55514
rect 113906 55462 113952 55514
rect 113656 55460 113712 55462
rect 113736 55460 113792 55462
rect 113816 55460 113872 55462
rect 113896 55460 113952 55462
rect 112920 54970 112976 54972
rect 113000 54970 113056 54972
rect 113080 54970 113136 54972
rect 113160 54970 113216 54972
rect 112920 54918 112966 54970
rect 112966 54918 112976 54970
rect 113000 54918 113030 54970
rect 113030 54918 113042 54970
rect 113042 54918 113056 54970
rect 113080 54918 113094 54970
rect 113094 54918 113106 54970
rect 113106 54918 113136 54970
rect 113160 54918 113170 54970
rect 113170 54918 113216 54970
rect 112920 54916 112976 54918
rect 113000 54916 113056 54918
rect 113080 54916 113136 54918
rect 113160 54916 113216 54918
rect 113656 54426 113712 54428
rect 113736 54426 113792 54428
rect 113816 54426 113872 54428
rect 113896 54426 113952 54428
rect 113656 54374 113702 54426
rect 113702 54374 113712 54426
rect 113736 54374 113766 54426
rect 113766 54374 113778 54426
rect 113778 54374 113792 54426
rect 113816 54374 113830 54426
rect 113830 54374 113842 54426
rect 113842 54374 113872 54426
rect 113896 54374 113906 54426
rect 113906 54374 113952 54426
rect 113656 54372 113712 54374
rect 113736 54372 113792 54374
rect 113816 54372 113872 54374
rect 113896 54372 113952 54374
rect 112920 53882 112976 53884
rect 113000 53882 113056 53884
rect 113080 53882 113136 53884
rect 113160 53882 113216 53884
rect 112920 53830 112966 53882
rect 112966 53830 112976 53882
rect 113000 53830 113030 53882
rect 113030 53830 113042 53882
rect 113042 53830 113056 53882
rect 113080 53830 113094 53882
rect 113094 53830 113106 53882
rect 113106 53830 113136 53882
rect 113160 53830 113170 53882
rect 113170 53830 113216 53882
rect 112920 53828 112976 53830
rect 113000 53828 113056 53830
rect 113080 53828 113136 53830
rect 113160 53828 113216 53830
rect 113656 53338 113712 53340
rect 113736 53338 113792 53340
rect 113816 53338 113872 53340
rect 113896 53338 113952 53340
rect 113656 53286 113702 53338
rect 113702 53286 113712 53338
rect 113736 53286 113766 53338
rect 113766 53286 113778 53338
rect 113778 53286 113792 53338
rect 113816 53286 113830 53338
rect 113830 53286 113842 53338
rect 113842 53286 113872 53338
rect 113896 53286 113906 53338
rect 113906 53286 113952 53338
rect 113656 53284 113712 53286
rect 113736 53284 113792 53286
rect 113816 53284 113872 53286
rect 113896 53284 113952 53286
rect 112920 52794 112976 52796
rect 113000 52794 113056 52796
rect 113080 52794 113136 52796
rect 113160 52794 113216 52796
rect 112920 52742 112966 52794
rect 112966 52742 112976 52794
rect 113000 52742 113030 52794
rect 113030 52742 113042 52794
rect 113042 52742 113056 52794
rect 113080 52742 113094 52794
rect 113094 52742 113106 52794
rect 113106 52742 113136 52794
rect 113160 52742 113170 52794
rect 113170 52742 113216 52794
rect 112920 52740 112976 52742
rect 113000 52740 113056 52742
rect 113080 52740 113136 52742
rect 113160 52740 113216 52742
rect 9678 44192 9734 44202
rect 9678 44146 9680 44192
rect 9680 44146 9732 44192
rect 9732 44146 9734 44192
rect 9678 42922 9734 42978
rect 9678 41154 9734 41210
rect 9678 40066 9734 40122
rect 9678 38434 9734 38490
rect 9494 37482 9550 37538
rect 9494 35760 9550 35770
rect 9494 35714 9496 35760
rect 9496 35714 9548 35760
rect 9548 35714 9550 35760
rect 106922 26560 106978 26616
rect 107014 24928 107070 24984
rect 109406 33260 109408 33280
rect 109408 33260 109460 33280
rect 109460 33260 109462 33280
rect 109406 33224 109462 33260
rect 113656 52250 113712 52252
rect 113736 52250 113792 52252
rect 113816 52250 113872 52252
rect 113896 52250 113952 52252
rect 113656 52198 113702 52250
rect 113702 52198 113712 52250
rect 113736 52198 113766 52250
rect 113766 52198 113778 52250
rect 113778 52198 113792 52250
rect 113816 52198 113830 52250
rect 113830 52198 113842 52250
rect 113842 52198 113872 52250
rect 113896 52198 113906 52250
rect 113906 52198 113952 52250
rect 113656 52196 113712 52198
rect 113736 52196 113792 52198
rect 113816 52196 113872 52198
rect 113896 52196 113952 52198
rect 112920 51706 112976 51708
rect 113000 51706 113056 51708
rect 113080 51706 113136 51708
rect 113160 51706 113216 51708
rect 112920 51654 112966 51706
rect 112966 51654 112976 51706
rect 113000 51654 113030 51706
rect 113030 51654 113042 51706
rect 113042 51654 113056 51706
rect 113080 51654 113094 51706
rect 113094 51654 113106 51706
rect 113106 51654 113136 51706
rect 113160 51654 113170 51706
rect 113170 51654 113216 51706
rect 112920 51652 112976 51654
rect 113000 51652 113056 51654
rect 113080 51652 113136 51654
rect 113160 51652 113216 51654
rect 113656 51162 113712 51164
rect 113736 51162 113792 51164
rect 113816 51162 113872 51164
rect 113896 51162 113952 51164
rect 113656 51110 113702 51162
rect 113702 51110 113712 51162
rect 113736 51110 113766 51162
rect 113766 51110 113778 51162
rect 113778 51110 113792 51162
rect 113816 51110 113830 51162
rect 113830 51110 113842 51162
rect 113842 51110 113872 51162
rect 113896 51110 113906 51162
rect 113906 51110 113952 51162
rect 113656 51108 113712 51110
rect 113736 51108 113792 51110
rect 113816 51108 113872 51110
rect 113896 51108 113952 51110
rect 112920 50618 112976 50620
rect 113000 50618 113056 50620
rect 113080 50618 113136 50620
rect 113160 50618 113216 50620
rect 112920 50566 112966 50618
rect 112966 50566 112976 50618
rect 113000 50566 113030 50618
rect 113030 50566 113042 50618
rect 113042 50566 113056 50618
rect 113080 50566 113094 50618
rect 113094 50566 113106 50618
rect 113106 50566 113136 50618
rect 113160 50566 113170 50618
rect 113170 50566 113216 50618
rect 112920 50564 112976 50566
rect 113000 50564 113056 50566
rect 113080 50564 113136 50566
rect 113160 50564 113216 50566
rect 113656 50074 113712 50076
rect 113736 50074 113792 50076
rect 113816 50074 113872 50076
rect 113896 50074 113952 50076
rect 113656 50022 113702 50074
rect 113702 50022 113712 50074
rect 113736 50022 113766 50074
rect 113766 50022 113778 50074
rect 113778 50022 113792 50074
rect 113816 50022 113830 50074
rect 113830 50022 113842 50074
rect 113842 50022 113872 50074
rect 113896 50022 113906 50074
rect 113906 50022 113952 50074
rect 113656 50020 113712 50022
rect 113736 50020 113792 50022
rect 113816 50020 113872 50022
rect 113896 50020 113952 50022
rect 112920 49530 112976 49532
rect 113000 49530 113056 49532
rect 113080 49530 113136 49532
rect 113160 49530 113216 49532
rect 112920 49478 112966 49530
rect 112966 49478 112976 49530
rect 113000 49478 113030 49530
rect 113030 49478 113042 49530
rect 113042 49478 113056 49530
rect 113080 49478 113094 49530
rect 113094 49478 113106 49530
rect 113106 49478 113136 49530
rect 113160 49478 113170 49530
rect 113170 49478 113216 49530
rect 112920 49476 112976 49478
rect 113000 49476 113056 49478
rect 113080 49476 113136 49478
rect 113160 49476 113216 49478
rect 113656 48986 113712 48988
rect 113736 48986 113792 48988
rect 113816 48986 113872 48988
rect 113896 48986 113952 48988
rect 113656 48934 113702 48986
rect 113702 48934 113712 48986
rect 113736 48934 113766 48986
rect 113766 48934 113778 48986
rect 113778 48934 113792 48986
rect 113816 48934 113830 48986
rect 113830 48934 113842 48986
rect 113842 48934 113872 48986
rect 113896 48934 113906 48986
rect 113906 48934 113952 48986
rect 113656 48932 113712 48934
rect 113736 48932 113792 48934
rect 113816 48932 113872 48934
rect 113896 48932 113952 48934
rect 112920 48442 112976 48444
rect 113000 48442 113056 48444
rect 113080 48442 113136 48444
rect 113160 48442 113216 48444
rect 112920 48390 112966 48442
rect 112966 48390 112976 48442
rect 113000 48390 113030 48442
rect 113030 48390 113042 48442
rect 113042 48390 113056 48442
rect 113080 48390 113094 48442
rect 113094 48390 113106 48442
rect 113106 48390 113136 48442
rect 113160 48390 113170 48442
rect 113170 48390 113216 48442
rect 112920 48388 112976 48390
rect 113000 48388 113056 48390
rect 113080 48388 113136 48390
rect 113160 48388 113216 48390
rect 113656 47898 113712 47900
rect 113736 47898 113792 47900
rect 113816 47898 113872 47900
rect 113896 47898 113952 47900
rect 113656 47846 113702 47898
rect 113702 47846 113712 47898
rect 113736 47846 113766 47898
rect 113766 47846 113778 47898
rect 113778 47846 113792 47898
rect 113816 47846 113830 47898
rect 113830 47846 113842 47898
rect 113842 47846 113872 47898
rect 113896 47846 113906 47898
rect 113906 47846 113952 47898
rect 113656 47844 113712 47846
rect 113736 47844 113792 47846
rect 113816 47844 113872 47846
rect 113896 47844 113952 47846
rect 112920 47354 112976 47356
rect 113000 47354 113056 47356
rect 113080 47354 113136 47356
rect 113160 47354 113216 47356
rect 112920 47302 112966 47354
rect 112966 47302 112976 47354
rect 113000 47302 113030 47354
rect 113030 47302 113042 47354
rect 113042 47302 113056 47354
rect 113080 47302 113094 47354
rect 113094 47302 113106 47354
rect 113106 47302 113136 47354
rect 113160 47302 113170 47354
rect 113170 47302 113216 47354
rect 112920 47300 112976 47302
rect 113000 47300 113056 47302
rect 113080 47300 113136 47302
rect 113160 47300 113216 47302
rect 113656 46810 113712 46812
rect 113736 46810 113792 46812
rect 113816 46810 113872 46812
rect 113896 46810 113952 46812
rect 113656 46758 113702 46810
rect 113702 46758 113712 46810
rect 113736 46758 113766 46810
rect 113766 46758 113778 46810
rect 113778 46758 113792 46810
rect 113816 46758 113830 46810
rect 113830 46758 113842 46810
rect 113842 46758 113872 46810
rect 113896 46758 113906 46810
rect 113906 46758 113952 46810
rect 113656 46756 113712 46758
rect 113736 46756 113792 46758
rect 113816 46756 113872 46758
rect 113896 46756 113952 46758
rect 112920 46266 112976 46268
rect 113000 46266 113056 46268
rect 113080 46266 113136 46268
rect 113160 46266 113216 46268
rect 112920 46214 112966 46266
rect 112966 46214 112976 46266
rect 113000 46214 113030 46266
rect 113030 46214 113042 46266
rect 113042 46214 113056 46266
rect 113080 46214 113094 46266
rect 113094 46214 113106 46266
rect 113106 46214 113136 46266
rect 113160 46214 113170 46266
rect 113170 46214 113216 46266
rect 112920 46212 112976 46214
rect 113000 46212 113056 46214
rect 113080 46212 113136 46214
rect 113160 46212 113216 46214
rect 113656 45722 113712 45724
rect 113736 45722 113792 45724
rect 113816 45722 113872 45724
rect 113896 45722 113952 45724
rect 113656 45670 113702 45722
rect 113702 45670 113712 45722
rect 113736 45670 113766 45722
rect 113766 45670 113778 45722
rect 113778 45670 113792 45722
rect 113816 45670 113830 45722
rect 113830 45670 113842 45722
rect 113842 45670 113872 45722
rect 113896 45670 113906 45722
rect 113906 45670 113952 45722
rect 113656 45668 113712 45670
rect 113736 45668 113792 45670
rect 113816 45668 113872 45670
rect 113896 45668 113952 45670
rect 112920 45178 112976 45180
rect 113000 45178 113056 45180
rect 113080 45178 113136 45180
rect 113160 45178 113216 45180
rect 112920 45126 112966 45178
rect 112966 45126 112976 45178
rect 113000 45126 113030 45178
rect 113030 45126 113042 45178
rect 113042 45126 113056 45178
rect 113080 45126 113094 45178
rect 113094 45126 113106 45178
rect 113106 45126 113136 45178
rect 113160 45126 113170 45178
rect 113170 45126 113216 45178
rect 112920 45124 112976 45126
rect 113000 45124 113056 45126
rect 113080 45124 113136 45126
rect 113160 45124 113216 45126
rect 113656 44634 113712 44636
rect 113736 44634 113792 44636
rect 113816 44634 113872 44636
rect 113896 44634 113952 44636
rect 113656 44582 113702 44634
rect 113702 44582 113712 44634
rect 113736 44582 113766 44634
rect 113766 44582 113778 44634
rect 113778 44582 113792 44634
rect 113816 44582 113830 44634
rect 113830 44582 113842 44634
rect 113842 44582 113872 44634
rect 113896 44582 113906 44634
rect 113906 44582 113952 44634
rect 113656 44580 113712 44582
rect 113736 44580 113792 44582
rect 113816 44580 113872 44582
rect 113896 44580 113952 44582
rect 112920 44090 112976 44092
rect 113000 44090 113056 44092
rect 113080 44090 113136 44092
rect 113160 44090 113216 44092
rect 112920 44038 112966 44090
rect 112966 44038 112976 44090
rect 113000 44038 113030 44090
rect 113030 44038 113042 44090
rect 113042 44038 113056 44090
rect 113080 44038 113094 44090
rect 113094 44038 113106 44090
rect 113106 44038 113136 44090
rect 113160 44038 113170 44090
rect 113170 44038 113216 44090
rect 112920 44036 112976 44038
rect 113000 44036 113056 44038
rect 113080 44036 113136 44038
rect 113160 44036 113216 44038
rect 113656 43546 113712 43548
rect 113736 43546 113792 43548
rect 113816 43546 113872 43548
rect 113896 43546 113952 43548
rect 113656 43494 113702 43546
rect 113702 43494 113712 43546
rect 113736 43494 113766 43546
rect 113766 43494 113778 43546
rect 113778 43494 113792 43546
rect 113816 43494 113830 43546
rect 113830 43494 113842 43546
rect 113842 43494 113872 43546
rect 113896 43494 113906 43546
rect 113906 43494 113952 43546
rect 113656 43492 113712 43494
rect 113736 43492 113792 43494
rect 113816 43492 113872 43494
rect 113896 43492 113952 43494
rect 112920 43002 112976 43004
rect 113000 43002 113056 43004
rect 113080 43002 113136 43004
rect 113160 43002 113216 43004
rect 112920 42950 112966 43002
rect 112966 42950 112976 43002
rect 113000 42950 113030 43002
rect 113030 42950 113042 43002
rect 113042 42950 113056 43002
rect 113080 42950 113094 43002
rect 113094 42950 113106 43002
rect 113106 42950 113136 43002
rect 113160 42950 113170 43002
rect 113170 42950 113216 43002
rect 112920 42948 112976 42950
rect 113000 42948 113056 42950
rect 113080 42948 113136 42950
rect 113160 42948 113216 42950
rect 113656 42458 113712 42460
rect 113736 42458 113792 42460
rect 113816 42458 113872 42460
rect 113896 42458 113952 42460
rect 113656 42406 113702 42458
rect 113702 42406 113712 42458
rect 113736 42406 113766 42458
rect 113766 42406 113778 42458
rect 113778 42406 113792 42458
rect 113816 42406 113830 42458
rect 113830 42406 113842 42458
rect 113842 42406 113872 42458
rect 113896 42406 113906 42458
rect 113906 42406 113952 42458
rect 113656 42404 113712 42406
rect 113736 42404 113792 42406
rect 113816 42404 113872 42406
rect 113896 42404 113952 42406
rect 112920 41914 112976 41916
rect 113000 41914 113056 41916
rect 113080 41914 113136 41916
rect 113160 41914 113216 41916
rect 112920 41862 112966 41914
rect 112966 41862 112976 41914
rect 113000 41862 113030 41914
rect 113030 41862 113042 41914
rect 113042 41862 113056 41914
rect 113080 41862 113094 41914
rect 113094 41862 113106 41914
rect 113106 41862 113136 41914
rect 113160 41862 113170 41914
rect 113170 41862 113216 41914
rect 112920 41860 112976 41862
rect 113000 41860 113056 41862
rect 113080 41860 113136 41862
rect 113160 41860 113216 41862
rect 113656 41370 113712 41372
rect 113736 41370 113792 41372
rect 113816 41370 113872 41372
rect 113896 41370 113952 41372
rect 113656 41318 113702 41370
rect 113702 41318 113712 41370
rect 113736 41318 113766 41370
rect 113766 41318 113778 41370
rect 113778 41318 113792 41370
rect 113816 41318 113830 41370
rect 113830 41318 113842 41370
rect 113842 41318 113872 41370
rect 113896 41318 113906 41370
rect 113906 41318 113952 41370
rect 113656 41316 113712 41318
rect 113736 41316 113792 41318
rect 113816 41316 113872 41318
rect 113896 41316 113952 41318
rect 112920 40826 112976 40828
rect 113000 40826 113056 40828
rect 113080 40826 113136 40828
rect 113160 40826 113216 40828
rect 112920 40774 112966 40826
rect 112966 40774 112976 40826
rect 113000 40774 113030 40826
rect 113030 40774 113042 40826
rect 113042 40774 113056 40826
rect 113080 40774 113094 40826
rect 113094 40774 113106 40826
rect 113106 40774 113136 40826
rect 113160 40774 113170 40826
rect 113170 40774 113216 40826
rect 112920 40772 112976 40774
rect 113000 40772 113056 40774
rect 113080 40772 113136 40774
rect 113160 40772 113216 40774
rect 112920 39738 112976 39740
rect 113000 39738 113056 39740
rect 113080 39738 113136 39740
rect 113160 39738 113216 39740
rect 112920 39686 112966 39738
rect 112966 39686 112976 39738
rect 113000 39686 113030 39738
rect 113030 39686 113042 39738
rect 113042 39686 113056 39738
rect 113080 39686 113094 39738
rect 113094 39686 113106 39738
rect 113106 39686 113136 39738
rect 113160 39686 113170 39738
rect 113170 39686 113216 39738
rect 112920 39684 112976 39686
rect 113000 39684 113056 39686
rect 113080 39684 113136 39686
rect 113160 39684 113216 39686
rect 112920 38650 112976 38652
rect 113000 38650 113056 38652
rect 113080 38650 113136 38652
rect 113160 38650 113216 38652
rect 112920 38598 112966 38650
rect 112966 38598 112976 38650
rect 113000 38598 113030 38650
rect 113030 38598 113042 38650
rect 113042 38598 113056 38650
rect 113080 38598 113094 38650
rect 113094 38598 113106 38650
rect 113106 38598 113136 38650
rect 113160 38598 113170 38650
rect 113170 38598 113216 38650
rect 112920 38596 112976 38598
rect 113000 38596 113056 38598
rect 113080 38596 113136 38598
rect 113160 38596 113216 38598
rect 113656 40282 113712 40284
rect 113736 40282 113792 40284
rect 113816 40282 113872 40284
rect 113896 40282 113952 40284
rect 113656 40230 113702 40282
rect 113702 40230 113712 40282
rect 113736 40230 113766 40282
rect 113766 40230 113778 40282
rect 113778 40230 113792 40282
rect 113816 40230 113830 40282
rect 113830 40230 113842 40282
rect 113842 40230 113872 40282
rect 113896 40230 113906 40282
rect 113906 40230 113952 40282
rect 113656 40228 113712 40230
rect 113736 40228 113792 40230
rect 113816 40228 113872 40230
rect 113896 40228 113952 40230
rect 113656 39194 113712 39196
rect 113736 39194 113792 39196
rect 113816 39194 113872 39196
rect 113896 39194 113952 39196
rect 113656 39142 113702 39194
rect 113702 39142 113712 39194
rect 113736 39142 113766 39194
rect 113766 39142 113778 39194
rect 113778 39142 113792 39194
rect 113816 39142 113830 39194
rect 113830 39142 113842 39194
rect 113842 39142 113872 39194
rect 113896 39142 113906 39194
rect 113906 39142 113952 39194
rect 113656 39140 113712 39142
rect 113736 39140 113792 39142
rect 113816 39140 113872 39142
rect 113896 39140 113952 39142
rect 113656 38106 113712 38108
rect 113736 38106 113792 38108
rect 113816 38106 113872 38108
rect 113896 38106 113952 38108
rect 113656 38054 113702 38106
rect 113702 38054 113712 38106
rect 113736 38054 113766 38106
rect 113766 38054 113778 38106
rect 113778 38054 113792 38106
rect 113816 38054 113830 38106
rect 113830 38054 113842 38106
rect 113842 38054 113872 38106
rect 113896 38054 113906 38106
rect 113906 38054 113952 38106
rect 113656 38052 113712 38054
rect 113736 38052 113792 38054
rect 113816 38052 113872 38054
rect 113896 38052 113952 38054
rect 112920 37562 112976 37564
rect 113000 37562 113056 37564
rect 113080 37562 113136 37564
rect 113160 37562 113216 37564
rect 112920 37510 112966 37562
rect 112966 37510 112976 37562
rect 113000 37510 113030 37562
rect 113030 37510 113042 37562
rect 113042 37510 113056 37562
rect 113080 37510 113094 37562
rect 113094 37510 113106 37562
rect 113106 37510 113136 37562
rect 113160 37510 113170 37562
rect 113170 37510 113216 37562
rect 112920 37508 112976 37510
rect 113000 37508 113056 37510
rect 113080 37508 113136 37510
rect 113160 37508 113216 37510
rect 113454 36760 113510 36816
rect 112920 36474 112976 36476
rect 113000 36474 113056 36476
rect 113080 36474 113136 36476
rect 113160 36474 113216 36476
rect 112920 36422 112966 36474
rect 112966 36422 112976 36474
rect 113000 36422 113030 36474
rect 113030 36422 113042 36474
rect 113042 36422 113056 36474
rect 113080 36422 113094 36474
rect 113094 36422 113106 36474
rect 113106 36422 113136 36474
rect 113160 36422 113170 36474
rect 113170 36422 113216 36474
rect 112920 36420 112976 36422
rect 113000 36420 113056 36422
rect 113080 36420 113136 36422
rect 113160 36420 113216 36422
rect 107106 23568 107162 23624
rect 9678 17218 9734 17274
rect 9678 15586 9734 15642
rect 106462 11872 106518 11928
rect 15842 9832 15898 9888
rect 92754 9832 92810 9888
rect 111338 31184 111394 31240
rect 112920 35386 112976 35388
rect 113000 35386 113056 35388
rect 113080 35386 113136 35388
rect 113160 35386 113216 35388
rect 112920 35334 112966 35386
rect 112966 35334 112976 35386
rect 113000 35334 113030 35386
rect 113030 35334 113042 35386
rect 113042 35334 113056 35386
rect 113080 35334 113094 35386
rect 113094 35334 113106 35386
rect 113106 35334 113136 35386
rect 113160 35334 113170 35386
rect 113170 35334 113216 35386
rect 112920 35332 112976 35334
rect 113000 35332 113056 35334
rect 113080 35332 113136 35334
rect 113160 35332 113216 35334
rect 113656 37018 113712 37020
rect 113736 37018 113792 37020
rect 113816 37018 113872 37020
rect 113896 37018 113952 37020
rect 113656 36966 113702 37018
rect 113702 36966 113712 37018
rect 113736 36966 113766 37018
rect 113766 36966 113778 37018
rect 113778 36966 113792 37018
rect 113816 36966 113830 37018
rect 113830 36966 113842 37018
rect 113842 36966 113872 37018
rect 113896 36966 113906 37018
rect 113906 36966 113952 37018
rect 113656 36964 113712 36966
rect 113736 36964 113792 36966
rect 113816 36964 113872 36966
rect 113896 36964 113952 36966
rect 114006 36780 114062 36816
rect 114006 36760 114008 36780
rect 114008 36760 114060 36780
rect 114060 36760 114062 36780
rect 113656 35930 113712 35932
rect 113736 35930 113792 35932
rect 113816 35930 113872 35932
rect 113896 35930 113952 35932
rect 113656 35878 113702 35930
rect 113702 35878 113712 35930
rect 113736 35878 113766 35930
rect 113766 35878 113778 35930
rect 113778 35878 113792 35930
rect 113816 35878 113830 35930
rect 113830 35878 113842 35930
rect 113842 35878 113872 35930
rect 113896 35878 113906 35930
rect 113906 35878 113952 35930
rect 113656 35876 113712 35878
rect 113736 35876 113792 35878
rect 113816 35876 113872 35878
rect 113896 35876 113952 35878
rect 115110 36796 115112 36816
rect 115112 36796 115164 36816
rect 115164 36796 115166 36816
rect 115110 36760 115166 36796
rect 112920 34298 112976 34300
rect 113000 34298 113056 34300
rect 113080 34298 113136 34300
rect 113160 34298 113216 34300
rect 112920 34246 112966 34298
rect 112966 34246 112976 34298
rect 113000 34246 113030 34298
rect 113030 34246 113042 34298
rect 113042 34246 113056 34298
rect 113080 34246 113094 34298
rect 113094 34246 113106 34298
rect 113106 34246 113136 34298
rect 113160 34246 113170 34298
rect 113170 34246 113216 34298
rect 112920 34244 112976 34246
rect 113000 34244 113056 34246
rect 113080 34244 113136 34246
rect 113160 34244 113216 34246
rect 113656 34842 113712 34844
rect 113736 34842 113792 34844
rect 113816 34842 113872 34844
rect 113896 34842 113952 34844
rect 113656 34790 113702 34842
rect 113702 34790 113712 34842
rect 113736 34790 113766 34842
rect 113766 34790 113778 34842
rect 113778 34790 113792 34842
rect 113816 34790 113830 34842
rect 113830 34790 113842 34842
rect 113842 34790 113872 34842
rect 113896 34790 113906 34842
rect 113906 34790 113952 34842
rect 113656 34788 113712 34790
rect 113736 34788 113792 34790
rect 113816 34788 113872 34790
rect 113896 34788 113952 34790
rect 112920 33210 112976 33212
rect 113000 33210 113056 33212
rect 113080 33210 113136 33212
rect 113160 33210 113216 33212
rect 112920 33158 112966 33210
rect 112966 33158 112976 33210
rect 113000 33158 113030 33210
rect 113030 33158 113042 33210
rect 113042 33158 113056 33210
rect 113080 33158 113094 33210
rect 113094 33158 113106 33210
rect 113106 33158 113136 33210
rect 113160 33158 113170 33210
rect 113170 33158 113216 33210
rect 112920 33156 112976 33158
rect 113000 33156 113056 33158
rect 113080 33156 113136 33158
rect 113160 33156 113216 33158
rect 112920 32122 112976 32124
rect 113000 32122 113056 32124
rect 113080 32122 113136 32124
rect 113160 32122 113216 32124
rect 112920 32070 112966 32122
rect 112966 32070 112976 32122
rect 113000 32070 113030 32122
rect 113030 32070 113042 32122
rect 113042 32070 113056 32122
rect 113080 32070 113094 32122
rect 113094 32070 113106 32122
rect 113106 32070 113136 32122
rect 113160 32070 113170 32122
rect 113170 32070 113216 32122
rect 112920 32068 112976 32070
rect 113000 32068 113056 32070
rect 113080 32068 113136 32070
rect 113160 32068 113216 32070
rect 111890 31184 111946 31240
rect 112534 30776 112590 30832
rect 112920 31034 112976 31036
rect 113000 31034 113056 31036
rect 113080 31034 113136 31036
rect 113160 31034 113216 31036
rect 112920 30982 112966 31034
rect 112966 30982 112976 31034
rect 113000 30982 113030 31034
rect 113030 30982 113042 31034
rect 113042 30982 113056 31034
rect 113080 30982 113094 31034
rect 113094 30982 113106 31034
rect 113106 30982 113136 31034
rect 113160 30982 113170 31034
rect 113170 30982 113216 31034
rect 112920 30980 112976 30982
rect 113000 30980 113056 30982
rect 113080 30980 113136 30982
rect 113160 30980 113216 30982
rect 113086 30776 113142 30832
rect 114098 34604 114154 34640
rect 114098 34584 114100 34604
rect 114100 34584 114152 34604
rect 114152 34584 114154 34604
rect 113656 33754 113712 33756
rect 113736 33754 113792 33756
rect 113816 33754 113872 33756
rect 113896 33754 113952 33756
rect 113656 33702 113702 33754
rect 113702 33702 113712 33754
rect 113736 33702 113766 33754
rect 113766 33702 113778 33754
rect 113778 33702 113792 33754
rect 113816 33702 113830 33754
rect 113830 33702 113842 33754
rect 113842 33702 113872 33754
rect 113896 33702 113906 33754
rect 113906 33702 113952 33754
rect 113656 33700 113712 33702
rect 113736 33700 113792 33702
rect 113816 33700 113872 33702
rect 113896 33700 113952 33702
rect 113656 32666 113712 32668
rect 113736 32666 113792 32668
rect 113816 32666 113872 32668
rect 113896 32666 113952 32668
rect 113656 32614 113702 32666
rect 113702 32614 113712 32666
rect 113736 32614 113766 32666
rect 113766 32614 113778 32666
rect 113778 32614 113792 32666
rect 113816 32614 113830 32666
rect 113830 32614 113842 32666
rect 113842 32614 113872 32666
rect 113896 32614 113906 32666
rect 113906 32614 113952 32666
rect 113656 32612 113712 32614
rect 113736 32612 113792 32614
rect 113816 32612 113872 32614
rect 113896 32612 113952 32614
rect 114098 31900 114100 31920
rect 114100 31900 114152 31920
rect 114152 31900 114154 31920
rect 114098 31864 114154 31900
rect 113656 31578 113712 31580
rect 113736 31578 113792 31580
rect 113816 31578 113872 31580
rect 113896 31578 113952 31580
rect 113656 31526 113702 31578
rect 113702 31526 113712 31578
rect 113736 31526 113766 31578
rect 113766 31526 113778 31578
rect 113778 31526 113792 31578
rect 113816 31526 113830 31578
rect 113830 31526 113842 31578
rect 113842 31526 113872 31578
rect 113896 31526 113906 31578
rect 113906 31526 113952 31578
rect 113656 31524 113712 31526
rect 113736 31524 113792 31526
rect 113816 31524 113872 31526
rect 113896 31524 113952 31526
rect 114926 33940 114928 33960
rect 114928 33940 114980 33960
rect 114980 33940 114982 33960
rect 114926 33904 114982 33940
rect 112920 29946 112976 29948
rect 113000 29946 113056 29948
rect 113080 29946 113136 29948
rect 113160 29946 113216 29948
rect 112920 29894 112966 29946
rect 112966 29894 112976 29946
rect 113000 29894 113030 29946
rect 113030 29894 113042 29946
rect 113042 29894 113056 29946
rect 113080 29894 113094 29946
rect 113094 29894 113106 29946
rect 113106 29894 113136 29946
rect 113160 29894 113170 29946
rect 113170 29894 113216 29946
rect 112920 29892 112976 29894
rect 113000 29892 113056 29894
rect 113080 29892 113136 29894
rect 113160 29892 113216 29894
rect 112920 28858 112976 28860
rect 113000 28858 113056 28860
rect 113080 28858 113136 28860
rect 113160 28858 113216 28860
rect 112920 28806 112966 28858
rect 112966 28806 112976 28858
rect 113000 28806 113030 28858
rect 113030 28806 113042 28858
rect 113042 28806 113056 28858
rect 113080 28806 113094 28858
rect 113094 28806 113106 28858
rect 113106 28806 113136 28858
rect 113160 28806 113170 28858
rect 113170 28806 113216 28858
rect 112920 28804 112976 28806
rect 113000 28804 113056 28806
rect 113080 28804 113136 28806
rect 113160 28804 113216 28806
rect 114098 30776 114154 30832
rect 113822 30676 113824 30696
rect 113824 30676 113876 30696
rect 113876 30676 113878 30696
rect 113822 30640 113878 30676
rect 113656 30490 113712 30492
rect 113736 30490 113792 30492
rect 113816 30490 113872 30492
rect 113896 30490 113952 30492
rect 113656 30438 113702 30490
rect 113702 30438 113712 30490
rect 113736 30438 113766 30490
rect 113766 30438 113778 30490
rect 113778 30438 113792 30490
rect 113816 30438 113830 30490
rect 113830 30438 113842 30490
rect 113842 30438 113872 30490
rect 113896 30438 113906 30490
rect 113906 30438 113952 30490
rect 113656 30436 113712 30438
rect 113736 30436 113792 30438
rect 113816 30436 113872 30438
rect 113896 30436 113952 30438
rect 115294 33904 115350 33960
rect 115662 34604 115718 34640
rect 115662 34584 115664 34604
rect 115664 34584 115716 34604
rect 115716 34584 115718 34604
rect 114650 30676 114652 30696
rect 114652 30676 114704 30696
rect 114704 30676 114706 30696
rect 114650 30640 114706 30676
rect 113656 29402 113712 29404
rect 113736 29402 113792 29404
rect 113816 29402 113872 29404
rect 113896 29402 113952 29404
rect 113656 29350 113702 29402
rect 113702 29350 113712 29402
rect 113736 29350 113766 29402
rect 113766 29350 113778 29402
rect 113778 29350 113792 29402
rect 113816 29350 113830 29402
rect 113830 29350 113842 29402
rect 113842 29350 113872 29402
rect 113896 29350 113906 29402
rect 113906 29350 113952 29402
rect 113656 29348 113712 29350
rect 113736 29348 113792 29350
rect 113816 29348 113872 29350
rect 113896 29348 113952 29350
rect 113656 28314 113712 28316
rect 113736 28314 113792 28316
rect 113816 28314 113872 28316
rect 113896 28314 113952 28316
rect 113656 28262 113702 28314
rect 113702 28262 113712 28314
rect 113736 28262 113766 28314
rect 113766 28262 113778 28314
rect 113778 28262 113792 28314
rect 113816 28262 113830 28314
rect 113830 28262 113842 28314
rect 113842 28262 113872 28314
rect 113896 28262 113906 28314
rect 113906 28262 113952 28314
rect 113656 28260 113712 28262
rect 113736 28260 113792 28262
rect 113816 28260 113872 28262
rect 113896 28260 113952 28262
rect 112920 27770 112976 27772
rect 113000 27770 113056 27772
rect 113080 27770 113136 27772
rect 113160 27770 113216 27772
rect 112920 27718 112966 27770
rect 112966 27718 112976 27770
rect 113000 27718 113030 27770
rect 113030 27718 113042 27770
rect 113042 27718 113056 27770
rect 113080 27718 113094 27770
rect 113094 27718 113106 27770
rect 113106 27718 113136 27770
rect 113160 27718 113170 27770
rect 113170 27718 113216 27770
rect 112920 27716 112976 27718
rect 113000 27716 113056 27718
rect 113080 27716 113136 27718
rect 113160 27716 113216 27718
rect 113656 27226 113712 27228
rect 113736 27226 113792 27228
rect 113816 27226 113872 27228
rect 113896 27226 113952 27228
rect 113656 27174 113702 27226
rect 113702 27174 113712 27226
rect 113736 27174 113766 27226
rect 113766 27174 113778 27226
rect 113778 27174 113792 27226
rect 113816 27174 113830 27226
rect 113830 27174 113842 27226
rect 113842 27174 113872 27226
rect 113896 27174 113906 27226
rect 113906 27174 113952 27226
rect 113656 27172 113712 27174
rect 113736 27172 113792 27174
rect 113816 27172 113872 27174
rect 113896 27172 113952 27174
rect 115294 32836 115350 32872
rect 115294 32816 115296 32836
rect 115296 32816 115348 32836
rect 115348 32816 115350 32836
rect 115846 33496 115902 33552
rect 116122 33940 116124 33960
rect 116124 33940 116176 33960
rect 116176 33940 116178 33960
rect 116122 33904 116178 33940
rect 116214 33532 116216 33552
rect 116216 33532 116268 33552
rect 116268 33532 116270 33552
rect 116214 33496 116270 33532
rect 115754 31864 115810 31920
rect 115110 30812 115112 30832
rect 115112 30812 115164 30832
rect 115164 30812 115166 30832
rect 115110 30776 115166 30812
rect 116122 31728 116178 31784
rect 116490 32816 116546 32872
rect 116766 32428 116822 32464
rect 116766 32408 116768 32428
rect 116768 32408 116820 32428
rect 116820 32408 116822 32428
rect 116582 32308 116584 32328
rect 116584 32308 116636 32328
rect 116636 32308 116638 32328
rect 116582 32272 116638 32308
rect 112920 26682 112976 26684
rect 113000 26682 113056 26684
rect 113080 26682 113136 26684
rect 113160 26682 113216 26684
rect 112920 26630 112966 26682
rect 112966 26630 112976 26682
rect 113000 26630 113030 26682
rect 113030 26630 113042 26682
rect 113042 26630 113056 26682
rect 113080 26630 113094 26682
rect 113094 26630 113106 26682
rect 113106 26630 113136 26682
rect 113160 26630 113170 26682
rect 113170 26630 113216 26682
rect 112920 26628 112976 26630
rect 113000 26628 113056 26630
rect 113080 26628 113136 26630
rect 113160 26628 113216 26630
rect 117134 31728 117190 31784
rect 117318 32428 117374 32464
rect 117318 32408 117320 32428
rect 117320 32408 117372 32428
rect 117372 32408 117374 32428
rect 117502 32272 117558 32328
rect 118514 32000 118570 32056
rect 118514 31340 118570 31376
rect 118514 31320 118516 31340
rect 118516 31320 118568 31340
rect 118568 31320 118570 31340
rect 118514 30640 118570 30696
rect 117318 28600 117374 28656
rect 118238 29280 118294 29336
rect 118238 27920 118294 27976
rect 118606 29960 118662 30016
rect 118514 28600 118570 28656
rect 118514 27240 118570 27296
rect 113656 26138 113712 26140
rect 113736 26138 113792 26140
rect 113816 26138 113872 26140
rect 113896 26138 113952 26140
rect 113656 26086 113702 26138
rect 113702 26086 113712 26138
rect 113736 26086 113766 26138
rect 113766 26086 113778 26138
rect 113778 26086 113792 26138
rect 113816 26086 113830 26138
rect 113830 26086 113842 26138
rect 113842 26086 113872 26138
rect 113896 26086 113906 26138
rect 113906 26086 113952 26138
rect 113656 26084 113712 26086
rect 113736 26084 113792 26086
rect 113816 26084 113872 26086
rect 113896 26084 113952 26086
rect 112920 25594 112976 25596
rect 113000 25594 113056 25596
rect 113080 25594 113136 25596
rect 113160 25594 113216 25596
rect 112920 25542 112966 25594
rect 112966 25542 112976 25594
rect 113000 25542 113030 25594
rect 113030 25542 113042 25594
rect 113042 25542 113056 25594
rect 113080 25542 113094 25594
rect 113094 25542 113106 25594
rect 113106 25542 113136 25594
rect 113160 25542 113170 25594
rect 113170 25542 113216 25594
rect 112920 25540 112976 25542
rect 113000 25540 113056 25542
rect 113080 25540 113136 25542
rect 113160 25540 113216 25542
rect 113656 25050 113712 25052
rect 113736 25050 113792 25052
rect 113816 25050 113872 25052
rect 113896 25050 113952 25052
rect 113656 24998 113702 25050
rect 113702 24998 113712 25050
rect 113736 24998 113766 25050
rect 113766 24998 113778 25050
rect 113778 24998 113792 25050
rect 113816 24998 113830 25050
rect 113830 24998 113842 25050
rect 113842 24998 113872 25050
rect 113896 24998 113906 25050
rect 113906 24998 113952 25050
rect 113656 24996 113712 24998
rect 113736 24996 113792 24998
rect 113816 24996 113872 24998
rect 113896 24996 113952 24998
rect 112920 24506 112976 24508
rect 113000 24506 113056 24508
rect 113080 24506 113136 24508
rect 113160 24506 113216 24508
rect 112920 24454 112966 24506
rect 112966 24454 112976 24506
rect 113000 24454 113030 24506
rect 113030 24454 113042 24506
rect 113042 24454 113056 24506
rect 113080 24454 113094 24506
rect 113094 24454 113106 24506
rect 113106 24454 113136 24506
rect 113160 24454 113170 24506
rect 113170 24454 113216 24506
rect 112920 24452 112976 24454
rect 113000 24452 113056 24454
rect 113080 24452 113136 24454
rect 113160 24452 113216 24454
rect 113656 23962 113712 23964
rect 113736 23962 113792 23964
rect 113816 23962 113872 23964
rect 113896 23962 113952 23964
rect 113656 23910 113702 23962
rect 113702 23910 113712 23962
rect 113736 23910 113766 23962
rect 113766 23910 113778 23962
rect 113778 23910 113792 23962
rect 113816 23910 113830 23962
rect 113830 23910 113842 23962
rect 113842 23910 113872 23962
rect 113896 23910 113906 23962
rect 113906 23910 113952 23962
rect 113656 23908 113712 23910
rect 113736 23908 113792 23910
rect 113816 23908 113872 23910
rect 113896 23908 113952 23910
rect 112920 23418 112976 23420
rect 113000 23418 113056 23420
rect 113080 23418 113136 23420
rect 113160 23418 113216 23420
rect 112920 23366 112966 23418
rect 112966 23366 112976 23418
rect 113000 23366 113030 23418
rect 113030 23366 113042 23418
rect 113042 23366 113056 23418
rect 113080 23366 113094 23418
rect 113094 23366 113106 23418
rect 113106 23366 113136 23418
rect 113160 23366 113170 23418
rect 113170 23366 113216 23418
rect 112920 23364 112976 23366
rect 113000 23364 113056 23366
rect 113080 23364 113136 23366
rect 113160 23364 113216 23366
rect 113656 22874 113712 22876
rect 113736 22874 113792 22876
rect 113816 22874 113872 22876
rect 113896 22874 113952 22876
rect 113656 22822 113702 22874
rect 113702 22822 113712 22874
rect 113736 22822 113766 22874
rect 113766 22822 113778 22874
rect 113778 22822 113792 22874
rect 113816 22822 113830 22874
rect 113830 22822 113842 22874
rect 113842 22822 113872 22874
rect 113896 22822 113906 22874
rect 113906 22822 113952 22874
rect 113656 22820 113712 22822
rect 113736 22820 113792 22822
rect 113816 22820 113872 22822
rect 113896 22820 113952 22822
rect 112920 22330 112976 22332
rect 113000 22330 113056 22332
rect 113080 22330 113136 22332
rect 113160 22330 113216 22332
rect 112920 22278 112966 22330
rect 112966 22278 112976 22330
rect 113000 22278 113030 22330
rect 113030 22278 113042 22330
rect 113042 22278 113056 22330
rect 113080 22278 113094 22330
rect 113094 22278 113106 22330
rect 113106 22278 113136 22330
rect 113160 22278 113170 22330
rect 113170 22278 113216 22330
rect 112920 22276 112976 22278
rect 113000 22276 113056 22278
rect 113080 22276 113136 22278
rect 113160 22276 113216 22278
rect 113656 21786 113712 21788
rect 113736 21786 113792 21788
rect 113816 21786 113872 21788
rect 113896 21786 113952 21788
rect 113656 21734 113702 21786
rect 113702 21734 113712 21786
rect 113736 21734 113766 21786
rect 113766 21734 113778 21786
rect 113778 21734 113792 21786
rect 113816 21734 113830 21786
rect 113830 21734 113842 21786
rect 113842 21734 113872 21786
rect 113896 21734 113906 21786
rect 113906 21734 113952 21786
rect 113656 21732 113712 21734
rect 113736 21732 113792 21734
rect 113816 21732 113872 21734
rect 113896 21732 113952 21734
rect 112920 21242 112976 21244
rect 113000 21242 113056 21244
rect 113080 21242 113136 21244
rect 113160 21242 113216 21244
rect 112920 21190 112966 21242
rect 112966 21190 112976 21242
rect 113000 21190 113030 21242
rect 113030 21190 113042 21242
rect 113042 21190 113056 21242
rect 113080 21190 113094 21242
rect 113094 21190 113106 21242
rect 113106 21190 113136 21242
rect 113160 21190 113170 21242
rect 113170 21190 113216 21242
rect 112920 21188 112976 21190
rect 113000 21188 113056 21190
rect 113080 21188 113136 21190
rect 113160 21188 113216 21190
rect 113656 20698 113712 20700
rect 113736 20698 113792 20700
rect 113816 20698 113872 20700
rect 113896 20698 113952 20700
rect 113656 20646 113702 20698
rect 113702 20646 113712 20698
rect 113736 20646 113766 20698
rect 113766 20646 113778 20698
rect 113778 20646 113792 20698
rect 113816 20646 113830 20698
rect 113830 20646 113842 20698
rect 113842 20646 113872 20698
rect 113896 20646 113906 20698
rect 113906 20646 113952 20698
rect 113656 20644 113712 20646
rect 113736 20644 113792 20646
rect 113816 20644 113872 20646
rect 113896 20644 113952 20646
rect 112920 20154 112976 20156
rect 113000 20154 113056 20156
rect 113080 20154 113136 20156
rect 113160 20154 113216 20156
rect 112920 20102 112966 20154
rect 112966 20102 112976 20154
rect 113000 20102 113030 20154
rect 113030 20102 113042 20154
rect 113042 20102 113056 20154
rect 113080 20102 113094 20154
rect 113094 20102 113106 20154
rect 113106 20102 113136 20154
rect 113160 20102 113170 20154
rect 113170 20102 113216 20154
rect 112920 20100 112976 20102
rect 113000 20100 113056 20102
rect 113080 20100 113136 20102
rect 113160 20100 113216 20102
rect 113656 19610 113712 19612
rect 113736 19610 113792 19612
rect 113816 19610 113872 19612
rect 113896 19610 113952 19612
rect 113656 19558 113702 19610
rect 113702 19558 113712 19610
rect 113736 19558 113766 19610
rect 113766 19558 113778 19610
rect 113778 19558 113792 19610
rect 113816 19558 113830 19610
rect 113830 19558 113842 19610
rect 113842 19558 113872 19610
rect 113896 19558 113906 19610
rect 113906 19558 113952 19610
rect 113656 19556 113712 19558
rect 113736 19556 113792 19558
rect 113816 19556 113872 19558
rect 113896 19556 113952 19558
rect 112920 19066 112976 19068
rect 113000 19066 113056 19068
rect 113080 19066 113136 19068
rect 113160 19066 113216 19068
rect 112920 19014 112966 19066
rect 112966 19014 112976 19066
rect 113000 19014 113030 19066
rect 113030 19014 113042 19066
rect 113042 19014 113056 19066
rect 113080 19014 113094 19066
rect 113094 19014 113106 19066
rect 113106 19014 113136 19066
rect 113160 19014 113170 19066
rect 113170 19014 113216 19066
rect 112920 19012 112976 19014
rect 113000 19012 113056 19014
rect 113080 19012 113136 19014
rect 113160 19012 113216 19014
rect 113656 18522 113712 18524
rect 113736 18522 113792 18524
rect 113816 18522 113872 18524
rect 113896 18522 113952 18524
rect 113656 18470 113702 18522
rect 113702 18470 113712 18522
rect 113736 18470 113766 18522
rect 113766 18470 113778 18522
rect 113778 18470 113792 18522
rect 113816 18470 113830 18522
rect 113830 18470 113842 18522
rect 113842 18470 113872 18522
rect 113896 18470 113906 18522
rect 113906 18470 113952 18522
rect 113656 18468 113712 18470
rect 113736 18468 113792 18470
rect 113816 18468 113872 18470
rect 113896 18468 113952 18470
rect 112920 17978 112976 17980
rect 113000 17978 113056 17980
rect 113080 17978 113136 17980
rect 113160 17978 113216 17980
rect 112920 17926 112966 17978
rect 112966 17926 112976 17978
rect 113000 17926 113030 17978
rect 113030 17926 113042 17978
rect 113042 17926 113056 17978
rect 113080 17926 113094 17978
rect 113094 17926 113106 17978
rect 113106 17926 113136 17978
rect 113160 17926 113170 17978
rect 113170 17926 113216 17978
rect 112920 17924 112976 17926
rect 113000 17924 113056 17926
rect 113080 17924 113136 17926
rect 113160 17924 113216 17926
rect 113656 17434 113712 17436
rect 113736 17434 113792 17436
rect 113816 17434 113872 17436
rect 113896 17434 113952 17436
rect 113656 17382 113702 17434
rect 113702 17382 113712 17434
rect 113736 17382 113766 17434
rect 113766 17382 113778 17434
rect 113778 17382 113792 17434
rect 113816 17382 113830 17434
rect 113830 17382 113842 17434
rect 113842 17382 113872 17434
rect 113896 17382 113906 17434
rect 113906 17382 113952 17434
rect 113656 17380 113712 17382
rect 113736 17380 113792 17382
rect 113816 17380 113872 17382
rect 113896 17380 113952 17382
rect 112920 16890 112976 16892
rect 113000 16890 113056 16892
rect 113080 16890 113136 16892
rect 113160 16890 113216 16892
rect 112920 16838 112966 16890
rect 112966 16838 112976 16890
rect 113000 16838 113030 16890
rect 113030 16838 113042 16890
rect 113042 16838 113056 16890
rect 113080 16838 113094 16890
rect 113094 16838 113106 16890
rect 113106 16838 113136 16890
rect 113160 16838 113170 16890
rect 113170 16838 113216 16890
rect 112920 16836 112976 16838
rect 113000 16836 113056 16838
rect 113080 16836 113136 16838
rect 113160 16836 113216 16838
rect 113656 16346 113712 16348
rect 113736 16346 113792 16348
rect 113816 16346 113872 16348
rect 113896 16346 113952 16348
rect 113656 16294 113702 16346
rect 113702 16294 113712 16346
rect 113736 16294 113766 16346
rect 113766 16294 113778 16346
rect 113778 16294 113792 16346
rect 113816 16294 113830 16346
rect 113830 16294 113842 16346
rect 113842 16294 113872 16346
rect 113896 16294 113906 16346
rect 113906 16294 113952 16346
rect 113656 16292 113712 16294
rect 113736 16292 113792 16294
rect 113816 16292 113872 16294
rect 113896 16292 113952 16294
rect 112920 15802 112976 15804
rect 113000 15802 113056 15804
rect 113080 15802 113136 15804
rect 113160 15802 113216 15804
rect 112920 15750 112966 15802
rect 112966 15750 112976 15802
rect 113000 15750 113030 15802
rect 113030 15750 113042 15802
rect 113042 15750 113056 15802
rect 113080 15750 113094 15802
rect 113094 15750 113106 15802
rect 113106 15750 113136 15802
rect 113160 15750 113170 15802
rect 113170 15750 113216 15802
rect 112920 15748 112976 15750
rect 113000 15748 113056 15750
rect 113080 15748 113136 15750
rect 113160 15748 113216 15750
rect 113656 15258 113712 15260
rect 113736 15258 113792 15260
rect 113816 15258 113872 15260
rect 113896 15258 113952 15260
rect 113656 15206 113702 15258
rect 113702 15206 113712 15258
rect 113736 15206 113766 15258
rect 113766 15206 113778 15258
rect 113778 15206 113792 15258
rect 113816 15206 113830 15258
rect 113830 15206 113842 15258
rect 113842 15206 113872 15258
rect 113896 15206 113906 15258
rect 113906 15206 113952 15258
rect 113656 15204 113712 15206
rect 113736 15204 113792 15206
rect 113816 15204 113872 15206
rect 113896 15204 113952 15206
rect 112920 14714 112976 14716
rect 113000 14714 113056 14716
rect 113080 14714 113136 14716
rect 113160 14714 113216 14716
rect 112920 14662 112966 14714
rect 112966 14662 112976 14714
rect 113000 14662 113030 14714
rect 113030 14662 113042 14714
rect 113042 14662 113056 14714
rect 113080 14662 113094 14714
rect 113094 14662 113106 14714
rect 113106 14662 113136 14714
rect 113160 14662 113170 14714
rect 113170 14662 113216 14714
rect 112920 14660 112976 14662
rect 113000 14660 113056 14662
rect 113080 14660 113136 14662
rect 113160 14660 113216 14662
rect 113656 14170 113712 14172
rect 113736 14170 113792 14172
rect 113816 14170 113872 14172
rect 113896 14170 113952 14172
rect 113656 14118 113702 14170
rect 113702 14118 113712 14170
rect 113736 14118 113766 14170
rect 113766 14118 113778 14170
rect 113778 14118 113792 14170
rect 113816 14118 113830 14170
rect 113830 14118 113842 14170
rect 113842 14118 113872 14170
rect 113896 14118 113906 14170
rect 113906 14118 113952 14170
rect 113656 14116 113712 14118
rect 113736 14116 113792 14118
rect 113816 14116 113872 14118
rect 113896 14116 113952 14118
rect 112920 13626 112976 13628
rect 113000 13626 113056 13628
rect 113080 13626 113136 13628
rect 113160 13626 113216 13628
rect 112920 13574 112966 13626
rect 112966 13574 112976 13626
rect 113000 13574 113030 13626
rect 113030 13574 113042 13626
rect 113042 13574 113056 13626
rect 113080 13574 113094 13626
rect 113094 13574 113106 13626
rect 113106 13574 113136 13626
rect 113160 13574 113170 13626
rect 113170 13574 113216 13626
rect 112920 13572 112976 13574
rect 113000 13572 113056 13574
rect 113080 13572 113136 13574
rect 113160 13572 113216 13574
rect 113656 13082 113712 13084
rect 113736 13082 113792 13084
rect 113816 13082 113872 13084
rect 113896 13082 113952 13084
rect 113656 13030 113702 13082
rect 113702 13030 113712 13082
rect 113736 13030 113766 13082
rect 113766 13030 113778 13082
rect 113778 13030 113792 13082
rect 113816 13030 113830 13082
rect 113830 13030 113842 13082
rect 113842 13030 113872 13082
rect 113896 13030 113906 13082
rect 113906 13030 113952 13082
rect 113656 13028 113712 13030
rect 113736 13028 113792 13030
rect 113816 13028 113872 13030
rect 113896 13028 113952 13030
rect 112920 12538 112976 12540
rect 113000 12538 113056 12540
rect 113080 12538 113136 12540
rect 113160 12538 113216 12540
rect 112920 12486 112966 12538
rect 112966 12486 112976 12538
rect 113000 12486 113030 12538
rect 113030 12486 113042 12538
rect 113042 12486 113056 12538
rect 113080 12486 113094 12538
rect 113094 12486 113106 12538
rect 113106 12486 113136 12538
rect 113160 12486 113170 12538
rect 113170 12486 113216 12538
rect 112920 12484 112976 12486
rect 113000 12484 113056 12486
rect 113080 12484 113136 12486
rect 113160 12484 113216 12486
rect 113656 11994 113712 11996
rect 113736 11994 113792 11996
rect 113816 11994 113872 11996
rect 113896 11994 113952 11996
rect 113656 11942 113702 11994
rect 113702 11942 113712 11994
rect 113736 11942 113766 11994
rect 113766 11942 113778 11994
rect 113778 11942 113792 11994
rect 113816 11942 113830 11994
rect 113830 11942 113842 11994
rect 113842 11942 113872 11994
rect 113896 11942 113906 11994
rect 113906 11942 113952 11994
rect 113656 11940 113712 11942
rect 113736 11940 113792 11942
rect 113816 11940 113872 11942
rect 113896 11940 113952 11942
rect 112920 11450 112976 11452
rect 113000 11450 113056 11452
rect 113080 11450 113136 11452
rect 113160 11450 113216 11452
rect 112920 11398 112966 11450
rect 112966 11398 112976 11450
rect 113000 11398 113030 11450
rect 113030 11398 113042 11450
rect 113042 11398 113056 11450
rect 113080 11398 113094 11450
rect 113094 11398 113106 11450
rect 113106 11398 113136 11450
rect 113160 11398 113170 11450
rect 113170 11398 113216 11450
rect 112920 11396 112976 11398
rect 113000 11396 113056 11398
rect 113080 11396 113136 11398
rect 113160 11396 113216 11398
rect 113656 10906 113712 10908
rect 113736 10906 113792 10908
rect 113816 10906 113872 10908
rect 113896 10906 113952 10908
rect 113656 10854 113702 10906
rect 113702 10854 113712 10906
rect 113736 10854 113766 10906
rect 113766 10854 113778 10906
rect 113778 10854 113792 10906
rect 113816 10854 113830 10906
rect 113830 10854 113842 10906
rect 113842 10854 113872 10906
rect 113896 10854 113906 10906
rect 113906 10854 113952 10906
rect 113656 10852 113712 10854
rect 113736 10852 113792 10854
rect 113816 10852 113872 10854
rect 113896 10852 113952 10854
rect 112920 10362 112976 10364
rect 113000 10362 113056 10364
rect 113080 10362 113136 10364
rect 113160 10362 113216 10364
rect 112920 10310 112966 10362
rect 112966 10310 112976 10362
rect 113000 10310 113030 10362
rect 113030 10310 113042 10362
rect 113042 10310 113056 10362
rect 113080 10310 113094 10362
rect 113094 10310 113106 10362
rect 113106 10310 113136 10362
rect 113160 10310 113170 10362
rect 113170 10310 113216 10362
rect 112920 10308 112976 10310
rect 113000 10308 113056 10310
rect 113080 10308 113136 10310
rect 113160 10308 113216 10310
rect 108762 9968 108818 10024
rect 26974 9696 27030 9752
rect 27802 9696 27858 9752
rect 29550 9696 29606 9752
rect 30194 9696 30250 9752
rect 51630 9696 51686 9752
rect 52458 9696 52514 9752
rect 53562 9696 53618 9752
rect 55034 9696 55090 9752
rect 56138 9696 56194 9752
rect 57426 9696 57482 9752
rect 58254 9696 58310 9752
rect 59542 9696 59598 9752
rect 60830 9696 60886 9752
rect 67730 9696 67786 9752
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 25870 8200 25926 8256
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 31666 8200 31722 8256
rect 32954 8200 33010 8256
rect 33782 8200 33838 8256
rect 34794 8200 34850 8256
rect 36174 8200 36230 8256
rect 37462 8200 37518 8256
rect 38290 8200 38346 8256
rect 40866 8200 40922 8256
rect 41970 8200 42026 8256
rect 43258 8200 43314 8256
rect 44546 8200 44602 8256
rect 46662 8200 46718 8256
rect 47766 8200 47822 8256
rect 49054 8200 49110 8256
rect 50342 8200 50398 8256
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 40038 2644 40094 2680
rect 45834 7112 45890 7168
rect 61934 8200 61990 8256
rect 63222 8200 63278 8256
rect 64050 8200 64106 8256
rect 65338 8200 65394 8256
rect 66718 8200 66774 8256
rect 66320 7642 66376 7644
rect 66400 7642 66456 7644
rect 66480 7642 66536 7644
rect 66560 7642 66616 7644
rect 66320 7590 66366 7642
rect 66366 7590 66376 7642
rect 66400 7590 66430 7642
rect 66430 7590 66442 7642
rect 66442 7590 66456 7642
rect 66480 7590 66494 7642
rect 66494 7590 66506 7642
rect 66506 7590 66536 7642
rect 66560 7590 66570 7642
rect 66570 7590 66616 7642
rect 66320 7588 66376 7590
rect 66400 7588 66456 7590
rect 66480 7588 66536 7590
rect 66560 7588 66616 7590
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 66320 6554 66376 6556
rect 66400 6554 66456 6556
rect 66480 6554 66536 6556
rect 66560 6554 66616 6556
rect 66320 6502 66366 6554
rect 66366 6502 66376 6554
rect 66400 6502 66430 6554
rect 66430 6502 66442 6554
rect 66442 6502 66456 6554
rect 66480 6502 66494 6554
rect 66494 6502 66506 6554
rect 66506 6502 66536 6554
rect 66560 6502 66570 6554
rect 66570 6502 66616 6554
rect 66320 6500 66376 6502
rect 66400 6500 66456 6502
rect 66480 6500 66536 6502
rect 66560 6500 66616 6502
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 66320 5466 66376 5468
rect 66400 5466 66456 5468
rect 66480 5466 66536 5468
rect 66560 5466 66616 5468
rect 66320 5414 66366 5466
rect 66366 5414 66376 5466
rect 66400 5414 66430 5466
rect 66430 5414 66442 5466
rect 66442 5414 66456 5466
rect 66480 5414 66494 5466
rect 66494 5414 66506 5466
rect 66506 5414 66536 5466
rect 66560 5414 66570 5466
rect 66570 5414 66616 5466
rect 66320 5412 66376 5414
rect 66400 5412 66456 5414
rect 66480 5412 66536 5414
rect 66560 5412 66616 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 66320 4378 66376 4380
rect 66400 4378 66456 4380
rect 66480 4378 66536 4380
rect 66560 4378 66616 4380
rect 66320 4326 66366 4378
rect 66366 4326 66376 4378
rect 66400 4326 66430 4378
rect 66430 4326 66442 4378
rect 66442 4326 66456 4378
rect 66480 4326 66494 4378
rect 66494 4326 66506 4378
rect 66506 4326 66536 4378
rect 66560 4326 66570 4378
rect 66570 4326 66616 4378
rect 66320 4324 66376 4326
rect 66400 4324 66456 4326
rect 66480 4324 66536 4326
rect 66560 4324 66616 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 66320 3290 66376 3292
rect 66400 3290 66456 3292
rect 66480 3290 66536 3292
rect 66560 3290 66616 3292
rect 66320 3238 66366 3290
rect 66366 3238 66376 3290
rect 66400 3238 66430 3290
rect 66430 3238 66442 3290
rect 66442 3238 66456 3290
rect 66480 3238 66494 3290
rect 66494 3238 66506 3290
rect 66506 3238 66536 3290
rect 66560 3238 66570 3290
rect 66570 3238 66616 3290
rect 66320 3236 66376 3238
rect 66400 3236 66456 3238
rect 66480 3236 66536 3238
rect 66560 3236 66616 3238
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 93398 9832 93454 9888
rect 93030 9696 93086 9752
rect 93214 8200 93270 8256
rect 113656 9818 113712 9820
rect 113736 9818 113792 9820
rect 113816 9818 113872 9820
rect 113896 9818 113952 9820
rect 113656 9766 113702 9818
rect 113702 9766 113712 9818
rect 113736 9766 113766 9818
rect 113766 9766 113778 9818
rect 113778 9766 113792 9818
rect 113816 9766 113830 9818
rect 113830 9766 113842 9818
rect 113842 9766 113872 9818
rect 113896 9766 113906 9818
rect 113906 9766 113952 9818
rect 113656 9764 113712 9766
rect 113736 9764 113792 9766
rect 113816 9764 113872 9766
rect 113896 9764 113952 9766
rect 112920 9274 112976 9276
rect 113000 9274 113056 9276
rect 113080 9274 113136 9276
rect 113160 9274 113216 9276
rect 112920 9222 112966 9274
rect 112966 9222 112976 9274
rect 113000 9222 113030 9274
rect 113030 9222 113042 9274
rect 113042 9222 113056 9274
rect 113080 9222 113094 9274
rect 113094 9222 113106 9274
rect 113106 9222 113136 9274
rect 113160 9222 113170 9274
rect 113170 9222 113216 9274
rect 112920 9220 112976 9222
rect 113000 9220 113056 9222
rect 113080 9220 113136 9222
rect 113160 9220 113216 9222
rect 113656 8730 113712 8732
rect 113736 8730 113792 8732
rect 113816 8730 113872 8732
rect 113896 8730 113952 8732
rect 113656 8678 113702 8730
rect 113702 8678 113712 8730
rect 113736 8678 113766 8730
rect 113766 8678 113778 8730
rect 113778 8678 113792 8730
rect 113816 8678 113830 8730
rect 113830 8678 113842 8730
rect 113842 8678 113872 8730
rect 113896 8678 113906 8730
rect 113906 8678 113952 8730
rect 113656 8676 113712 8678
rect 113736 8676 113792 8678
rect 113816 8676 113872 8678
rect 113896 8676 113952 8678
rect 112920 8186 112976 8188
rect 113000 8186 113056 8188
rect 113080 8186 113136 8188
rect 113160 8186 113216 8188
rect 112920 8134 112966 8186
rect 112966 8134 112976 8186
rect 113000 8134 113030 8186
rect 113030 8134 113042 8186
rect 113042 8134 113056 8186
rect 113080 8134 113094 8186
rect 113094 8134 113106 8186
rect 113106 8134 113136 8186
rect 113160 8134 113170 8186
rect 113170 8134 113216 8186
rect 112920 8132 112976 8134
rect 113000 8132 113056 8134
rect 113080 8132 113136 8134
rect 113160 8132 113216 8134
rect 97040 7642 97096 7644
rect 97120 7642 97176 7644
rect 97200 7642 97256 7644
rect 97280 7642 97336 7644
rect 97040 7590 97086 7642
rect 97086 7590 97096 7642
rect 97120 7590 97150 7642
rect 97150 7590 97162 7642
rect 97162 7590 97176 7642
rect 97200 7590 97214 7642
rect 97214 7590 97226 7642
rect 97226 7590 97256 7642
rect 97280 7590 97290 7642
rect 97290 7590 97336 7642
rect 97040 7588 97096 7590
rect 97120 7588 97176 7590
rect 97200 7588 97256 7590
rect 97280 7588 97336 7590
rect 113656 7642 113712 7644
rect 113736 7642 113792 7644
rect 113816 7642 113872 7644
rect 113896 7642 113952 7644
rect 113656 7590 113702 7642
rect 113702 7590 113712 7642
rect 113736 7590 113766 7642
rect 113766 7590 113778 7642
rect 113778 7590 113792 7642
rect 113816 7590 113830 7642
rect 113830 7590 113842 7642
rect 113842 7590 113872 7642
rect 113896 7590 113906 7642
rect 113906 7590 113952 7642
rect 113656 7588 113712 7590
rect 113736 7588 113792 7590
rect 113816 7588 113872 7590
rect 113896 7588 113952 7590
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 112920 7098 112976 7100
rect 113000 7098 113056 7100
rect 113080 7098 113136 7100
rect 113160 7098 113216 7100
rect 112920 7046 112966 7098
rect 112966 7046 112976 7098
rect 113000 7046 113030 7098
rect 113030 7046 113042 7098
rect 113042 7046 113056 7098
rect 113080 7046 113094 7098
rect 113094 7046 113106 7098
rect 113106 7046 113136 7098
rect 113160 7046 113170 7098
rect 113170 7046 113216 7098
rect 112920 7044 112976 7046
rect 113000 7044 113056 7046
rect 113080 7044 113136 7046
rect 113160 7044 113216 7046
rect 97040 6554 97096 6556
rect 97120 6554 97176 6556
rect 97200 6554 97256 6556
rect 97280 6554 97336 6556
rect 97040 6502 97086 6554
rect 97086 6502 97096 6554
rect 97120 6502 97150 6554
rect 97150 6502 97162 6554
rect 97162 6502 97176 6554
rect 97200 6502 97214 6554
rect 97214 6502 97226 6554
rect 97226 6502 97256 6554
rect 97280 6502 97290 6554
rect 97290 6502 97336 6554
rect 97040 6500 97096 6502
rect 97120 6500 97176 6502
rect 97200 6500 97256 6502
rect 97280 6500 97336 6502
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 97040 5466 97096 5468
rect 97120 5466 97176 5468
rect 97200 5466 97256 5468
rect 97280 5466 97336 5468
rect 97040 5414 97086 5466
rect 97086 5414 97096 5466
rect 97120 5414 97150 5466
rect 97150 5414 97162 5466
rect 97162 5414 97176 5466
rect 97200 5414 97214 5466
rect 97214 5414 97226 5466
rect 97226 5414 97256 5466
rect 97280 5414 97290 5466
rect 97290 5414 97336 5466
rect 97040 5412 97096 5414
rect 97120 5412 97176 5414
rect 97200 5412 97256 5414
rect 97280 5412 97336 5414
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 97040 4378 97096 4380
rect 97120 4378 97176 4380
rect 97200 4378 97256 4380
rect 97280 4378 97336 4380
rect 97040 4326 97086 4378
rect 97086 4326 97096 4378
rect 97120 4326 97150 4378
rect 97150 4326 97162 4378
rect 97162 4326 97176 4378
rect 97200 4326 97214 4378
rect 97214 4326 97226 4378
rect 97226 4326 97256 4378
rect 97280 4326 97290 4378
rect 97290 4326 97336 4378
rect 97040 4324 97096 4326
rect 97120 4324 97176 4326
rect 97200 4324 97256 4326
rect 97280 4324 97336 4326
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 97040 3290 97096 3292
rect 97120 3290 97176 3292
rect 97200 3290 97256 3292
rect 97280 3290 97336 3292
rect 97040 3238 97086 3290
rect 97086 3238 97096 3290
rect 97120 3238 97150 3290
rect 97150 3238 97162 3290
rect 97162 3238 97176 3290
rect 97200 3238 97214 3290
rect 97214 3238 97226 3290
rect 97226 3238 97256 3290
rect 97280 3238 97290 3290
rect 97290 3238 97336 3290
rect 97040 3236 97096 3238
rect 97120 3236 97176 3238
rect 97200 3236 97256 3238
rect 97280 3236 97336 3238
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 40038 2624 40040 2644
rect 40040 2624 40092 2644
rect 40092 2624 40094 2644
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 66320 2202 66376 2204
rect 66400 2202 66456 2204
rect 66480 2202 66536 2204
rect 66560 2202 66616 2204
rect 66320 2150 66366 2202
rect 66366 2150 66376 2202
rect 66400 2150 66430 2202
rect 66430 2150 66442 2202
rect 66442 2150 66456 2202
rect 66480 2150 66494 2202
rect 66494 2150 66506 2202
rect 66506 2150 66536 2202
rect 66560 2150 66570 2202
rect 66570 2150 66616 2202
rect 66320 2148 66376 2150
rect 66400 2148 66456 2150
rect 66480 2148 66536 2150
rect 66560 2148 66616 2150
rect 97040 2202 97096 2204
rect 97120 2202 97176 2204
rect 97200 2202 97256 2204
rect 97280 2202 97336 2204
rect 97040 2150 97086 2202
rect 97086 2150 97096 2202
rect 97120 2150 97150 2202
rect 97150 2150 97162 2202
rect 97162 2150 97176 2202
rect 97200 2150 97214 2202
rect 97214 2150 97226 2202
rect 97226 2150 97256 2202
rect 97280 2150 97290 2202
rect 97290 2150 97336 2202
rect 97040 2148 97096 2150
rect 97120 2148 97176 2150
rect 97200 2148 97256 2150
rect 97280 2148 97336 2150
<< metal3 >>
rect 4210 97408 4526 97409
rect 4210 97344 4216 97408
rect 4280 97344 4296 97408
rect 4360 97344 4376 97408
rect 4440 97344 4456 97408
rect 4520 97344 4526 97408
rect 4210 97343 4526 97344
rect 34930 97408 35246 97409
rect 34930 97344 34936 97408
rect 35000 97344 35016 97408
rect 35080 97344 35096 97408
rect 35160 97344 35176 97408
rect 35240 97344 35246 97408
rect 34930 97343 35246 97344
rect 65650 97408 65966 97409
rect 65650 97344 65656 97408
rect 65720 97344 65736 97408
rect 65800 97344 65816 97408
rect 65880 97344 65896 97408
rect 65960 97344 65966 97408
rect 65650 97343 65966 97344
rect 96370 97408 96686 97409
rect 96370 97344 96376 97408
rect 96440 97344 96456 97408
rect 96520 97344 96536 97408
rect 96600 97344 96616 97408
rect 96680 97344 96686 97408
rect 96370 97343 96686 97344
rect 4870 96864 5186 96865
rect 4870 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5186 96864
rect 4870 96799 5186 96800
rect 35590 96864 35906 96865
rect 35590 96800 35596 96864
rect 35660 96800 35676 96864
rect 35740 96800 35756 96864
rect 35820 96800 35836 96864
rect 35900 96800 35906 96864
rect 35590 96799 35906 96800
rect 66310 96864 66626 96865
rect 66310 96800 66316 96864
rect 66380 96800 66396 96864
rect 66460 96800 66476 96864
rect 66540 96800 66556 96864
rect 66620 96800 66626 96864
rect 66310 96799 66626 96800
rect 97030 96864 97346 96865
rect 97030 96800 97036 96864
rect 97100 96800 97116 96864
rect 97180 96800 97196 96864
rect 97260 96800 97276 96864
rect 97340 96800 97346 96864
rect 97030 96799 97346 96800
rect 4210 96320 4526 96321
rect 4210 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4526 96320
rect 4210 96255 4526 96256
rect 34930 96320 35246 96321
rect 34930 96256 34936 96320
rect 35000 96256 35016 96320
rect 35080 96256 35096 96320
rect 35160 96256 35176 96320
rect 35240 96256 35246 96320
rect 34930 96255 35246 96256
rect 65650 96320 65966 96321
rect 65650 96256 65656 96320
rect 65720 96256 65736 96320
rect 65800 96256 65816 96320
rect 65880 96256 65896 96320
rect 65960 96256 65966 96320
rect 65650 96255 65966 96256
rect 96370 96320 96686 96321
rect 96370 96256 96376 96320
rect 96440 96256 96456 96320
rect 96520 96256 96536 96320
rect 96600 96256 96616 96320
rect 96680 96256 96686 96320
rect 96370 96255 96686 96256
rect 4870 95776 5186 95777
rect 4870 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5186 95776
rect 4870 95711 5186 95712
rect 35590 95776 35906 95777
rect 35590 95712 35596 95776
rect 35660 95712 35676 95776
rect 35740 95712 35756 95776
rect 35820 95712 35836 95776
rect 35900 95712 35906 95776
rect 35590 95711 35906 95712
rect 66310 95776 66626 95777
rect 66310 95712 66316 95776
rect 66380 95712 66396 95776
rect 66460 95712 66476 95776
rect 66540 95712 66556 95776
rect 66620 95712 66626 95776
rect 66310 95711 66626 95712
rect 97030 95776 97346 95777
rect 97030 95712 97036 95776
rect 97100 95712 97116 95776
rect 97180 95712 97196 95776
rect 97260 95712 97276 95776
rect 97340 95712 97346 95776
rect 97030 95711 97346 95712
rect 4210 95232 4526 95233
rect 4210 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4526 95232
rect 4210 95167 4526 95168
rect 34930 95232 35246 95233
rect 34930 95168 34936 95232
rect 35000 95168 35016 95232
rect 35080 95168 35096 95232
rect 35160 95168 35176 95232
rect 35240 95168 35246 95232
rect 34930 95167 35246 95168
rect 65650 95232 65966 95233
rect 65650 95168 65656 95232
rect 65720 95168 65736 95232
rect 65800 95168 65816 95232
rect 65880 95168 65896 95232
rect 65960 95168 65966 95232
rect 65650 95167 65966 95168
rect 96370 95232 96686 95233
rect 96370 95168 96376 95232
rect 96440 95168 96456 95232
rect 96520 95168 96536 95232
rect 96600 95168 96616 95232
rect 96680 95168 96686 95232
rect 96370 95167 96686 95168
rect 4870 94688 5186 94689
rect 4870 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5186 94688
rect 4870 94623 5186 94624
rect 35590 94688 35906 94689
rect 35590 94624 35596 94688
rect 35660 94624 35676 94688
rect 35740 94624 35756 94688
rect 35820 94624 35836 94688
rect 35900 94624 35906 94688
rect 35590 94623 35906 94624
rect 66310 94688 66626 94689
rect 66310 94624 66316 94688
rect 66380 94624 66396 94688
rect 66460 94624 66476 94688
rect 66540 94624 66556 94688
rect 66620 94624 66626 94688
rect 66310 94623 66626 94624
rect 97030 94688 97346 94689
rect 97030 94624 97036 94688
rect 97100 94624 97116 94688
rect 97180 94624 97196 94688
rect 97260 94624 97276 94688
rect 97340 94624 97346 94688
rect 97030 94623 97346 94624
rect 4210 94144 4526 94145
rect 4210 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4526 94144
rect 4210 94079 4526 94080
rect 34930 94144 35246 94145
rect 34930 94080 34936 94144
rect 35000 94080 35016 94144
rect 35080 94080 35096 94144
rect 35160 94080 35176 94144
rect 35240 94080 35246 94144
rect 34930 94079 35246 94080
rect 65650 94144 65966 94145
rect 65650 94080 65656 94144
rect 65720 94080 65736 94144
rect 65800 94080 65816 94144
rect 65880 94080 65896 94144
rect 65960 94080 65966 94144
rect 65650 94079 65966 94080
rect 96370 94144 96686 94145
rect 96370 94080 96376 94144
rect 96440 94080 96456 94144
rect 96520 94080 96536 94144
rect 96600 94080 96616 94144
rect 96680 94080 96686 94144
rect 96370 94079 96686 94080
rect 49366 93876 49372 93940
rect 49436 93938 49442 93940
rect 55581 93938 55647 93941
rect 49436 93936 55647 93938
rect 49436 93880 55586 93936
rect 55642 93880 55647 93936
rect 49436 93878 55647 93880
rect 49436 93876 49442 93878
rect 55581 93875 55647 93878
rect 65885 93802 65951 93805
rect 67265 93802 67331 93805
rect 65885 93800 67331 93802
rect 65885 93744 65890 93800
rect 65946 93744 67270 93800
rect 67326 93744 67331 93800
rect 65885 93742 67331 93744
rect 65885 93739 65951 93742
rect 67265 93739 67331 93742
rect 4870 93600 5186 93601
rect 4870 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5186 93600
rect 4870 93535 5186 93536
rect 35590 93600 35906 93601
rect 35590 93536 35596 93600
rect 35660 93536 35676 93600
rect 35740 93536 35756 93600
rect 35820 93536 35836 93600
rect 35900 93536 35906 93600
rect 35590 93535 35906 93536
rect 66310 93600 66626 93601
rect 66310 93536 66316 93600
rect 66380 93536 66396 93600
rect 66460 93536 66476 93600
rect 66540 93536 66556 93600
rect 66620 93536 66626 93600
rect 66310 93535 66626 93536
rect 97030 93600 97346 93601
rect 97030 93536 97036 93600
rect 97100 93536 97116 93600
rect 97180 93536 97196 93600
rect 97260 93536 97276 93600
rect 97340 93536 97346 93600
rect 97030 93535 97346 93536
rect 42006 93196 42012 93260
rect 42076 93258 42082 93260
rect 49325 93258 49391 93261
rect 42076 93256 49391 93258
rect 42076 93200 49330 93256
rect 49386 93200 49391 93256
rect 42076 93198 49391 93200
rect 42076 93196 42082 93198
rect 49325 93195 49391 93198
rect 64873 93258 64939 93261
rect 69197 93258 69263 93261
rect 64873 93256 69263 93258
rect 64873 93200 64878 93256
rect 64934 93200 69202 93256
rect 69258 93200 69263 93256
rect 64873 93198 69263 93200
rect 64873 93195 64939 93198
rect 69197 93195 69263 93198
rect 4210 93056 4526 93057
rect 4210 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4526 93056
rect 4210 92991 4526 92992
rect 34930 93056 35246 93057
rect 34930 92992 34936 93056
rect 35000 92992 35016 93056
rect 35080 92992 35096 93056
rect 35160 92992 35176 93056
rect 35240 92992 35246 93056
rect 34930 92991 35246 92992
rect 65650 93056 65966 93057
rect 65650 92992 65656 93056
rect 65720 92992 65736 93056
rect 65800 92992 65816 93056
rect 65880 92992 65896 93056
rect 65960 92992 65966 93056
rect 65650 92991 65966 92992
rect 96370 93056 96686 93057
rect 96370 92992 96376 93056
rect 96440 92992 96456 93056
rect 96520 92992 96536 93056
rect 96600 92992 96616 93056
rect 96680 92992 96686 93056
rect 96370 92991 96686 92992
rect 56910 92924 56916 92988
rect 56980 92986 56986 92988
rect 63493 92986 63559 92989
rect 56980 92984 63559 92986
rect 56980 92928 63498 92984
rect 63554 92928 63559 92984
rect 56980 92926 63559 92928
rect 56980 92924 56986 92926
rect 63493 92923 63559 92926
rect 44582 92788 44588 92852
rect 44652 92850 44658 92852
rect 50613 92850 50679 92853
rect 44652 92848 50679 92850
rect 44652 92792 50618 92848
rect 50674 92792 50679 92848
rect 44652 92790 50679 92792
rect 44652 92788 44658 92790
rect 50613 92787 50679 92790
rect 51942 92788 51948 92852
rect 52012 92850 52018 92852
rect 57973 92850 58039 92853
rect 58433 92850 58499 92853
rect 52012 92848 58499 92850
rect 52012 92792 57978 92848
rect 58034 92792 58438 92848
rect 58494 92792 58499 92848
rect 52012 92790 58499 92792
rect 52012 92788 52018 92790
rect 57973 92787 58039 92790
rect 58433 92787 58499 92790
rect 39614 92652 39620 92716
rect 39684 92714 39690 92716
rect 47117 92714 47183 92717
rect 52545 92714 52611 92717
rect 39684 92712 47183 92714
rect 39684 92656 47122 92712
rect 47178 92656 47183 92712
rect 39684 92654 47183 92656
rect 39684 92652 39690 92654
rect 47117 92651 47183 92654
rect 48086 92712 52611 92714
rect 48086 92656 52550 92712
rect 52606 92656 52611 92712
rect 48086 92654 52611 92656
rect 38142 92516 38148 92580
rect 38212 92578 38218 92580
rect 44173 92578 44239 92581
rect 38212 92576 44239 92578
rect 38212 92520 44178 92576
rect 44234 92520 44239 92576
rect 38212 92518 44239 92520
rect 38212 92516 38218 92518
rect 44173 92515 44239 92518
rect 45870 92516 45876 92580
rect 45940 92578 45946 92580
rect 48086 92578 48146 92654
rect 52545 92651 52611 92654
rect 59813 92714 59879 92717
rect 61878 92714 61884 92716
rect 59813 92712 61884 92714
rect 59813 92656 59818 92712
rect 59874 92656 61884 92712
rect 59813 92654 61884 92656
rect 59813 92651 59879 92654
rect 61878 92652 61884 92654
rect 61948 92652 61954 92716
rect 45940 92518 48146 92578
rect 45940 92516 45946 92518
rect 48262 92516 48268 92580
rect 48332 92578 48338 92580
rect 54017 92578 54083 92581
rect 48332 92576 54083 92578
rect 48332 92520 54022 92576
rect 54078 92520 54083 92576
rect 48332 92518 54083 92520
rect 48332 92516 48338 92518
rect 54017 92515 54083 92518
rect 56593 92578 56659 92581
rect 63493 92578 63559 92581
rect 56593 92576 63559 92578
rect 56593 92520 56598 92576
rect 56654 92520 63498 92576
rect 63554 92520 63559 92576
rect 56593 92518 63559 92520
rect 56593 92515 56659 92518
rect 63493 92515 63559 92518
rect 63769 92578 63835 92581
rect 69197 92580 69263 92581
rect 64270 92578 64276 92580
rect 63769 92576 64276 92578
rect 63769 92520 63774 92576
rect 63830 92520 64276 92576
rect 63769 92518 64276 92520
rect 63769 92515 63835 92518
rect 64270 92516 64276 92518
rect 64340 92516 64346 92580
rect 69197 92576 69244 92580
rect 69308 92578 69314 92580
rect 70485 92578 70551 92581
rect 70710 92578 70716 92580
rect 69197 92520 69202 92576
rect 69197 92516 69244 92520
rect 69308 92518 69354 92578
rect 70485 92576 70716 92578
rect 70485 92520 70490 92576
rect 70546 92520 70716 92576
rect 70485 92518 70716 92520
rect 69308 92516 69314 92518
rect 69197 92515 69263 92516
rect 70485 92515 70551 92518
rect 70710 92516 70716 92518
rect 70780 92516 70786 92580
rect 4870 92512 5186 92513
rect 4870 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5186 92512
rect 4870 92447 5186 92448
rect 35590 92512 35906 92513
rect 35590 92448 35596 92512
rect 35660 92448 35676 92512
rect 35740 92448 35756 92512
rect 35820 92448 35836 92512
rect 35900 92448 35906 92512
rect 35590 92447 35906 92448
rect 66310 92512 66626 92513
rect 66310 92448 66316 92512
rect 66380 92448 66396 92512
rect 66460 92448 66476 92512
rect 66540 92448 66556 92512
rect 66620 92448 66626 92512
rect 66310 92447 66626 92448
rect 97030 92512 97346 92513
rect 97030 92448 97036 92512
rect 97100 92448 97116 92512
rect 97180 92448 97196 92512
rect 97260 92448 97276 92512
rect 97340 92448 97346 92512
rect 97030 92447 97346 92448
rect 113646 92512 113962 92513
rect 113646 92448 113652 92512
rect 113716 92448 113732 92512
rect 113796 92448 113812 92512
rect 113876 92448 113892 92512
rect 113956 92448 113962 92512
rect 113646 92447 113962 92448
rect 43294 92108 43300 92172
rect 43364 92170 43370 92172
rect 50245 92170 50311 92173
rect 43364 92168 50311 92170
rect 43364 92112 50250 92168
rect 50306 92112 50311 92168
rect 43364 92110 50311 92112
rect 43364 92108 43370 92110
rect 50245 92107 50311 92110
rect 50654 92108 50660 92172
rect 50724 92170 50730 92172
rect 52913 92170 52979 92173
rect 50724 92168 52979 92170
rect 50724 92112 52918 92168
rect 52974 92112 52979 92168
rect 50724 92110 52979 92112
rect 50724 92108 50730 92110
rect 52913 92107 52979 92110
rect 53230 92108 53236 92172
rect 53300 92170 53306 92172
rect 58709 92170 58775 92173
rect 53300 92168 58775 92170
rect 53300 92112 58714 92168
rect 58770 92112 58775 92168
rect 53300 92110 58775 92112
rect 53300 92108 53306 92110
rect 58709 92107 58775 92110
rect 46790 91972 46796 92036
rect 46860 92034 46866 92036
rect 53189 92034 53255 92037
rect 46860 92032 53255 92034
rect 46860 91976 53194 92032
rect 53250 91976 53255 92032
rect 46860 91974 53255 91976
rect 46860 91972 46866 91974
rect 53189 91971 53255 91974
rect 4210 91968 4526 91969
rect 4210 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4526 91968
rect 4210 91903 4526 91904
rect 34930 91968 35246 91969
rect 34930 91904 34936 91968
rect 35000 91904 35016 91968
rect 35080 91904 35096 91968
rect 35160 91904 35176 91968
rect 35240 91904 35246 91968
rect 34930 91903 35246 91904
rect 65650 91968 65966 91969
rect 65650 91904 65656 91968
rect 65720 91904 65736 91968
rect 65800 91904 65816 91968
rect 65880 91904 65896 91968
rect 65960 91904 65966 91968
rect 65650 91903 65966 91904
rect 96370 91968 96686 91969
rect 96370 91904 96376 91968
rect 96440 91904 96456 91968
rect 96520 91904 96536 91968
rect 96600 91904 96616 91968
rect 96680 91904 96686 91968
rect 96370 91903 96686 91904
rect 112910 91968 113226 91969
rect 112910 91904 112916 91968
rect 112980 91904 112996 91968
rect 113060 91904 113076 91968
rect 113140 91904 113156 91968
rect 113220 91904 113226 91968
rect 112910 91903 113226 91904
rect 4870 91424 5186 91425
rect 4870 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5186 91424
rect 4870 91359 5186 91360
rect 113646 91424 113962 91425
rect 113646 91360 113652 91424
rect 113716 91360 113732 91424
rect 113796 91360 113812 91424
rect 113876 91360 113892 91424
rect 113956 91360 113962 91424
rect 113646 91359 113962 91360
rect 100017 91220 100083 91221
rect 99966 91218 99972 91220
rect 99926 91158 99972 91218
rect 100036 91216 100083 91220
rect 100078 91160 100083 91216
rect 99966 91156 99972 91158
rect 100036 91156 100083 91160
rect 100017 91155 100083 91156
rect 62849 91082 62915 91085
rect 73245 91084 73311 91085
rect 74165 91084 74231 91085
rect 62982 91082 62988 91084
rect 62849 91080 62988 91082
rect 62849 91024 62854 91080
rect 62910 91024 62988 91080
rect 62849 91022 62988 91024
rect 62849 91019 62915 91022
rect 62982 91020 62988 91022
rect 63052 91020 63058 91084
rect 73245 91080 73292 91084
rect 73356 91082 73362 91084
rect 73245 91024 73250 91080
rect 73245 91020 73292 91024
rect 73356 91022 73402 91082
rect 74165 91080 74212 91084
rect 74276 91082 74282 91084
rect 74165 91024 74170 91080
rect 73356 91020 73362 91022
rect 74165 91020 74212 91024
rect 74276 91022 74322 91082
rect 74276 91020 74282 91022
rect 73245 91019 73311 91020
rect 74165 91019 74231 91020
rect 4210 90880 4526 90881
rect 4210 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4526 90880
rect 4210 90815 4526 90816
rect 112910 90880 113226 90881
rect 112910 90816 112916 90880
rect 112980 90816 112996 90880
rect 113060 90816 113076 90880
rect 113140 90816 113156 90880
rect 113220 90816 113226 90880
rect 112910 90815 113226 90816
rect 4870 90336 5186 90337
rect 4870 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5186 90336
rect 4870 90271 5186 90272
rect 113646 90336 113962 90337
rect 113646 90272 113652 90336
rect 113716 90272 113732 90336
rect 113796 90272 113812 90336
rect 113876 90272 113892 90336
rect 113956 90272 113962 90336
rect 113646 90271 113962 90272
rect 58157 89996 58223 89997
rect 58144 89994 58150 89996
rect 58066 89934 58150 89994
rect 58214 89992 58223 89996
rect 58218 89936 58223 89992
rect 58144 89932 58150 89934
rect 58214 89932 58223 89936
rect 58157 89931 58223 89932
rect 59445 89996 59511 89997
rect 59445 89992 59510 89996
rect 59445 89936 59450 89992
rect 59506 89936 59510 89992
rect 59445 89932 59510 89936
rect 59574 89994 59580 89996
rect 59574 89934 59602 89994
rect 59574 89932 59580 89934
rect 59445 89931 59511 89932
rect 55560 89796 55566 89860
rect 55630 89858 55636 89860
rect 59261 89858 59327 89861
rect 55630 89856 59327 89858
rect 55630 89800 59266 89856
rect 59322 89800 59327 89856
rect 55630 89798 59327 89800
rect 55630 89796 55636 89798
rect 59261 89795 59327 89798
rect 4210 89792 4526 89793
rect 4210 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4526 89792
rect 4210 89727 4526 89728
rect 112910 89792 113226 89793
rect 112910 89728 112916 89792
rect 112980 89728 112996 89792
rect 113060 89728 113076 89792
rect 113140 89728 113156 89792
rect 113220 89728 113226 89792
rect 112910 89727 113226 89728
rect 40600 89660 40606 89724
rect 40670 89722 40676 89724
rect 46841 89722 46907 89725
rect 40670 89720 46907 89722
rect 40670 89664 46846 89720
rect 46902 89664 46907 89720
rect 40670 89662 46907 89664
rect 40670 89660 40676 89662
rect 46841 89659 46907 89662
rect 54336 89660 54342 89724
rect 54406 89722 54412 89724
rect 59353 89722 59419 89725
rect 60592 89722 60598 89724
rect 54406 89662 55230 89722
rect 54406 89660 54412 89662
rect 55170 89586 55230 89662
rect 59353 89720 60598 89722
rect 59353 89664 59358 89720
rect 59414 89664 60598 89720
rect 59353 89662 60598 89664
rect 59353 89659 59419 89662
rect 60592 89660 60598 89662
rect 60662 89660 60668 89724
rect 65241 89722 65307 89725
rect 66805 89724 66871 89725
rect 65624 89722 65630 89724
rect 65241 89720 65630 89722
rect 65241 89664 65246 89720
rect 65302 89664 65630 89720
rect 65241 89662 65630 89664
rect 65241 89659 65307 89662
rect 65624 89660 65630 89662
rect 65694 89660 65700 89724
rect 66805 89720 66854 89724
rect 66918 89722 66924 89724
rect 67541 89722 67607 89725
rect 71865 89724 71931 89725
rect 68208 89722 68214 89724
rect 66805 89664 66810 89720
rect 66805 89660 66854 89664
rect 66918 89662 66962 89722
rect 67541 89720 68214 89722
rect 67541 89664 67546 89720
rect 67602 89664 68214 89720
rect 67541 89662 68214 89664
rect 66918 89660 66924 89662
rect 66805 89659 66871 89660
rect 67541 89659 67607 89662
rect 68208 89660 68214 89662
rect 68278 89660 68284 89724
rect 71865 89720 71886 89724
rect 71950 89722 71956 89724
rect 73705 89722 73771 89725
rect 75552 89722 75558 89724
rect 71865 89664 71870 89720
rect 71865 89660 71886 89664
rect 71950 89662 72022 89722
rect 73705 89720 75558 89722
rect 73705 89664 73710 89720
rect 73766 89664 75558 89720
rect 73705 89662 75558 89664
rect 71950 89660 71956 89662
rect 71865 89659 71931 89660
rect 73705 89659 73771 89662
rect 75552 89660 75558 89662
rect 75622 89660 75628 89724
rect 75913 89722 75979 89725
rect 89437 89724 89503 89725
rect 76912 89722 76918 89724
rect 75913 89720 76918 89722
rect 75913 89664 75918 89720
rect 75974 89664 76918 89720
rect 75913 89662 76918 89664
rect 75913 89659 75979 89662
rect 76912 89660 76918 89662
rect 76982 89660 76988 89724
rect 89424 89722 89430 89724
rect 89346 89662 89430 89722
rect 89494 89722 89503 89724
rect 89494 89720 93870 89722
rect 89498 89664 93870 89720
rect 89424 89660 89430 89662
rect 89494 89662 93870 89664
rect 89494 89660 89503 89662
rect 89437 89659 89503 89660
rect 60549 89586 60615 89589
rect 55170 89584 60615 89586
rect 55170 89528 60554 89584
rect 60610 89528 60615 89584
rect 55170 89526 60615 89528
rect 93810 89586 93870 89662
rect 106917 89586 106983 89589
rect 93810 89584 106983 89586
rect 93810 89528 106922 89584
rect 106978 89528 106983 89584
rect 93810 89526 106983 89528
rect 60549 89523 60615 89526
rect 106917 89523 106983 89526
rect 4870 89248 5186 89249
rect 4870 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5186 89248
rect 4870 89183 5186 89184
rect 113646 89248 113962 89249
rect 113646 89184 113652 89248
rect 113716 89184 113732 89248
rect 113796 89184 113812 89248
rect 113876 89184 113892 89248
rect 113956 89184 113962 89248
rect 113646 89183 113962 89184
rect 4210 88704 4526 88705
rect 4210 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4526 88704
rect 4210 88639 4526 88640
rect 112910 88704 113226 88705
rect 112910 88640 112916 88704
rect 112980 88640 112996 88704
rect 113060 88640 113076 88704
rect 113140 88640 113156 88704
rect 113220 88640 113226 88704
rect 112910 88639 113226 88640
rect 4870 88160 5186 88161
rect 4870 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5186 88160
rect 4870 88095 5186 88096
rect 113646 88160 113962 88161
rect 113646 88096 113652 88160
rect 113716 88096 113732 88160
rect 113796 88096 113812 88160
rect 113876 88096 113892 88160
rect 113956 88096 113962 88160
rect 113646 88095 113962 88096
rect 4210 87616 4526 87617
rect 4210 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4526 87616
rect 4210 87551 4526 87552
rect 112910 87616 113226 87617
rect 112910 87552 112916 87616
rect 112980 87552 112996 87616
rect 113060 87552 113076 87616
rect 113140 87552 113156 87616
rect 113220 87552 113226 87616
rect 112910 87551 113226 87552
rect 4870 87072 5186 87073
rect 4870 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5186 87072
rect 4870 87007 5186 87008
rect 113646 87072 113962 87073
rect 113646 87008 113652 87072
rect 113716 87008 113732 87072
rect 113796 87008 113812 87072
rect 113876 87008 113892 87072
rect 113956 87008 113962 87072
rect 113646 87007 113962 87008
rect 4210 86528 4526 86529
rect 4210 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4526 86528
rect 112910 86528 113226 86529
rect 106181 86500 106247 86503
rect 4210 86463 4526 86464
rect 105892 86498 106247 86500
rect 105892 86442 106186 86498
rect 106242 86442 106247 86498
rect 112910 86464 112916 86528
rect 112980 86464 112996 86528
rect 113060 86464 113076 86528
rect 113140 86464 113156 86528
rect 113220 86464 113226 86528
rect 112910 86463 113226 86464
rect 105892 86440 106247 86442
rect 106181 86437 106247 86440
rect 4870 85984 5186 85985
rect 4870 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5186 85984
rect 4870 85919 5186 85920
rect 113646 85984 113962 85985
rect 113646 85920 113652 85984
rect 113716 85920 113732 85984
rect 113796 85920 113812 85984
rect 113876 85920 113892 85984
rect 113956 85920 113962 85984
rect 113646 85919 113962 85920
rect 4210 85440 4526 85441
rect 4210 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4526 85440
rect 4210 85375 4526 85376
rect 112910 85440 113226 85441
rect 112910 85376 112916 85440
rect 112980 85376 112996 85440
rect 113060 85376 113076 85440
rect 113140 85376 113156 85440
rect 113220 85376 113226 85440
rect 112910 85375 113226 85376
rect 4870 84896 5186 84897
rect 4870 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5186 84896
rect 4870 84831 5186 84832
rect 113646 84896 113962 84897
rect 113646 84832 113652 84896
rect 113716 84832 113732 84896
rect 113796 84832 113812 84896
rect 113876 84832 113892 84896
rect 113956 84832 113962 84896
rect 113646 84831 113962 84832
rect 4210 84352 4526 84353
rect 4210 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4526 84352
rect 4210 84287 4526 84288
rect 112910 84352 113226 84353
rect 112910 84288 112916 84352
rect 112980 84288 112996 84352
rect 113060 84288 113076 84352
rect 113140 84288 113156 84352
rect 113220 84288 113226 84352
rect 112910 84287 113226 84288
rect 4870 83808 5186 83809
rect 4870 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5186 83808
rect 4870 83743 5186 83744
rect 113646 83808 113962 83809
rect 113646 83744 113652 83808
rect 113716 83744 113732 83808
rect 113796 83744 113812 83808
rect 113876 83744 113892 83808
rect 113956 83744 113962 83808
rect 113646 83743 113962 83744
rect 4210 83264 4526 83265
rect 4210 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4526 83264
rect 4210 83199 4526 83200
rect 112910 83264 113226 83265
rect 112910 83200 112916 83264
rect 112980 83200 112996 83264
rect 113060 83200 113076 83264
rect 113140 83200 113156 83264
rect 113220 83200 113226 83264
rect 112910 83199 113226 83200
rect 4870 82720 5186 82721
rect 4870 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5186 82720
rect 4870 82655 5186 82656
rect 113646 82720 113962 82721
rect 113646 82656 113652 82720
rect 113716 82656 113732 82720
rect 113796 82656 113812 82720
rect 113876 82656 113892 82720
rect 113956 82656 113962 82720
rect 113646 82655 113962 82656
rect 4210 82176 4526 82177
rect 4210 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4526 82176
rect 4210 82111 4526 82112
rect 112910 82176 113226 82177
rect 112910 82112 112916 82176
rect 112980 82112 112996 82176
rect 113060 82112 113076 82176
rect 113140 82112 113156 82176
rect 113220 82112 113226 82176
rect 112910 82111 113226 82112
rect 4870 81632 5186 81633
rect 4870 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5186 81632
rect 4870 81567 5186 81568
rect 113646 81632 113962 81633
rect 113646 81568 113652 81632
rect 113716 81568 113732 81632
rect 113796 81568 113812 81632
rect 113876 81568 113892 81632
rect 113956 81568 113962 81632
rect 113646 81567 113962 81568
rect 4210 81088 4526 81089
rect 4210 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4526 81088
rect 4210 81023 4526 81024
rect 112910 81088 113226 81089
rect 112910 81024 112916 81088
rect 112980 81024 112996 81088
rect 113060 81024 113076 81088
rect 113140 81024 113156 81088
rect 113220 81024 113226 81088
rect 112910 81023 113226 81024
rect 4870 80544 5186 80545
rect 4870 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5186 80544
rect 4870 80479 5186 80480
rect 113646 80544 113962 80545
rect 113646 80480 113652 80544
rect 113716 80480 113732 80544
rect 113796 80480 113812 80544
rect 113876 80480 113892 80544
rect 113956 80480 113962 80544
rect 113646 80479 113962 80480
rect 4210 80000 4526 80001
rect 4210 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4526 80000
rect 4210 79935 4526 79936
rect 112910 80000 113226 80001
rect 112910 79936 112916 80000
rect 112980 79936 112996 80000
rect 113060 79936 113076 80000
rect 113140 79936 113156 80000
rect 113220 79936 113226 80000
rect 112910 79935 113226 79936
rect 4870 79456 5186 79457
rect 4870 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5186 79456
rect 4870 79391 5186 79392
rect 113646 79456 113962 79457
rect 113646 79392 113652 79456
rect 113716 79392 113732 79456
rect 113796 79392 113812 79456
rect 113876 79392 113892 79456
rect 113956 79392 113962 79456
rect 113646 79391 113962 79392
rect 4210 78912 4526 78913
rect 4210 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4526 78912
rect 4210 78847 4526 78848
rect 112910 78912 113226 78913
rect 112910 78848 112916 78912
rect 112980 78848 112996 78912
rect 113060 78848 113076 78912
rect 113140 78848 113156 78912
rect 113220 78848 113226 78912
rect 112910 78847 113226 78848
rect 4870 78368 5186 78369
rect 4870 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5186 78368
rect 4870 78303 5186 78304
rect 113646 78368 113962 78369
rect 113646 78304 113652 78368
rect 113716 78304 113732 78368
rect 113796 78304 113812 78368
rect 113876 78304 113892 78368
rect 113956 78304 113962 78368
rect 113646 78303 113962 78304
rect 4210 77824 4526 77825
rect 4210 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4526 77824
rect 4210 77759 4526 77760
rect 112910 77824 113226 77825
rect 112910 77760 112916 77824
rect 112980 77760 112996 77824
rect 113060 77760 113076 77824
rect 113140 77760 113156 77824
rect 113220 77760 113226 77824
rect 112910 77759 113226 77760
rect 4870 77280 5186 77281
rect 4870 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5186 77280
rect 4870 77215 5186 77216
rect 113646 77280 113962 77281
rect 113646 77216 113652 77280
rect 113716 77216 113732 77280
rect 113796 77216 113812 77280
rect 113876 77216 113892 77280
rect 113956 77216 113962 77280
rect 113646 77215 113962 77216
rect 4210 76736 4526 76737
rect 4210 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4526 76736
rect 4210 76671 4526 76672
rect 112910 76736 113226 76737
rect 112910 76672 112916 76736
rect 112980 76672 112996 76736
rect 113060 76672 113076 76736
rect 113140 76672 113156 76736
rect 113220 76672 113226 76736
rect 112910 76671 113226 76672
rect 4870 76192 5186 76193
rect 4870 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5186 76192
rect 4870 76127 5186 76128
rect 113646 76192 113962 76193
rect 113646 76128 113652 76192
rect 113716 76128 113732 76192
rect 113796 76128 113812 76192
rect 113876 76128 113892 76192
rect 113956 76128 113962 76192
rect 113646 76127 113962 76128
rect 4210 75648 4526 75649
rect 4210 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4526 75648
rect 4210 75583 4526 75584
rect 112910 75648 113226 75649
rect 112910 75584 112916 75648
rect 112980 75584 112996 75648
rect 113060 75584 113076 75648
rect 113140 75584 113156 75648
rect 113220 75584 113226 75648
rect 112910 75583 113226 75584
rect 4870 75104 5186 75105
rect 4870 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5186 75104
rect 4870 75039 5186 75040
rect 113646 75104 113962 75105
rect 113646 75040 113652 75104
rect 113716 75040 113732 75104
rect 113796 75040 113812 75104
rect 113876 75040 113892 75104
rect 113956 75040 113962 75104
rect 113646 75039 113962 75040
rect 4210 74560 4526 74561
rect 4210 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4526 74560
rect 4210 74495 4526 74496
rect 112910 74560 113226 74561
rect 112910 74496 112916 74560
rect 112980 74496 112996 74560
rect 113060 74496 113076 74560
rect 113140 74496 113156 74560
rect 113220 74496 113226 74560
rect 112910 74495 113226 74496
rect 4870 74016 5186 74017
rect 4870 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5186 74016
rect 4870 73951 5186 73952
rect 113646 74016 113962 74017
rect 113646 73952 113652 74016
rect 113716 73952 113732 74016
rect 113796 73952 113812 74016
rect 113876 73952 113892 74016
rect 113956 73952 113962 74016
rect 113646 73951 113962 73952
rect 4210 73472 4526 73473
rect 4210 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4526 73472
rect 4210 73407 4526 73408
rect 112910 73472 113226 73473
rect 112910 73408 112916 73472
rect 112980 73408 112996 73472
rect 113060 73408 113076 73472
rect 113140 73408 113156 73472
rect 113220 73408 113226 73472
rect 112910 73407 113226 73408
rect 4870 72928 5186 72929
rect 4870 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5186 72928
rect 4870 72863 5186 72864
rect 113646 72928 113962 72929
rect 113646 72864 113652 72928
rect 113716 72864 113732 72928
rect 113796 72864 113812 72928
rect 113876 72864 113892 72928
rect 113956 72864 113962 72928
rect 113646 72863 113962 72864
rect 4210 72384 4526 72385
rect 4210 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4526 72384
rect 4210 72319 4526 72320
rect 112910 72384 113226 72385
rect 112910 72320 112916 72384
rect 112980 72320 112996 72384
rect 113060 72320 113076 72384
rect 113140 72320 113156 72384
rect 113220 72320 113226 72384
rect 112910 72319 113226 72320
rect 4870 71840 5186 71841
rect 4870 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5186 71840
rect 4870 71775 5186 71776
rect 113646 71840 113962 71841
rect 113646 71776 113652 71840
rect 113716 71776 113732 71840
rect 113796 71776 113812 71840
rect 113876 71776 113892 71840
rect 113956 71776 113962 71840
rect 113646 71775 113962 71776
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 112910 71296 113226 71297
rect 112910 71232 112916 71296
rect 112980 71232 112996 71296
rect 113060 71232 113076 71296
rect 113140 71232 113156 71296
rect 113220 71232 113226 71296
rect 112910 71231 113226 71232
rect 4870 70752 5186 70753
rect 4870 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5186 70752
rect 4870 70687 5186 70688
rect 113646 70752 113962 70753
rect 113646 70688 113652 70752
rect 113716 70688 113732 70752
rect 113796 70688 113812 70752
rect 113876 70688 113892 70752
rect 113956 70688 113962 70752
rect 113646 70687 113962 70688
rect 4210 70208 4526 70209
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 112910 70208 113226 70209
rect 112910 70144 112916 70208
rect 112980 70144 112996 70208
rect 113060 70144 113076 70208
rect 113140 70144 113156 70208
rect 113220 70144 113226 70208
rect 112910 70143 113226 70144
rect 4870 69664 5186 69665
rect 4870 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5186 69664
rect 4870 69599 5186 69600
rect 113646 69664 113962 69665
rect 113646 69600 113652 69664
rect 113716 69600 113732 69664
rect 113796 69600 113812 69664
rect 113876 69600 113892 69664
rect 113956 69600 113962 69664
rect 113646 69599 113962 69600
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 112910 69120 113226 69121
rect 112910 69056 112916 69120
rect 112980 69056 112996 69120
rect 113060 69056 113076 69120
rect 113140 69056 113156 69120
rect 113220 69056 113226 69120
rect 112910 69055 113226 69056
rect 4870 68576 5186 68577
rect 4870 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5186 68576
rect 4870 68511 5186 68512
rect 113646 68576 113962 68577
rect 113646 68512 113652 68576
rect 113716 68512 113732 68576
rect 113796 68512 113812 68576
rect 113876 68512 113892 68576
rect 113956 68512 113962 68576
rect 113646 68511 113962 68512
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 112910 68032 113226 68033
rect 112910 67968 112916 68032
rect 112980 67968 112996 68032
rect 113060 67968 113076 68032
rect 113140 67968 113156 68032
rect 113220 67968 113226 68032
rect 112910 67967 113226 67968
rect 4870 67488 5186 67489
rect 4870 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5186 67488
rect 4870 67423 5186 67424
rect 113646 67488 113962 67489
rect 113646 67424 113652 67488
rect 113716 67424 113732 67488
rect 113796 67424 113812 67488
rect 113876 67424 113892 67488
rect 113956 67424 113962 67488
rect 113646 67423 113962 67424
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 112910 66944 113226 66945
rect 112910 66880 112916 66944
rect 112980 66880 112996 66944
rect 113060 66880 113076 66944
rect 113140 66880 113156 66944
rect 113220 66880 113226 66944
rect 112910 66879 113226 66880
rect 4870 66400 5186 66401
rect 4870 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5186 66400
rect 4870 66335 5186 66336
rect 113646 66400 113962 66401
rect 113646 66336 113652 66400
rect 113716 66336 113732 66400
rect 113796 66336 113812 66400
rect 113876 66336 113892 66400
rect 113956 66336 113962 66400
rect 113646 66335 113962 66336
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 112910 65856 113226 65857
rect 112910 65792 112916 65856
rect 112980 65792 112996 65856
rect 113060 65792 113076 65856
rect 113140 65792 113156 65856
rect 113220 65792 113226 65856
rect 112910 65791 113226 65792
rect 4870 65312 5186 65313
rect 4870 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5186 65312
rect 4870 65247 5186 65248
rect 113646 65312 113962 65313
rect 113646 65248 113652 65312
rect 113716 65248 113732 65312
rect 113796 65248 113812 65312
rect 113876 65248 113892 65312
rect 113956 65248 113962 65312
rect 113646 65247 113962 65248
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 112910 64768 113226 64769
rect 112910 64704 112916 64768
rect 112980 64704 112996 64768
rect 113060 64704 113076 64768
rect 113140 64704 113156 64768
rect 113220 64704 113226 64768
rect 112910 64703 113226 64704
rect 4870 64224 5186 64225
rect 4870 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5186 64224
rect 4870 64159 5186 64160
rect 113646 64224 113962 64225
rect 113646 64160 113652 64224
rect 113716 64160 113732 64224
rect 113796 64160 113812 64224
rect 113876 64160 113892 64224
rect 113956 64160 113962 64224
rect 113646 64159 113962 64160
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 112910 63680 113226 63681
rect 112910 63616 112916 63680
rect 112980 63616 112996 63680
rect 113060 63616 113076 63680
rect 113140 63616 113156 63680
rect 113220 63616 113226 63680
rect 112910 63615 113226 63616
rect 4870 63136 5186 63137
rect 4870 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5186 63136
rect 4870 63071 5186 63072
rect 113646 63136 113962 63137
rect 113646 63072 113652 63136
rect 113716 63072 113732 63136
rect 113796 63072 113812 63136
rect 113876 63072 113892 63136
rect 113956 63072 113962 63136
rect 113646 63071 113962 63072
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 112910 62592 113226 62593
rect 112910 62528 112916 62592
rect 112980 62528 112996 62592
rect 113060 62528 113076 62592
rect 113140 62528 113156 62592
rect 113220 62528 113226 62592
rect 112910 62527 113226 62528
rect 4870 62048 5186 62049
rect 4870 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5186 62048
rect 4870 61983 5186 61984
rect 113646 62048 113962 62049
rect 113646 61984 113652 62048
rect 113716 61984 113732 62048
rect 113796 61984 113812 62048
rect 113876 61984 113892 62048
rect 113956 61984 113962 62048
rect 113646 61983 113962 61984
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 112910 61504 113226 61505
rect 112910 61440 112916 61504
rect 112980 61440 112996 61504
rect 113060 61440 113076 61504
rect 113140 61440 113156 61504
rect 113220 61440 113226 61504
rect 112910 61439 113226 61440
rect 4870 60960 5186 60961
rect 4870 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5186 60960
rect 4870 60895 5186 60896
rect 113646 60960 113962 60961
rect 113646 60896 113652 60960
rect 113716 60896 113732 60960
rect 113796 60896 113812 60960
rect 113876 60896 113892 60960
rect 113956 60896 113962 60960
rect 113646 60895 113962 60896
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 112910 60416 113226 60417
rect 112910 60352 112916 60416
rect 112980 60352 112996 60416
rect 113060 60352 113076 60416
rect 113140 60352 113156 60416
rect 113220 60352 113226 60416
rect 112910 60351 113226 60352
rect 4870 59872 5186 59873
rect 4870 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5186 59872
rect 4870 59807 5186 59808
rect 113646 59872 113962 59873
rect 113646 59808 113652 59872
rect 113716 59808 113732 59872
rect 113796 59808 113812 59872
rect 113876 59808 113892 59872
rect 113956 59808 113962 59872
rect 113646 59807 113962 59808
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 112910 59328 113226 59329
rect 112910 59264 112916 59328
rect 112980 59264 112996 59328
rect 113060 59264 113076 59328
rect 113140 59264 113156 59328
rect 113220 59264 113226 59328
rect 112910 59263 113226 59264
rect 4870 58784 5186 58785
rect 4870 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5186 58784
rect 4870 58719 5186 58720
rect 113646 58784 113962 58785
rect 113646 58720 113652 58784
rect 113716 58720 113732 58784
rect 113796 58720 113812 58784
rect 113876 58720 113892 58784
rect 113956 58720 113962 58784
rect 113646 58719 113962 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 112910 58240 113226 58241
rect 112910 58176 112916 58240
rect 112980 58176 112996 58240
rect 113060 58176 113076 58240
rect 113140 58176 113156 58240
rect 113220 58176 113226 58240
rect 112910 58175 113226 58176
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 113646 57696 113962 57697
rect 113646 57632 113652 57696
rect 113716 57632 113732 57696
rect 113796 57632 113812 57696
rect 113876 57632 113892 57696
rect 113956 57632 113962 57696
rect 113646 57631 113962 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 112910 57152 113226 57153
rect 112910 57088 112916 57152
rect 112980 57088 112996 57152
rect 113060 57088 113076 57152
rect 113140 57088 113156 57152
rect 113220 57088 113226 57152
rect 112910 57087 113226 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 113646 56608 113962 56609
rect 113646 56544 113652 56608
rect 113716 56544 113732 56608
rect 113796 56544 113812 56608
rect 113876 56544 113892 56608
rect 113956 56544 113962 56608
rect 113646 56543 113962 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 112910 56064 113226 56065
rect 112910 56000 112916 56064
rect 112980 56000 112996 56064
rect 113060 56000 113076 56064
rect 113140 56000 113156 56064
rect 113220 56000 113226 56064
rect 112910 55999 113226 56000
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 113646 55520 113962 55521
rect 113646 55456 113652 55520
rect 113716 55456 113732 55520
rect 113796 55456 113812 55520
rect 113876 55456 113892 55520
rect 113956 55456 113962 55520
rect 113646 55455 113962 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 112910 54976 113226 54977
rect 112910 54912 112916 54976
rect 112980 54912 112996 54976
rect 113060 54912 113076 54976
rect 113140 54912 113156 54976
rect 113220 54912 113226 54976
rect 112910 54911 113226 54912
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 113646 54432 113962 54433
rect 113646 54368 113652 54432
rect 113716 54368 113732 54432
rect 113796 54368 113812 54432
rect 113876 54368 113892 54432
rect 113956 54368 113962 54432
rect 113646 54367 113962 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 112910 53888 113226 53889
rect 112910 53824 112916 53888
rect 112980 53824 112996 53888
rect 113060 53824 113076 53888
rect 113140 53824 113156 53888
rect 113220 53824 113226 53888
rect 112910 53823 113226 53824
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 113646 53344 113962 53345
rect 113646 53280 113652 53344
rect 113716 53280 113732 53344
rect 113796 53280 113812 53344
rect 113876 53280 113892 53344
rect 113956 53280 113962 53344
rect 113646 53279 113962 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 112910 52800 113226 52801
rect 112910 52736 112916 52800
rect 112980 52736 112996 52800
rect 113060 52736 113076 52800
rect 113140 52736 113156 52800
rect 113220 52736 113226 52800
rect 112910 52735 113226 52736
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 113646 52256 113962 52257
rect 113646 52192 113652 52256
rect 113716 52192 113732 52256
rect 113796 52192 113812 52256
rect 113876 52192 113892 52256
rect 113956 52192 113962 52256
rect 113646 52191 113962 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 112910 51712 113226 51713
rect 112910 51648 112916 51712
rect 112980 51648 112996 51712
rect 113060 51648 113076 51712
rect 113140 51648 113156 51712
rect 113220 51648 113226 51712
rect 112910 51647 113226 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 113646 51168 113962 51169
rect 113646 51104 113652 51168
rect 113716 51104 113732 51168
rect 113796 51104 113812 51168
rect 113876 51104 113892 51168
rect 113956 51104 113962 51168
rect 113646 51103 113962 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 112910 50624 113226 50625
rect 112910 50560 112916 50624
rect 112980 50560 112996 50624
rect 113060 50560 113076 50624
rect 113140 50560 113156 50624
rect 113220 50560 113226 50624
rect 112910 50559 113226 50560
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 113646 50080 113962 50081
rect 113646 50016 113652 50080
rect 113716 50016 113732 50080
rect 113796 50016 113812 50080
rect 113876 50016 113892 50080
rect 113956 50016 113962 50080
rect 113646 50015 113962 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 112910 49536 113226 49537
rect 112910 49472 112916 49536
rect 112980 49472 112996 49536
rect 113060 49472 113076 49536
rect 113140 49472 113156 49536
rect 113220 49472 113226 49536
rect 112910 49471 113226 49472
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 113646 48992 113962 48993
rect 113646 48928 113652 48992
rect 113716 48928 113732 48992
rect 113796 48928 113812 48992
rect 113876 48928 113892 48992
rect 113956 48928 113962 48992
rect 113646 48927 113962 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 112910 48448 113226 48449
rect 112910 48384 112916 48448
rect 112980 48384 112996 48448
rect 113060 48384 113076 48448
rect 113140 48384 113156 48448
rect 113220 48384 113226 48448
rect 112910 48383 113226 48384
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 113646 47904 113962 47905
rect 113646 47840 113652 47904
rect 113716 47840 113732 47904
rect 113796 47840 113812 47904
rect 113876 47840 113892 47904
rect 113956 47840 113962 47904
rect 113646 47839 113962 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 112910 47360 113226 47361
rect 112910 47296 112916 47360
rect 112980 47296 112996 47360
rect 113060 47296 113076 47360
rect 113140 47296 113156 47360
rect 113220 47296 113226 47360
rect 112910 47295 113226 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 113646 46816 113962 46817
rect 113646 46752 113652 46816
rect 113716 46752 113732 46816
rect 113796 46752 113812 46816
rect 113876 46752 113892 46816
rect 113956 46752 113962 46816
rect 113646 46751 113962 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 112910 46272 113226 46273
rect 112910 46208 112916 46272
rect 112980 46208 112996 46272
rect 113060 46208 113076 46272
rect 113140 46208 113156 46272
rect 113220 46208 113226 46272
rect 112910 46207 113226 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 113646 45728 113962 45729
rect 113646 45664 113652 45728
rect 113716 45664 113732 45728
rect 113796 45664 113812 45728
rect 113876 45664 113892 45728
rect 113956 45664 113962 45728
rect 113646 45663 113962 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 112910 45184 113226 45185
rect 112910 45120 112916 45184
rect 112980 45120 112996 45184
rect 113060 45120 113076 45184
rect 113140 45120 113156 45184
rect 113220 45120 113226 45184
rect 112910 45119 113226 45120
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 113646 44640 113962 44641
rect 113646 44576 113652 44640
rect 113716 44576 113732 44640
rect 113796 44576 113812 44640
rect 113876 44576 113892 44640
rect 113956 44576 113962 44640
rect 113646 44575 113962 44576
rect 0 44298 800 44328
rect 1301 44298 1367 44301
rect 0 44296 1367 44298
rect 0 44240 1306 44296
rect 1362 44240 1367 44296
rect 0 44238 1367 44240
rect 0 44208 800 44238
rect 1301 44235 1367 44238
rect 9673 44204 9739 44207
rect 9673 44202 10028 44204
rect 9673 44146 9678 44202
rect 9734 44146 10028 44202
rect 9673 44144 10028 44146
rect 9673 44141 9739 44144
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 112910 44096 113226 44097
rect 112910 44032 112916 44096
rect 112980 44032 112996 44096
rect 113060 44032 113076 44096
rect 113140 44032 113156 44096
rect 113220 44032 113226 44096
rect 112910 44031 113226 44032
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 113646 43552 113962 43553
rect 113646 43488 113652 43552
rect 113716 43488 113732 43552
rect 113796 43488 113812 43552
rect 113876 43488 113892 43552
rect 113956 43488 113962 43552
rect 113646 43487 113962 43488
rect 4210 43008 4526 43009
rect 0 42938 800 42968
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 112910 43008 113226 43009
rect 4210 42943 4526 42944
rect 9673 42980 9739 42983
rect 9673 42978 10028 42980
rect 1301 42938 1367 42941
rect 0 42936 1367 42938
rect 0 42880 1306 42936
rect 1362 42880 1367 42936
rect 9673 42922 9678 42978
rect 9734 42922 10028 42978
rect 112910 42944 112916 43008
rect 112980 42944 112996 43008
rect 113060 42944 113076 43008
rect 113140 42944 113156 43008
rect 113220 42944 113226 43008
rect 112910 42943 113226 42944
rect 9673 42920 10028 42922
rect 9673 42917 9739 42920
rect 0 42878 1367 42880
rect 0 42848 800 42878
rect 1301 42875 1367 42878
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 113646 42464 113962 42465
rect 113646 42400 113652 42464
rect 113716 42400 113732 42464
rect 113796 42400 113812 42464
rect 113876 42400 113892 42464
rect 113956 42400 113962 42464
rect 113646 42399 113962 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 112910 41920 113226 41921
rect 112910 41856 112916 41920
rect 112980 41856 112996 41920
rect 113060 41856 113076 41920
rect 113140 41856 113156 41920
rect 113220 41856 113226 41920
rect 112910 41855 113226 41856
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 113646 41376 113962 41377
rect 113646 41312 113652 41376
rect 113716 41312 113732 41376
rect 113796 41312 113812 41376
rect 113876 41312 113892 41376
rect 113956 41312 113962 41376
rect 113646 41311 113962 41312
rect 9673 41212 9739 41215
rect 9673 41210 10028 41212
rect 9673 41154 9678 41210
rect 9734 41154 10028 41210
rect 9673 41152 10028 41154
rect 9673 41149 9739 41152
rect 0 40898 800 40928
rect 1301 40898 1367 40901
rect 0 40896 1367 40898
rect 0 40840 1306 40896
rect 1362 40840 1367 40896
rect 0 40838 1367 40840
rect 0 40808 800 40838
rect 1301 40835 1367 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 112910 40832 113226 40833
rect 112910 40768 112916 40832
rect 112980 40768 112996 40832
rect 113060 40768 113076 40832
rect 113140 40768 113156 40832
rect 113220 40768 113226 40832
rect 112910 40767 113226 40768
rect 4870 40288 5186 40289
rect 0 40218 800 40248
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 113646 40288 113962 40289
rect 113646 40224 113652 40288
rect 113716 40224 113732 40288
rect 113796 40224 113812 40288
rect 113876 40224 113892 40288
rect 113956 40224 113962 40288
rect 113646 40223 113962 40224
rect 1301 40218 1367 40221
rect 0 40216 1367 40218
rect 0 40160 1306 40216
rect 1362 40160 1367 40216
rect 0 40158 1367 40160
rect 0 40128 800 40158
rect 1301 40155 1367 40158
rect 9673 40124 9739 40127
rect 9673 40122 10028 40124
rect 9673 40066 9678 40122
rect 9734 40066 10028 40122
rect 9673 40064 10028 40066
rect 9673 40061 9739 40064
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 112910 39744 113226 39745
rect 112910 39680 112916 39744
rect 112980 39680 112996 39744
rect 113060 39680 113076 39744
rect 113140 39680 113156 39744
rect 113220 39680 113226 39744
rect 112910 39679 113226 39680
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 113646 39200 113962 39201
rect 113646 39136 113652 39200
rect 113716 39136 113732 39200
rect 113796 39136 113812 39200
rect 113876 39136 113892 39200
rect 113956 39136 113962 39200
rect 113646 39135 113962 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 112910 38656 113226 38657
rect 112910 38592 112916 38656
rect 112980 38592 112996 38656
rect 113060 38592 113076 38656
rect 113140 38592 113156 38656
rect 113220 38592 113226 38656
rect 112910 38591 113226 38592
rect 9673 38492 9739 38495
rect 9673 38490 10028 38492
rect 9673 38434 9678 38490
rect 9734 38434 10028 38490
rect 9673 38432 10028 38434
rect 9673 38429 9739 38432
rect 0 38178 800 38208
rect 1209 38178 1275 38181
rect 0 38176 1275 38178
rect 0 38120 1214 38176
rect 1270 38120 1275 38176
rect 0 38118 1275 38120
rect 0 38088 800 38118
rect 1209 38115 1275 38118
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 113646 38112 113962 38113
rect 113646 38048 113652 38112
rect 113716 38048 113732 38112
rect 113796 38048 113812 38112
rect 113876 38048 113892 38112
rect 113956 38048 113962 38112
rect 113646 38047 113962 38048
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 112910 37568 113226 37569
rect 4210 37503 4526 37504
rect 9489 37540 9555 37543
rect 9489 37538 10028 37540
rect 1301 37498 1367 37501
rect 0 37496 1367 37498
rect 0 37440 1306 37496
rect 1362 37440 1367 37496
rect 9489 37482 9494 37538
rect 9550 37482 10028 37538
rect 112910 37504 112916 37568
rect 112980 37504 112996 37568
rect 113060 37504 113076 37568
rect 113140 37504 113156 37568
rect 113220 37504 113226 37568
rect 112910 37503 113226 37504
rect 9489 37480 10028 37482
rect 9489 37477 9555 37480
rect 0 37438 1367 37440
rect 0 37408 800 37438
rect 1301 37435 1367 37438
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 113646 37024 113962 37025
rect 113646 36960 113652 37024
rect 113716 36960 113732 37024
rect 113796 36960 113812 37024
rect 113876 36960 113892 37024
rect 113956 36960 113962 37024
rect 113646 36959 113962 36960
rect 113449 36818 113515 36821
rect 114001 36818 114067 36821
rect 115105 36818 115171 36821
rect 113449 36816 115171 36818
rect 113449 36760 113454 36816
rect 113510 36760 114006 36816
rect 114062 36760 115110 36816
rect 115166 36760 115171 36816
rect 113449 36758 115171 36760
rect 113449 36755 113515 36758
rect 114001 36755 114067 36758
rect 115105 36755 115171 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 112910 36480 113226 36481
rect 112910 36416 112916 36480
rect 112980 36416 112996 36480
rect 113060 36416 113076 36480
rect 113140 36416 113156 36480
rect 113220 36416 113226 36480
rect 112910 36415 113226 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 113646 35936 113962 35937
rect 113646 35872 113652 35936
rect 113716 35872 113732 35936
rect 113796 35872 113812 35936
rect 113876 35872 113892 35936
rect 113956 35872 113962 35936
rect 113646 35871 113962 35872
rect 9489 35772 9555 35775
rect 9489 35770 10028 35772
rect 9489 35714 9494 35770
rect 9550 35714 10028 35770
rect 9489 35712 10028 35714
rect 9489 35709 9555 35712
rect 0 35458 800 35488
rect 1301 35458 1367 35461
rect 0 35456 1367 35458
rect 0 35400 1306 35456
rect 1362 35400 1367 35456
rect 0 35398 1367 35400
rect 0 35368 800 35398
rect 1301 35395 1367 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 112910 35392 113226 35393
rect 112910 35328 112916 35392
rect 112980 35328 112996 35392
rect 113060 35328 113076 35392
rect 113140 35328 113156 35392
rect 113220 35328 113226 35392
rect 112910 35327 113226 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 113646 34848 113962 34849
rect 113646 34784 113652 34848
rect 113716 34784 113732 34848
rect 113796 34784 113812 34848
rect 113876 34784 113892 34848
rect 113956 34784 113962 34848
rect 113646 34783 113962 34784
rect 114093 34642 114159 34645
rect 115657 34642 115723 34645
rect 114093 34640 115723 34642
rect 114093 34584 114098 34640
rect 114154 34584 115662 34640
rect 115718 34584 115723 34640
rect 114093 34582 115723 34584
rect 114093 34579 114159 34582
rect 115657 34579 115723 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 112910 34304 113226 34305
rect 112910 34240 112916 34304
rect 112980 34240 112996 34304
rect 113060 34240 113076 34304
rect 113140 34240 113156 34304
rect 113220 34240 113226 34304
rect 112910 34239 113226 34240
rect 114921 33962 114987 33965
rect 115289 33962 115355 33965
rect 116117 33962 116183 33965
rect 114921 33960 116183 33962
rect 114921 33904 114926 33960
rect 114982 33904 115294 33960
rect 115350 33904 116122 33960
rect 116178 33904 116183 33960
rect 114921 33902 116183 33904
rect 114921 33899 114987 33902
rect 115289 33899 115355 33902
rect 116117 33899 116183 33902
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 113646 33760 113962 33761
rect 113646 33696 113652 33760
rect 113716 33696 113732 33760
rect 113796 33696 113812 33760
rect 113876 33696 113892 33760
rect 113956 33696 113962 33760
rect 113646 33695 113962 33696
rect 115841 33554 115907 33557
rect 116209 33554 116275 33557
rect 115841 33552 116275 33554
rect 115841 33496 115846 33552
rect 115902 33496 116214 33552
rect 116270 33496 116275 33552
rect 115841 33494 116275 33496
rect 115841 33491 115907 33494
rect 116209 33491 116275 33494
rect 109401 33284 109467 33285
rect 109350 33220 109356 33284
rect 109420 33282 109467 33284
rect 109420 33280 109512 33282
rect 109462 33224 109512 33280
rect 109420 33222 109512 33224
rect 109420 33220 109467 33222
rect 109401 33219 109467 33220
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 112910 33216 113226 33217
rect 112910 33152 112916 33216
rect 112980 33152 112996 33216
rect 113060 33152 113076 33216
rect 113140 33152 113156 33216
rect 113220 33152 113226 33216
rect 112910 33151 113226 33152
rect 115289 32874 115355 32877
rect 116485 32874 116551 32877
rect 115289 32872 116551 32874
rect 115289 32816 115294 32872
rect 115350 32816 116490 32872
rect 116546 32816 116551 32872
rect 115289 32814 116551 32816
rect 115289 32811 115355 32814
rect 116485 32811 116551 32814
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 113646 32672 113962 32673
rect 113646 32608 113652 32672
rect 113716 32608 113732 32672
rect 113796 32608 113812 32672
rect 113876 32608 113892 32672
rect 113956 32608 113962 32672
rect 113646 32607 113962 32608
rect 116761 32466 116827 32469
rect 117313 32466 117379 32469
rect 116761 32464 117379 32466
rect 116761 32408 116766 32464
rect 116822 32408 117318 32464
rect 117374 32408 117379 32464
rect 116761 32406 117379 32408
rect 116761 32403 116827 32406
rect 117313 32403 117379 32406
rect 116577 32330 116643 32333
rect 117497 32330 117563 32333
rect 116577 32328 117563 32330
rect 116577 32272 116582 32328
rect 116638 32272 117502 32328
rect 117558 32272 117563 32328
rect 116577 32270 117563 32272
rect 116577 32267 116643 32270
rect 117497 32267 117563 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 112910 32128 113226 32129
rect 112910 32064 112916 32128
rect 112980 32064 112996 32128
rect 113060 32064 113076 32128
rect 113140 32064 113156 32128
rect 113220 32064 113226 32128
rect 112910 32063 113226 32064
rect 118509 32058 118575 32061
rect 119200 32058 120000 32088
rect 118509 32056 120000 32058
rect 118509 32000 118514 32056
rect 118570 32000 120000 32056
rect 118509 31998 120000 32000
rect 118509 31995 118575 31998
rect 119200 31968 120000 31998
rect 114093 31922 114159 31925
rect 115749 31922 115815 31925
rect 114093 31920 115815 31922
rect 114093 31864 114098 31920
rect 114154 31864 115754 31920
rect 115810 31864 115815 31920
rect 114093 31862 115815 31864
rect 114093 31859 114159 31862
rect 115749 31859 115815 31862
rect 116117 31786 116183 31789
rect 117129 31786 117195 31789
rect 116117 31784 117195 31786
rect 116117 31728 116122 31784
rect 116178 31728 117134 31784
rect 117190 31728 117195 31784
rect 116117 31726 117195 31728
rect 116117 31723 116183 31726
rect 117129 31723 117195 31726
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 113646 31584 113962 31585
rect 113646 31520 113652 31584
rect 113716 31520 113732 31584
rect 113796 31520 113812 31584
rect 113876 31520 113892 31584
rect 113956 31520 113962 31584
rect 113646 31519 113962 31520
rect 118509 31378 118575 31381
rect 119200 31378 120000 31408
rect 118509 31376 120000 31378
rect 118509 31320 118514 31376
rect 118570 31320 120000 31376
rect 118509 31318 120000 31320
rect 118509 31315 118575 31318
rect 119200 31288 120000 31318
rect 111333 31242 111399 31245
rect 111885 31242 111951 31245
rect 111333 31240 111951 31242
rect 111333 31184 111338 31240
rect 111394 31184 111890 31240
rect 111946 31184 111951 31240
rect 111333 31182 111951 31184
rect 111333 31179 111399 31182
rect 111885 31179 111951 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 112910 31040 113226 31041
rect 112910 30976 112916 31040
rect 112980 30976 112996 31040
rect 113060 30976 113076 31040
rect 113140 30976 113156 31040
rect 113220 30976 113226 31040
rect 112910 30975 113226 30976
rect 112529 30834 112595 30837
rect 113081 30834 113147 30837
rect 114093 30834 114159 30837
rect 115105 30834 115171 30837
rect 112529 30832 115171 30834
rect 112529 30776 112534 30832
rect 112590 30776 113086 30832
rect 113142 30776 114098 30832
rect 114154 30776 115110 30832
rect 115166 30776 115171 30832
rect 112529 30774 115171 30776
rect 112529 30771 112595 30774
rect 113081 30771 113147 30774
rect 114093 30771 114159 30774
rect 115105 30771 115171 30774
rect 113817 30698 113883 30701
rect 114645 30698 114711 30701
rect 113817 30696 114711 30698
rect 113817 30640 113822 30696
rect 113878 30640 114650 30696
rect 114706 30640 114711 30696
rect 113817 30638 114711 30640
rect 113817 30635 113883 30638
rect 114645 30635 114711 30638
rect 118509 30698 118575 30701
rect 119200 30698 120000 30728
rect 118509 30696 120000 30698
rect 118509 30640 118514 30696
rect 118570 30640 120000 30696
rect 118509 30638 120000 30640
rect 118509 30635 118575 30638
rect 119200 30608 120000 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 113646 30496 113962 30497
rect 113646 30432 113652 30496
rect 113716 30432 113732 30496
rect 113796 30432 113812 30496
rect 113876 30432 113892 30496
rect 113956 30432 113962 30496
rect 113646 30431 113962 30432
rect 118601 30018 118667 30021
rect 119200 30018 120000 30048
rect 118601 30016 120000 30018
rect 118601 29960 118606 30016
rect 118662 29960 120000 30016
rect 118601 29958 120000 29960
rect 118601 29955 118667 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 112910 29952 113226 29953
rect 112910 29888 112916 29952
rect 112980 29888 112996 29952
rect 113060 29888 113076 29952
rect 113140 29888 113156 29952
rect 113220 29888 113226 29952
rect 119200 29928 120000 29958
rect 112910 29887 113226 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 113646 29408 113962 29409
rect 113646 29344 113652 29408
rect 113716 29344 113732 29408
rect 113796 29344 113812 29408
rect 113876 29344 113892 29408
rect 113956 29344 113962 29408
rect 113646 29343 113962 29344
rect 118233 29338 118299 29341
rect 119200 29338 120000 29368
rect 118233 29336 120000 29338
rect 118233 29280 118238 29336
rect 118294 29280 120000 29336
rect 118233 29278 120000 29280
rect 118233 29275 118299 29278
rect 119200 29248 120000 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 112910 28864 113226 28865
rect 112910 28800 112916 28864
rect 112980 28800 112996 28864
rect 113060 28800 113076 28864
rect 113140 28800 113156 28864
rect 113220 28800 113226 28864
rect 112910 28799 113226 28800
rect 117313 28658 117379 28661
rect 118509 28658 118575 28661
rect 119200 28658 120000 28688
rect 117313 28656 120000 28658
rect 117313 28600 117318 28656
rect 117374 28600 118514 28656
rect 118570 28600 120000 28656
rect 117313 28598 120000 28600
rect 117313 28595 117379 28598
rect 118509 28595 118575 28598
rect 119200 28568 120000 28598
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 113646 28320 113962 28321
rect 113646 28256 113652 28320
rect 113716 28256 113732 28320
rect 113796 28256 113812 28320
rect 113876 28256 113892 28320
rect 113956 28256 113962 28320
rect 113646 28255 113962 28256
rect 118233 27978 118299 27981
rect 119200 27978 120000 28008
rect 118233 27976 120000 27978
rect 118233 27920 118238 27976
rect 118294 27920 120000 27976
rect 118233 27918 120000 27920
rect 118233 27915 118299 27918
rect 119200 27888 120000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 112910 27776 113226 27777
rect 112910 27712 112916 27776
rect 112980 27712 112996 27776
rect 113060 27712 113076 27776
rect 113140 27712 113156 27776
rect 113220 27712 113226 27776
rect 112910 27711 113226 27712
rect 118509 27298 118575 27301
rect 119200 27298 120000 27328
rect 118509 27296 120000 27298
rect 118509 27240 118514 27296
rect 118570 27240 120000 27296
rect 118509 27238 120000 27240
rect 118509 27235 118575 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 113646 27232 113962 27233
rect 113646 27168 113652 27232
rect 113716 27168 113732 27232
rect 113796 27168 113812 27232
rect 113876 27168 113892 27232
rect 113956 27168 113962 27232
rect 119200 27208 120000 27238
rect 113646 27167 113962 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 112910 26688 113226 26689
rect 4210 26623 4526 26624
rect 105892 26618 106474 26660
rect 112910 26624 112916 26688
rect 112980 26624 112996 26688
rect 113060 26624 113076 26688
rect 113140 26624 113156 26688
rect 113220 26624 113226 26688
rect 112910 26623 113226 26624
rect 106917 26618 106983 26621
rect 105892 26616 106983 26618
rect 105892 26600 106922 26616
rect 106414 26560 106922 26600
rect 106978 26560 106983 26616
rect 106414 26558 106983 26560
rect 106917 26555 106983 26558
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 113646 26144 113962 26145
rect 113646 26080 113652 26144
rect 113716 26080 113732 26144
rect 113796 26080 113812 26144
rect 113876 26080 113892 26144
rect 113956 26080 113962 26144
rect 113646 26079 113962 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 112910 25600 113226 25601
rect 112910 25536 112916 25600
rect 112980 25536 112996 25600
rect 113060 25536 113076 25600
rect 113140 25536 113156 25600
rect 113220 25536 113226 25600
rect 112910 25535 113226 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 113646 25056 113962 25057
rect 4870 24991 5186 24992
rect 105892 24986 106474 25028
rect 113646 24992 113652 25056
rect 113716 24992 113732 25056
rect 113796 24992 113812 25056
rect 113876 24992 113892 25056
rect 113956 24992 113962 25056
rect 113646 24991 113962 24992
rect 107009 24986 107075 24989
rect 105892 24984 107075 24986
rect 105892 24968 107014 24984
rect 106414 24928 107014 24968
rect 107070 24928 107075 24984
rect 106414 24926 107075 24928
rect 107009 24923 107075 24926
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 112910 24512 113226 24513
rect 112910 24448 112916 24512
rect 112980 24448 112996 24512
rect 113060 24448 113076 24512
rect 113140 24448 113156 24512
rect 113220 24448 113226 24512
rect 112910 24447 113226 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 113646 23968 113962 23969
rect 113646 23904 113652 23968
rect 113716 23904 113732 23968
rect 113796 23904 113812 23968
rect 113876 23904 113892 23968
rect 113956 23904 113962 23968
rect 113646 23903 113962 23904
rect 105892 23626 106474 23668
rect 107101 23626 107167 23629
rect 105892 23624 107167 23626
rect 105892 23608 107106 23624
rect 106414 23568 107106 23608
rect 107162 23568 107167 23624
rect 106414 23566 107167 23568
rect 107101 23563 107167 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 112910 23424 113226 23425
rect 112910 23360 112916 23424
rect 112980 23360 112996 23424
rect 113060 23360 113076 23424
rect 113140 23360 113156 23424
rect 113220 23360 113226 23424
rect 112910 23359 113226 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 113646 22880 113962 22881
rect 113646 22816 113652 22880
rect 113716 22816 113732 22880
rect 113796 22816 113812 22880
rect 113876 22816 113892 22880
rect 113956 22816 113962 22880
rect 113646 22815 113962 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 112910 22336 113226 22337
rect 112910 22272 112916 22336
rect 112980 22272 112996 22336
rect 113060 22272 113076 22336
rect 113140 22272 113156 22336
rect 113220 22272 113226 22336
rect 112910 22271 113226 22272
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 113646 21792 113962 21793
rect 113646 21728 113652 21792
rect 113716 21728 113732 21792
rect 113796 21728 113812 21792
rect 113876 21728 113892 21792
rect 113956 21728 113962 21792
rect 113646 21727 113962 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 112910 21248 113226 21249
rect 112910 21184 112916 21248
rect 112980 21184 112996 21248
rect 113060 21184 113076 21248
rect 113140 21184 113156 21248
rect 113220 21184 113226 21248
rect 112910 21183 113226 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 113646 20704 113962 20705
rect 113646 20640 113652 20704
rect 113716 20640 113732 20704
rect 113796 20640 113812 20704
rect 113876 20640 113892 20704
rect 113956 20640 113962 20704
rect 113646 20639 113962 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 112910 20160 113226 20161
rect 112910 20096 112916 20160
rect 112980 20096 112996 20160
rect 113060 20096 113076 20160
rect 113140 20096 113156 20160
rect 113220 20096 113226 20160
rect 112910 20095 113226 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 113646 19616 113962 19617
rect 113646 19552 113652 19616
rect 113716 19552 113732 19616
rect 113796 19552 113812 19616
rect 113876 19552 113892 19616
rect 113956 19552 113962 19616
rect 113646 19551 113962 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 112910 19072 113226 19073
rect 112910 19008 112916 19072
rect 112980 19008 112996 19072
rect 113060 19008 113076 19072
rect 113140 19008 113156 19072
rect 113220 19008 113226 19072
rect 112910 19007 113226 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 113646 18528 113962 18529
rect 113646 18464 113652 18528
rect 113716 18464 113732 18528
rect 113796 18464 113812 18528
rect 113876 18464 113892 18528
rect 113956 18464 113962 18528
rect 113646 18463 113962 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 112910 17984 113226 17985
rect 112910 17920 112916 17984
rect 112980 17920 112996 17984
rect 113060 17920 113076 17984
rect 113140 17920 113156 17984
rect 113220 17920 113226 17984
rect 112910 17919 113226 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 113646 17440 113962 17441
rect 113646 17376 113652 17440
rect 113716 17376 113732 17440
rect 113796 17376 113812 17440
rect 113876 17376 113892 17440
rect 113956 17376 113962 17440
rect 113646 17375 113962 17376
rect 9673 17276 9739 17279
rect 9673 17274 10028 17276
rect 9673 17218 9678 17274
rect 9734 17218 10028 17274
rect 9673 17216 10028 17218
rect 9673 17213 9739 17216
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 112910 16896 113226 16897
rect 112910 16832 112916 16896
rect 112980 16832 112996 16896
rect 113060 16832 113076 16896
rect 113140 16832 113156 16896
rect 113220 16832 113226 16896
rect 112910 16831 113226 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 113646 16352 113962 16353
rect 113646 16288 113652 16352
rect 113716 16288 113732 16352
rect 113796 16288 113812 16352
rect 113876 16288 113892 16352
rect 113956 16288 113962 16352
rect 113646 16287 113962 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 112910 15808 113226 15809
rect 112910 15744 112916 15808
rect 112980 15744 112996 15808
rect 113060 15744 113076 15808
rect 113140 15744 113156 15808
rect 113220 15744 113226 15808
rect 112910 15743 113226 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 9673 15644 9739 15647
rect 9673 15642 10028 15644
rect 9673 15586 9678 15642
rect 9734 15586 10028 15642
rect 9673 15584 10028 15586
rect 9673 15581 9739 15584
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 113646 15264 113962 15265
rect 113646 15200 113652 15264
rect 113716 15200 113732 15264
rect 113796 15200 113812 15264
rect 113876 15200 113892 15264
rect 113956 15200 113962 15264
rect 113646 15199 113962 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 112910 14720 113226 14721
rect 112910 14656 112916 14720
rect 112980 14656 112996 14720
rect 113060 14656 113076 14720
rect 113140 14656 113156 14720
rect 113220 14656 113226 14720
rect 112910 14655 113226 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 113646 14176 113962 14177
rect 113646 14112 113652 14176
rect 113716 14112 113732 14176
rect 113796 14112 113812 14176
rect 113876 14112 113892 14176
rect 113956 14112 113962 14176
rect 113646 14111 113962 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 112910 13632 113226 13633
rect 112910 13568 112916 13632
rect 112980 13568 112996 13632
rect 113060 13568 113076 13632
rect 113140 13568 113156 13632
rect 113220 13568 113226 13632
rect 112910 13567 113226 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 113646 13088 113962 13089
rect 113646 13024 113652 13088
rect 113716 13024 113732 13088
rect 113796 13024 113812 13088
rect 113876 13024 113892 13088
rect 113956 13024 113962 13088
rect 113646 13023 113962 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 112910 12544 113226 12545
rect 112910 12480 112916 12544
rect 112980 12480 112996 12544
rect 113060 12480 113076 12544
rect 113140 12480 113156 12544
rect 113220 12480 113226 12544
rect 112910 12479 113226 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 113646 12000 113962 12001
rect 113646 11936 113652 12000
rect 113716 11936 113732 12000
rect 113796 11936 113812 12000
rect 113876 11936 113892 12000
rect 113956 11936 113962 12000
rect 113646 11935 113962 11936
rect 106457 11930 106523 11933
rect 109350 11930 109356 11932
rect 106457 11928 109356 11930
rect 106457 11872 106462 11928
rect 106518 11872 109356 11928
rect 106457 11870 109356 11872
rect 106457 11867 106523 11870
rect 109350 11868 109356 11870
rect 109420 11868 109426 11932
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 112910 11456 113226 11457
rect 112910 11392 112916 11456
rect 112980 11392 112996 11456
rect 113060 11392 113076 11456
rect 113140 11392 113156 11456
rect 113220 11392 113226 11456
rect 112910 11391 113226 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 113646 10912 113962 10913
rect 113646 10848 113652 10912
rect 113716 10848 113732 10912
rect 113796 10848 113812 10912
rect 113876 10848 113892 10912
rect 113956 10848 113962 10912
rect 113646 10847 113962 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 112910 10368 113226 10369
rect 112910 10304 112916 10368
rect 112980 10304 112996 10368
rect 113060 10304 113076 10368
rect 113140 10304 113156 10368
rect 113220 10304 113226 10368
rect 112910 10303 113226 10304
rect 93342 10026 93348 10028
rect 92968 9966 93348 10026
rect 15837 9892 15903 9893
rect 92749 9892 92815 9893
rect 92968 9892 93028 9966
rect 93342 9964 93348 9966
rect 93412 10026 93418 10028
rect 108757 10026 108823 10029
rect 93412 10024 108823 10026
rect 93412 9968 108762 10024
rect 108818 9968 108823 10024
rect 93412 9966 108823 9968
rect 93412 9964 93418 9966
rect 108757 9963 108823 9966
rect 15837 9888 15854 9892
rect 15918 9890 15924 9892
rect 92688 9890 92694 9892
rect 15837 9832 15842 9888
rect 15837 9828 15854 9832
rect 15918 9830 15994 9890
rect 92658 9830 92694 9890
rect 92758 9888 92815 9892
rect 92810 9832 92815 9888
rect 15918 9828 15924 9830
rect 92688 9828 92694 9830
rect 92758 9828 92815 9832
rect 92960 9828 92966 9892
rect 93030 9828 93036 9892
rect 93096 9828 93102 9892
rect 93166 9890 93172 9892
rect 93393 9890 93459 9893
rect 93166 9888 93459 9890
rect 93166 9832 93398 9888
rect 93454 9832 93459 9888
rect 93166 9830 93459 9832
rect 93166 9828 93172 9830
rect 15837 9827 15903 9828
rect 92749 9827 92815 9828
rect 93393 9827 93459 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 113646 9824 113962 9825
rect 113646 9760 113652 9824
rect 113716 9760 113732 9824
rect 113796 9760 113812 9824
rect 113876 9760 113892 9824
rect 113956 9760 113962 9824
rect 113646 9759 113962 9760
rect 26728 9692 26734 9756
rect 26798 9754 26804 9756
rect 26969 9754 27035 9757
rect 27797 9756 27863 9757
rect 27797 9754 27822 9756
rect 26798 9752 27035 9754
rect 26798 9696 26974 9752
rect 27030 9696 27035 9752
rect 26798 9694 27035 9696
rect 27730 9752 27822 9754
rect 27730 9696 27802 9752
rect 27730 9694 27822 9696
rect 26798 9692 26804 9694
rect 26969 9691 27035 9694
rect 27797 9692 27822 9694
rect 27886 9692 27892 9756
rect 29176 9692 29182 9756
rect 29246 9754 29252 9756
rect 29545 9754 29611 9757
rect 30189 9756 30255 9757
rect 29246 9752 29611 9754
rect 29246 9696 29550 9752
rect 29606 9696 29611 9752
rect 29246 9694 29611 9696
rect 29246 9692 29252 9694
rect 27797 9691 27863 9692
rect 29545 9691 29611 9694
rect 30128 9692 30134 9756
rect 30198 9754 30255 9756
rect 30198 9752 30290 9754
rect 30250 9696 30290 9752
rect 30198 9694 30290 9696
rect 30198 9692 30255 9694
rect 51344 9692 51350 9756
rect 51414 9754 51420 9756
rect 51625 9754 51691 9757
rect 52453 9756 52519 9757
rect 53557 9756 53623 9757
rect 52432 9754 52438 9756
rect 51414 9752 51691 9754
rect 51414 9696 51630 9752
rect 51686 9696 51691 9752
rect 51414 9694 51691 9696
rect 52362 9694 52438 9754
rect 52502 9752 52519 9756
rect 53520 9754 53526 9756
rect 52514 9696 52519 9752
rect 51414 9692 51420 9694
rect 30189 9691 30255 9692
rect 51625 9691 51691 9694
rect 52432 9692 52438 9694
rect 52502 9692 52519 9696
rect 53466 9694 53526 9754
rect 53590 9752 53623 9756
rect 53618 9696 53623 9752
rect 53520 9692 53526 9694
rect 53590 9692 53623 9696
rect 54880 9692 54886 9756
rect 54950 9754 54956 9756
rect 55029 9754 55095 9757
rect 54950 9752 55095 9754
rect 54950 9696 55034 9752
rect 55090 9696 55095 9752
rect 54950 9694 55095 9696
rect 54950 9692 54956 9694
rect 52453 9691 52519 9692
rect 53557 9691 53623 9692
rect 55029 9691 55095 9694
rect 55968 9692 55974 9756
rect 56038 9754 56044 9756
rect 56133 9754 56199 9757
rect 56038 9752 56199 9754
rect 56038 9696 56138 9752
rect 56194 9696 56199 9752
rect 56038 9694 56199 9696
rect 56038 9692 56044 9694
rect 56133 9691 56199 9694
rect 57056 9692 57062 9756
rect 57126 9754 57132 9756
rect 57421 9754 57487 9757
rect 57126 9752 57487 9754
rect 57126 9696 57426 9752
rect 57482 9696 57487 9752
rect 57126 9694 57487 9696
rect 57126 9692 57132 9694
rect 57421 9691 57487 9694
rect 58249 9756 58315 9757
rect 58249 9752 58286 9756
rect 58350 9754 58356 9756
rect 58249 9696 58254 9752
rect 58249 9692 58286 9696
rect 58350 9694 58406 9754
rect 58350 9692 58356 9694
rect 59368 9692 59374 9756
rect 59438 9754 59444 9756
rect 59537 9754 59603 9757
rect 60825 9756 60891 9757
rect 67725 9756 67791 9757
rect 60774 9754 60780 9756
rect 59438 9752 59603 9754
rect 59438 9696 59542 9752
rect 59598 9696 59603 9752
rect 59438 9694 59603 9696
rect 60734 9694 60780 9754
rect 60844 9752 60891 9756
rect 67664 9754 67670 9756
rect 60886 9696 60891 9752
rect 59438 9692 59444 9694
rect 58249 9691 58315 9692
rect 59537 9691 59603 9694
rect 60774 9692 60780 9694
rect 60844 9692 60891 9696
rect 67634 9694 67670 9754
rect 67734 9752 67791 9756
rect 67786 9696 67791 9752
rect 67664 9692 67670 9694
rect 67734 9692 67791 9696
rect 92824 9692 92830 9756
rect 92894 9754 92900 9756
rect 93025 9754 93091 9757
rect 92894 9752 93091 9754
rect 92894 9696 93030 9752
rect 93086 9696 93091 9752
rect 92894 9694 93091 9696
rect 92894 9692 92900 9694
rect 60825 9691 60891 9692
rect 67725 9691 67791 9692
rect 93025 9691 93091 9694
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 112910 9280 113226 9281
rect 112910 9216 112916 9280
rect 112980 9216 112996 9280
rect 113060 9216 113076 9280
rect 113140 9216 113156 9280
rect 113220 9216 113226 9280
rect 112910 9215 113226 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 113646 8736 113962 8737
rect 113646 8672 113652 8736
rect 113716 8672 113732 8736
rect 113796 8672 113812 8736
rect 113876 8672 113892 8736
rect 113956 8672 113962 8736
rect 113646 8671 113962 8672
rect 25446 8196 25452 8260
rect 25516 8258 25522 8260
rect 25865 8258 25931 8261
rect 25516 8256 25931 8258
rect 25516 8200 25870 8256
rect 25926 8200 25931 8256
rect 25516 8198 25931 8200
rect 25516 8196 25522 8198
rect 25865 8195 25931 8198
rect 31334 8196 31340 8260
rect 31404 8258 31410 8260
rect 31661 8258 31727 8261
rect 31404 8256 31727 8258
rect 31404 8200 31666 8256
rect 31722 8200 31727 8256
rect 31404 8198 31727 8200
rect 31404 8196 31410 8198
rect 31661 8195 31727 8198
rect 32622 8196 32628 8260
rect 32692 8258 32698 8260
rect 32949 8258 33015 8261
rect 33777 8260 33843 8261
rect 33726 8258 33732 8260
rect 32692 8256 33015 8258
rect 32692 8200 32954 8256
rect 33010 8200 33015 8256
rect 32692 8198 33015 8200
rect 33686 8198 33732 8258
rect 33796 8256 33843 8260
rect 33838 8200 33843 8256
rect 32692 8196 32698 8198
rect 32949 8195 33015 8198
rect 33726 8196 33732 8198
rect 33796 8196 33843 8200
rect 33777 8195 33843 8196
rect 34789 8258 34855 8261
rect 36169 8260 36235 8261
rect 35014 8258 35020 8260
rect 34789 8256 35020 8258
rect 34789 8200 34794 8256
rect 34850 8200 35020 8256
rect 34789 8198 35020 8200
rect 34789 8195 34855 8198
rect 35014 8196 35020 8198
rect 35084 8196 35090 8260
rect 36118 8258 36124 8260
rect 36078 8198 36124 8258
rect 36188 8256 36235 8260
rect 36230 8200 36235 8256
rect 36118 8196 36124 8198
rect 36188 8196 36235 8200
rect 37222 8196 37228 8260
rect 37292 8258 37298 8260
rect 37457 8258 37523 8261
rect 37292 8256 37523 8258
rect 37292 8200 37462 8256
rect 37518 8200 37523 8256
rect 37292 8198 37523 8200
rect 37292 8196 37298 8198
rect 36169 8195 36235 8196
rect 37457 8195 37523 8198
rect 38285 8260 38351 8261
rect 38285 8256 38332 8260
rect 38396 8258 38402 8260
rect 38285 8200 38290 8256
rect 38285 8196 38332 8200
rect 38396 8198 38442 8258
rect 38396 8196 38402 8198
rect 40718 8196 40724 8260
rect 40788 8258 40794 8260
rect 40861 8258 40927 8261
rect 40788 8256 40927 8258
rect 40788 8200 40866 8256
rect 40922 8200 40927 8256
rect 40788 8198 40927 8200
rect 40788 8196 40794 8198
rect 38285 8195 38351 8196
rect 40861 8195 40927 8198
rect 41822 8196 41828 8260
rect 41892 8258 41898 8260
rect 41965 8258 42031 8261
rect 41892 8256 42031 8258
rect 41892 8200 41970 8256
rect 42026 8200 42031 8256
rect 41892 8198 42031 8200
rect 41892 8196 41898 8198
rect 41965 8195 42031 8198
rect 43110 8196 43116 8260
rect 43180 8258 43186 8260
rect 43253 8258 43319 8261
rect 43180 8256 43319 8258
rect 43180 8200 43258 8256
rect 43314 8200 43319 8256
rect 43180 8198 43319 8200
rect 43180 8196 43186 8198
rect 43253 8195 43319 8198
rect 44214 8196 44220 8260
rect 44284 8258 44290 8260
rect 44541 8258 44607 8261
rect 46657 8260 46723 8261
rect 47761 8260 47827 8261
rect 49049 8260 49115 8261
rect 50337 8260 50403 8261
rect 61929 8260 61995 8261
rect 46606 8258 46612 8260
rect 44284 8256 44607 8258
rect 44284 8200 44546 8256
rect 44602 8200 44607 8256
rect 44284 8198 44607 8200
rect 46566 8198 46612 8258
rect 46676 8256 46723 8260
rect 47710 8258 47716 8260
rect 46718 8200 46723 8256
rect 44284 8196 44290 8198
rect 44541 8195 44607 8198
rect 46606 8196 46612 8198
rect 46676 8196 46723 8200
rect 47670 8198 47716 8258
rect 47780 8256 47827 8260
rect 48998 8258 49004 8260
rect 47822 8200 47827 8256
rect 47710 8196 47716 8198
rect 47780 8196 47827 8200
rect 48958 8198 49004 8258
rect 49068 8256 49115 8260
rect 50286 8258 50292 8260
rect 49110 8200 49115 8256
rect 48998 8196 49004 8198
rect 49068 8196 49115 8200
rect 50246 8198 50292 8258
rect 50356 8256 50403 8260
rect 61878 8258 61884 8260
rect 50398 8200 50403 8256
rect 50286 8196 50292 8198
rect 50356 8196 50403 8200
rect 61838 8198 61884 8258
rect 61948 8256 61995 8260
rect 61990 8200 61995 8256
rect 61878 8196 61884 8198
rect 61948 8196 61995 8200
rect 62982 8196 62988 8260
rect 63052 8258 63058 8260
rect 63217 8258 63283 8261
rect 63052 8256 63283 8258
rect 63052 8200 63222 8256
rect 63278 8200 63283 8256
rect 63052 8198 63283 8200
rect 63052 8196 63058 8198
rect 46657 8195 46723 8196
rect 47761 8195 47827 8196
rect 49049 8195 49115 8196
rect 50337 8195 50403 8196
rect 61929 8195 61995 8196
rect 63217 8195 63283 8198
rect 64045 8260 64111 8261
rect 64045 8256 64092 8260
rect 64156 8258 64162 8260
rect 64045 8200 64050 8256
rect 64045 8196 64092 8200
rect 64156 8198 64202 8258
rect 64156 8196 64162 8198
rect 65190 8196 65196 8260
rect 65260 8258 65266 8260
rect 65333 8258 65399 8261
rect 66713 8260 66779 8261
rect 66662 8258 66668 8260
rect 65260 8256 65399 8258
rect 65260 8200 65338 8256
rect 65394 8200 65399 8256
rect 65260 8198 65399 8200
rect 66622 8198 66668 8258
rect 66732 8256 66779 8260
rect 66774 8200 66779 8256
rect 65260 8196 65266 8198
rect 64045 8195 64111 8196
rect 65333 8195 65399 8198
rect 66662 8196 66668 8198
rect 66732 8196 66779 8200
rect 66713 8195 66779 8196
rect 93209 8258 93275 8261
rect 93342 8258 93348 8260
rect 93209 8256 93348 8258
rect 93209 8200 93214 8256
rect 93270 8200 93348 8256
rect 93209 8198 93348 8200
rect 93209 8195 93275 8198
rect 93342 8196 93348 8198
rect 93412 8196 93418 8260
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 112910 8192 113226 8193
rect 112910 8128 112916 8192
rect 112980 8128 112996 8192
rect 113060 8128 113076 8192
rect 113140 8128 113156 8192
rect 113220 8128 113226 8192
rect 112910 8127 113226 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 66310 7648 66626 7649
rect 66310 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66626 7648
rect 66310 7583 66626 7584
rect 97030 7648 97346 7649
rect 97030 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97346 7648
rect 97030 7583 97346 7584
rect 113646 7648 113962 7649
rect 113646 7584 113652 7648
rect 113716 7584 113732 7648
rect 113796 7584 113812 7648
rect 113876 7584 113892 7648
rect 113956 7584 113962 7648
rect 113646 7583 113962 7584
rect 45502 7108 45508 7172
rect 45572 7170 45578 7172
rect 45829 7170 45895 7173
rect 45572 7168 45895 7170
rect 45572 7112 45834 7168
rect 45890 7112 45895 7168
rect 45572 7110 45895 7112
rect 45572 7108 45578 7110
rect 45829 7107 45895 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 96370 7104 96686 7105
rect 96370 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96686 7104
rect 96370 7039 96686 7040
rect 112910 7104 113226 7105
rect 112910 7040 112916 7104
rect 112980 7040 112996 7104
rect 113060 7040 113076 7104
rect 113140 7040 113156 7104
rect 113220 7040 113226 7104
rect 112910 7039 113226 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 66310 6560 66626 6561
rect 66310 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66626 6560
rect 66310 6495 66626 6496
rect 97030 6560 97346 6561
rect 97030 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97346 6560
rect 97030 6495 97346 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 96370 6016 96686 6017
rect 96370 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96686 6016
rect 96370 5951 96686 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 66310 5472 66626 5473
rect 66310 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66626 5472
rect 66310 5407 66626 5408
rect 97030 5472 97346 5473
rect 97030 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97346 5472
rect 97030 5407 97346 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 96370 4928 96686 4929
rect 96370 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96686 4928
rect 96370 4863 96686 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 66310 4384 66626 4385
rect 66310 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66626 4384
rect 66310 4319 66626 4320
rect 97030 4384 97346 4385
rect 97030 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97346 4384
rect 97030 4319 97346 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 96370 3840 96686 3841
rect 96370 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96686 3840
rect 96370 3775 96686 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 66310 3296 66626 3297
rect 66310 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66626 3296
rect 66310 3231 66626 3232
rect 97030 3296 97346 3297
rect 97030 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97346 3296
rect 97030 3231 97346 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 96370 2752 96686 2753
rect 96370 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96686 2752
rect 96370 2687 96686 2688
rect 39614 2620 39620 2684
rect 39684 2682 39690 2684
rect 40033 2682 40099 2685
rect 39684 2680 40099 2682
rect 39684 2624 40038 2680
rect 40094 2624 40099 2680
rect 39684 2622 40099 2624
rect 39684 2620 39690 2622
rect 40033 2619 40099 2622
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 66310 2208 66626 2209
rect 66310 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66626 2208
rect 66310 2143 66626 2144
rect 97030 2208 97346 2209
rect 97030 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97346 2208
rect 97030 2143 97346 2144
<< via3 >>
rect 4216 97404 4280 97408
rect 4216 97348 4220 97404
rect 4220 97348 4276 97404
rect 4276 97348 4280 97404
rect 4216 97344 4280 97348
rect 4296 97404 4360 97408
rect 4296 97348 4300 97404
rect 4300 97348 4356 97404
rect 4356 97348 4360 97404
rect 4296 97344 4360 97348
rect 4376 97404 4440 97408
rect 4376 97348 4380 97404
rect 4380 97348 4436 97404
rect 4436 97348 4440 97404
rect 4376 97344 4440 97348
rect 4456 97404 4520 97408
rect 4456 97348 4460 97404
rect 4460 97348 4516 97404
rect 4516 97348 4520 97404
rect 4456 97344 4520 97348
rect 34936 97404 35000 97408
rect 34936 97348 34940 97404
rect 34940 97348 34996 97404
rect 34996 97348 35000 97404
rect 34936 97344 35000 97348
rect 35016 97404 35080 97408
rect 35016 97348 35020 97404
rect 35020 97348 35076 97404
rect 35076 97348 35080 97404
rect 35016 97344 35080 97348
rect 35096 97404 35160 97408
rect 35096 97348 35100 97404
rect 35100 97348 35156 97404
rect 35156 97348 35160 97404
rect 35096 97344 35160 97348
rect 35176 97404 35240 97408
rect 35176 97348 35180 97404
rect 35180 97348 35236 97404
rect 35236 97348 35240 97404
rect 35176 97344 35240 97348
rect 65656 97404 65720 97408
rect 65656 97348 65660 97404
rect 65660 97348 65716 97404
rect 65716 97348 65720 97404
rect 65656 97344 65720 97348
rect 65736 97404 65800 97408
rect 65736 97348 65740 97404
rect 65740 97348 65796 97404
rect 65796 97348 65800 97404
rect 65736 97344 65800 97348
rect 65816 97404 65880 97408
rect 65816 97348 65820 97404
rect 65820 97348 65876 97404
rect 65876 97348 65880 97404
rect 65816 97344 65880 97348
rect 65896 97404 65960 97408
rect 65896 97348 65900 97404
rect 65900 97348 65956 97404
rect 65956 97348 65960 97404
rect 65896 97344 65960 97348
rect 96376 97404 96440 97408
rect 96376 97348 96380 97404
rect 96380 97348 96436 97404
rect 96436 97348 96440 97404
rect 96376 97344 96440 97348
rect 96456 97404 96520 97408
rect 96456 97348 96460 97404
rect 96460 97348 96516 97404
rect 96516 97348 96520 97404
rect 96456 97344 96520 97348
rect 96536 97404 96600 97408
rect 96536 97348 96540 97404
rect 96540 97348 96596 97404
rect 96596 97348 96600 97404
rect 96536 97344 96600 97348
rect 96616 97404 96680 97408
rect 96616 97348 96620 97404
rect 96620 97348 96676 97404
rect 96676 97348 96680 97404
rect 96616 97344 96680 97348
rect 4876 96860 4940 96864
rect 4876 96804 4880 96860
rect 4880 96804 4936 96860
rect 4936 96804 4940 96860
rect 4876 96800 4940 96804
rect 4956 96860 5020 96864
rect 4956 96804 4960 96860
rect 4960 96804 5016 96860
rect 5016 96804 5020 96860
rect 4956 96800 5020 96804
rect 5036 96860 5100 96864
rect 5036 96804 5040 96860
rect 5040 96804 5096 96860
rect 5096 96804 5100 96860
rect 5036 96800 5100 96804
rect 5116 96860 5180 96864
rect 5116 96804 5120 96860
rect 5120 96804 5176 96860
rect 5176 96804 5180 96860
rect 5116 96800 5180 96804
rect 35596 96860 35660 96864
rect 35596 96804 35600 96860
rect 35600 96804 35656 96860
rect 35656 96804 35660 96860
rect 35596 96800 35660 96804
rect 35676 96860 35740 96864
rect 35676 96804 35680 96860
rect 35680 96804 35736 96860
rect 35736 96804 35740 96860
rect 35676 96800 35740 96804
rect 35756 96860 35820 96864
rect 35756 96804 35760 96860
rect 35760 96804 35816 96860
rect 35816 96804 35820 96860
rect 35756 96800 35820 96804
rect 35836 96860 35900 96864
rect 35836 96804 35840 96860
rect 35840 96804 35896 96860
rect 35896 96804 35900 96860
rect 35836 96800 35900 96804
rect 66316 96860 66380 96864
rect 66316 96804 66320 96860
rect 66320 96804 66376 96860
rect 66376 96804 66380 96860
rect 66316 96800 66380 96804
rect 66396 96860 66460 96864
rect 66396 96804 66400 96860
rect 66400 96804 66456 96860
rect 66456 96804 66460 96860
rect 66396 96800 66460 96804
rect 66476 96860 66540 96864
rect 66476 96804 66480 96860
rect 66480 96804 66536 96860
rect 66536 96804 66540 96860
rect 66476 96800 66540 96804
rect 66556 96860 66620 96864
rect 66556 96804 66560 96860
rect 66560 96804 66616 96860
rect 66616 96804 66620 96860
rect 66556 96800 66620 96804
rect 97036 96860 97100 96864
rect 97036 96804 97040 96860
rect 97040 96804 97096 96860
rect 97096 96804 97100 96860
rect 97036 96800 97100 96804
rect 97116 96860 97180 96864
rect 97116 96804 97120 96860
rect 97120 96804 97176 96860
rect 97176 96804 97180 96860
rect 97116 96800 97180 96804
rect 97196 96860 97260 96864
rect 97196 96804 97200 96860
rect 97200 96804 97256 96860
rect 97256 96804 97260 96860
rect 97196 96800 97260 96804
rect 97276 96860 97340 96864
rect 97276 96804 97280 96860
rect 97280 96804 97336 96860
rect 97336 96804 97340 96860
rect 97276 96800 97340 96804
rect 4216 96316 4280 96320
rect 4216 96260 4220 96316
rect 4220 96260 4276 96316
rect 4276 96260 4280 96316
rect 4216 96256 4280 96260
rect 4296 96316 4360 96320
rect 4296 96260 4300 96316
rect 4300 96260 4356 96316
rect 4356 96260 4360 96316
rect 4296 96256 4360 96260
rect 4376 96316 4440 96320
rect 4376 96260 4380 96316
rect 4380 96260 4436 96316
rect 4436 96260 4440 96316
rect 4376 96256 4440 96260
rect 4456 96316 4520 96320
rect 4456 96260 4460 96316
rect 4460 96260 4516 96316
rect 4516 96260 4520 96316
rect 4456 96256 4520 96260
rect 34936 96316 35000 96320
rect 34936 96260 34940 96316
rect 34940 96260 34996 96316
rect 34996 96260 35000 96316
rect 34936 96256 35000 96260
rect 35016 96316 35080 96320
rect 35016 96260 35020 96316
rect 35020 96260 35076 96316
rect 35076 96260 35080 96316
rect 35016 96256 35080 96260
rect 35096 96316 35160 96320
rect 35096 96260 35100 96316
rect 35100 96260 35156 96316
rect 35156 96260 35160 96316
rect 35096 96256 35160 96260
rect 35176 96316 35240 96320
rect 35176 96260 35180 96316
rect 35180 96260 35236 96316
rect 35236 96260 35240 96316
rect 35176 96256 35240 96260
rect 65656 96316 65720 96320
rect 65656 96260 65660 96316
rect 65660 96260 65716 96316
rect 65716 96260 65720 96316
rect 65656 96256 65720 96260
rect 65736 96316 65800 96320
rect 65736 96260 65740 96316
rect 65740 96260 65796 96316
rect 65796 96260 65800 96316
rect 65736 96256 65800 96260
rect 65816 96316 65880 96320
rect 65816 96260 65820 96316
rect 65820 96260 65876 96316
rect 65876 96260 65880 96316
rect 65816 96256 65880 96260
rect 65896 96316 65960 96320
rect 65896 96260 65900 96316
rect 65900 96260 65956 96316
rect 65956 96260 65960 96316
rect 65896 96256 65960 96260
rect 96376 96316 96440 96320
rect 96376 96260 96380 96316
rect 96380 96260 96436 96316
rect 96436 96260 96440 96316
rect 96376 96256 96440 96260
rect 96456 96316 96520 96320
rect 96456 96260 96460 96316
rect 96460 96260 96516 96316
rect 96516 96260 96520 96316
rect 96456 96256 96520 96260
rect 96536 96316 96600 96320
rect 96536 96260 96540 96316
rect 96540 96260 96596 96316
rect 96596 96260 96600 96316
rect 96536 96256 96600 96260
rect 96616 96316 96680 96320
rect 96616 96260 96620 96316
rect 96620 96260 96676 96316
rect 96676 96260 96680 96316
rect 96616 96256 96680 96260
rect 4876 95772 4940 95776
rect 4876 95716 4880 95772
rect 4880 95716 4936 95772
rect 4936 95716 4940 95772
rect 4876 95712 4940 95716
rect 4956 95772 5020 95776
rect 4956 95716 4960 95772
rect 4960 95716 5016 95772
rect 5016 95716 5020 95772
rect 4956 95712 5020 95716
rect 5036 95772 5100 95776
rect 5036 95716 5040 95772
rect 5040 95716 5096 95772
rect 5096 95716 5100 95772
rect 5036 95712 5100 95716
rect 5116 95772 5180 95776
rect 5116 95716 5120 95772
rect 5120 95716 5176 95772
rect 5176 95716 5180 95772
rect 5116 95712 5180 95716
rect 35596 95772 35660 95776
rect 35596 95716 35600 95772
rect 35600 95716 35656 95772
rect 35656 95716 35660 95772
rect 35596 95712 35660 95716
rect 35676 95772 35740 95776
rect 35676 95716 35680 95772
rect 35680 95716 35736 95772
rect 35736 95716 35740 95772
rect 35676 95712 35740 95716
rect 35756 95772 35820 95776
rect 35756 95716 35760 95772
rect 35760 95716 35816 95772
rect 35816 95716 35820 95772
rect 35756 95712 35820 95716
rect 35836 95772 35900 95776
rect 35836 95716 35840 95772
rect 35840 95716 35896 95772
rect 35896 95716 35900 95772
rect 35836 95712 35900 95716
rect 66316 95772 66380 95776
rect 66316 95716 66320 95772
rect 66320 95716 66376 95772
rect 66376 95716 66380 95772
rect 66316 95712 66380 95716
rect 66396 95772 66460 95776
rect 66396 95716 66400 95772
rect 66400 95716 66456 95772
rect 66456 95716 66460 95772
rect 66396 95712 66460 95716
rect 66476 95772 66540 95776
rect 66476 95716 66480 95772
rect 66480 95716 66536 95772
rect 66536 95716 66540 95772
rect 66476 95712 66540 95716
rect 66556 95772 66620 95776
rect 66556 95716 66560 95772
rect 66560 95716 66616 95772
rect 66616 95716 66620 95772
rect 66556 95712 66620 95716
rect 97036 95772 97100 95776
rect 97036 95716 97040 95772
rect 97040 95716 97096 95772
rect 97096 95716 97100 95772
rect 97036 95712 97100 95716
rect 97116 95772 97180 95776
rect 97116 95716 97120 95772
rect 97120 95716 97176 95772
rect 97176 95716 97180 95772
rect 97116 95712 97180 95716
rect 97196 95772 97260 95776
rect 97196 95716 97200 95772
rect 97200 95716 97256 95772
rect 97256 95716 97260 95772
rect 97196 95712 97260 95716
rect 97276 95772 97340 95776
rect 97276 95716 97280 95772
rect 97280 95716 97336 95772
rect 97336 95716 97340 95772
rect 97276 95712 97340 95716
rect 4216 95228 4280 95232
rect 4216 95172 4220 95228
rect 4220 95172 4276 95228
rect 4276 95172 4280 95228
rect 4216 95168 4280 95172
rect 4296 95228 4360 95232
rect 4296 95172 4300 95228
rect 4300 95172 4356 95228
rect 4356 95172 4360 95228
rect 4296 95168 4360 95172
rect 4376 95228 4440 95232
rect 4376 95172 4380 95228
rect 4380 95172 4436 95228
rect 4436 95172 4440 95228
rect 4376 95168 4440 95172
rect 4456 95228 4520 95232
rect 4456 95172 4460 95228
rect 4460 95172 4516 95228
rect 4516 95172 4520 95228
rect 4456 95168 4520 95172
rect 34936 95228 35000 95232
rect 34936 95172 34940 95228
rect 34940 95172 34996 95228
rect 34996 95172 35000 95228
rect 34936 95168 35000 95172
rect 35016 95228 35080 95232
rect 35016 95172 35020 95228
rect 35020 95172 35076 95228
rect 35076 95172 35080 95228
rect 35016 95168 35080 95172
rect 35096 95228 35160 95232
rect 35096 95172 35100 95228
rect 35100 95172 35156 95228
rect 35156 95172 35160 95228
rect 35096 95168 35160 95172
rect 35176 95228 35240 95232
rect 35176 95172 35180 95228
rect 35180 95172 35236 95228
rect 35236 95172 35240 95228
rect 35176 95168 35240 95172
rect 65656 95228 65720 95232
rect 65656 95172 65660 95228
rect 65660 95172 65716 95228
rect 65716 95172 65720 95228
rect 65656 95168 65720 95172
rect 65736 95228 65800 95232
rect 65736 95172 65740 95228
rect 65740 95172 65796 95228
rect 65796 95172 65800 95228
rect 65736 95168 65800 95172
rect 65816 95228 65880 95232
rect 65816 95172 65820 95228
rect 65820 95172 65876 95228
rect 65876 95172 65880 95228
rect 65816 95168 65880 95172
rect 65896 95228 65960 95232
rect 65896 95172 65900 95228
rect 65900 95172 65956 95228
rect 65956 95172 65960 95228
rect 65896 95168 65960 95172
rect 96376 95228 96440 95232
rect 96376 95172 96380 95228
rect 96380 95172 96436 95228
rect 96436 95172 96440 95228
rect 96376 95168 96440 95172
rect 96456 95228 96520 95232
rect 96456 95172 96460 95228
rect 96460 95172 96516 95228
rect 96516 95172 96520 95228
rect 96456 95168 96520 95172
rect 96536 95228 96600 95232
rect 96536 95172 96540 95228
rect 96540 95172 96596 95228
rect 96596 95172 96600 95228
rect 96536 95168 96600 95172
rect 96616 95228 96680 95232
rect 96616 95172 96620 95228
rect 96620 95172 96676 95228
rect 96676 95172 96680 95228
rect 96616 95168 96680 95172
rect 4876 94684 4940 94688
rect 4876 94628 4880 94684
rect 4880 94628 4936 94684
rect 4936 94628 4940 94684
rect 4876 94624 4940 94628
rect 4956 94684 5020 94688
rect 4956 94628 4960 94684
rect 4960 94628 5016 94684
rect 5016 94628 5020 94684
rect 4956 94624 5020 94628
rect 5036 94684 5100 94688
rect 5036 94628 5040 94684
rect 5040 94628 5096 94684
rect 5096 94628 5100 94684
rect 5036 94624 5100 94628
rect 5116 94684 5180 94688
rect 5116 94628 5120 94684
rect 5120 94628 5176 94684
rect 5176 94628 5180 94684
rect 5116 94624 5180 94628
rect 35596 94684 35660 94688
rect 35596 94628 35600 94684
rect 35600 94628 35656 94684
rect 35656 94628 35660 94684
rect 35596 94624 35660 94628
rect 35676 94684 35740 94688
rect 35676 94628 35680 94684
rect 35680 94628 35736 94684
rect 35736 94628 35740 94684
rect 35676 94624 35740 94628
rect 35756 94684 35820 94688
rect 35756 94628 35760 94684
rect 35760 94628 35816 94684
rect 35816 94628 35820 94684
rect 35756 94624 35820 94628
rect 35836 94684 35900 94688
rect 35836 94628 35840 94684
rect 35840 94628 35896 94684
rect 35896 94628 35900 94684
rect 35836 94624 35900 94628
rect 66316 94684 66380 94688
rect 66316 94628 66320 94684
rect 66320 94628 66376 94684
rect 66376 94628 66380 94684
rect 66316 94624 66380 94628
rect 66396 94684 66460 94688
rect 66396 94628 66400 94684
rect 66400 94628 66456 94684
rect 66456 94628 66460 94684
rect 66396 94624 66460 94628
rect 66476 94684 66540 94688
rect 66476 94628 66480 94684
rect 66480 94628 66536 94684
rect 66536 94628 66540 94684
rect 66476 94624 66540 94628
rect 66556 94684 66620 94688
rect 66556 94628 66560 94684
rect 66560 94628 66616 94684
rect 66616 94628 66620 94684
rect 66556 94624 66620 94628
rect 97036 94684 97100 94688
rect 97036 94628 97040 94684
rect 97040 94628 97096 94684
rect 97096 94628 97100 94684
rect 97036 94624 97100 94628
rect 97116 94684 97180 94688
rect 97116 94628 97120 94684
rect 97120 94628 97176 94684
rect 97176 94628 97180 94684
rect 97116 94624 97180 94628
rect 97196 94684 97260 94688
rect 97196 94628 97200 94684
rect 97200 94628 97256 94684
rect 97256 94628 97260 94684
rect 97196 94624 97260 94628
rect 97276 94684 97340 94688
rect 97276 94628 97280 94684
rect 97280 94628 97336 94684
rect 97336 94628 97340 94684
rect 97276 94624 97340 94628
rect 4216 94140 4280 94144
rect 4216 94084 4220 94140
rect 4220 94084 4276 94140
rect 4276 94084 4280 94140
rect 4216 94080 4280 94084
rect 4296 94140 4360 94144
rect 4296 94084 4300 94140
rect 4300 94084 4356 94140
rect 4356 94084 4360 94140
rect 4296 94080 4360 94084
rect 4376 94140 4440 94144
rect 4376 94084 4380 94140
rect 4380 94084 4436 94140
rect 4436 94084 4440 94140
rect 4376 94080 4440 94084
rect 4456 94140 4520 94144
rect 4456 94084 4460 94140
rect 4460 94084 4516 94140
rect 4516 94084 4520 94140
rect 4456 94080 4520 94084
rect 34936 94140 35000 94144
rect 34936 94084 34940 94140
rect 34940 94084 34996 94140
rect 34996 94084 35000 94140
rect 34936 94080 35000 94084
rect 35016 94140 35080 94144
rect 35016 94084 35020 94140
rect 35020 94084 35076 94140
rect 35076 94084 35080 94140
rect 35016 94080 35080 94084
rect 35096 94140 35160 94144
rect 35096 94084 35100 94140
rect 35100 94084 35156 94140
rect 35156 94084 35160 94140
rect 35096 94080 35160 94084
rect 35176 94140 35240 94144
rect 35176 94084 35180 94140
rect 35180 94084 35236 94140
rect 35236 94084 35240 94140
rect 35176 94080 35240 94084
rect 65656 94140 65720 94144
rect 65656 94084 65660 94140
rect 65660 94084 65716 94140
rect 65716 94084 65720 94140
rect 65656 94080 65720 94084
rect 65736 94140 65800 94144
rect 65736 94084 65740 94140
rect 65740 94084 65796 94140
rect 65796 94084 65800 94140
rect 65736 94080 65800 94084
rect 65816 94140 65880 94144
rect 65816 94084 65820 94140
rect 65820 94084 65876 94140
rect 65876 94084 65880 94140
rect 65816 94080 65880 94084
rect 65896 94140 65960 94144
rect 65896 94084 65900 94140
rect 65900 94084 65956 94140
rect 65956 94084 65960 94140
rect 65896 94080 65960 94084
rect 96376 94140 96440 94144
rect 96376 94084 96380 94140
rect 96380 94084 96436 94140
rect 96436 94084 96440 94140
rect 96376 94080 96440 94084
rect 96456 94140 96520 94144
rect 96456 94084 96460 94140
rect 96460 94084 96516 94140
rect 96516 94084 96520 94140
rect 96456 94080 96520 94084
rect 96536 94140 96600 94144
rect 96536 94084 96540 94140
rect 96540 94084 96596 94140
rect 96596 94084 96600 94140
rect 96536 94080 96600 94084
rect 96616 94140 96680 94144
rect 96616 94084 96620 94140
rect 96620 94084 96676 94140
rect 96676 94084 96680 94140
rect 96616 94080 96680 94084
rect 49372 93876 49436 93940
rect 4876 93596 4940 93600
rect 4876 93540 4880 93596
rect 4880 93540 4936 93596
rect 4936 93540 4940 93596
rect 4876 93536 4940 93540
rect 4956 93596 5020 93600
rect 4956 93540 4960 93596
rect 4960 93540 5016 93596
rect 5016 93540 5020 93596
rect 4956 93536 5020 93540
rect 5036 93596 5100 93600
rect 5036 93540 5040 93596
rect 5040 93540 5096 93596
rect 5096 93540 5100 93596
rect 5036 93536 5100 93540
rect 5116 93596 5180 93600
rect 5116 93540 5120 93596
rect 5120 93540 5176 93596
rect 5176 93540 5180 93596
rect 5116 93536 5180 93540
rect 35596 93596 35660 93600
rect 35596 93540 35600 93596
rect 35600 93540 35656 93596
rect 35656 93540 35660 93596
rect 35596 93536 35660 93540
rect 35676 93596 35740 93600
rect 35676 93540 35680 93596
rect 35680 93540 35736 93596
rect 35736 93540 35740 93596
rect 35676 93536 35740 93540
rect 35756 93596 35820 93600
rect 35756 93540 35760 93596
rect 35760 93540 35816 93596
rect 35816 93540 35820 93596
rect 35756 93536 35820 93540
rect 35836 93596 35900 93600
rect 35836 93540 35840 93596
rect 35840 93540 35896 93596
rect 35896 93540 35900 93596
rect 35836 93536 35900 93540
rect 66316 93596 66380 93600
rect 66316 93540 66320 93596
rect 66320 93540 66376 93596
rect 66376 93540 66380 93596
rect 66316 93536 66380 93540
rect 66396 93596 66460 93600
rect 66396 93540 66400 93596
rect 66400 93540 66456 93596
rect 66456 93540 66460 93596
rect 66396 93536 66460 93540
rect 66476 93596 66540 93600
rect 66476 93540 66480 93596
rect 66480 93540 66536 93596
rect 66536 93540 66540 93596
rect 66476 93536 66540 93540
rect 66556 93596 66620 93600
rect 66556 93540 66560 93596
rect 66560 93540 66616 93596
rect 66616 93540 66620 93596
rect 66556 93536 66620 93540
rect 97036 93596 97100 93600
rect 97036 93540 97040 93596
rect 97040 93540 97096 93596
rect 97096 93540 97100 93596
rect 97036 93536 97100 93540
rect 97116 93596 97180 93600
rect 97116 93540 97120 93596
rect 97120 93540 97176 93596
rect 97176 93540 97180 93596
rect 97116 93536 97180 93540
rect 97196 93596 97260 93600
rect 97196 93540 97200 93596
rect 97200 93540 97256 93596
rect 97256 93540 97260 93596
rect 97196 93536 97260 93540
rect 97276 93596 97340 93600
rect 97276 93540 97280 93596
rect 97280 93540 97336 93596
rect 97336 93540 97340 93596
rect 97276 93536 97340 93540
rect 42012 93196 42076 93260
rect 4216 93052 4280 93056
rect 4216 92996 4220 93052
rect 4220 92996 4276 93052
rect 4276 92996 4280 93052
rect 4216 92992 4280 92996
rect 4296 93052 4360 93056
rect 4296 92996 4300 93052
rect 4300 92996 4356 93052
rect 4356 92996 4360 93052
rect 4296 92992 4360 92996
rect 4376 93052 4440 93056
rect 4376 92996 4380 93052
rect 4380 92996 4436 93052
rect 4436 92996 4440 93052
rect 4376 92992 4440 92996
rect 4456 93052 4520 93056
rect 4456 92996 4460 93052
rect 4460 92996 4516 93052
rect 4516 92996 4520 93052
rect 4456 92992 4520 92996
rect 34936 93052 35000 93056
rect 34936 92996 34940 93052
rect 34940 92996 34996 93052
rect 34996 92996 35000 93052
rect 34936 92992 35000 92996
rect 35016 93052 35080 93056
rect 35016 92996 35020 93052
rect 35020 92996 35076 93052
rect 35076 92996 35080 93052
rect 35016 92992 35080 92996
rect 35096 93052 35160 93056
rect 35096 92996 35100 93052
rect 35100 92996 35156 93052
rect 35156 92996 35160 93052
rect 35096 92992 35160 92996
rect 35176 93052 35240 93056
rect 35176 92996 35180 93052
rect 35180 92996 35236 93052
rect 35236 92996 35240 93052
rect 35176 92992 35240 92996
rect 65656 93052 65720 93056
rect 65656 92996 65660 93052
rect 65660 92996 65716 93052
rect 65716 92996 65720 93052
rect 65656 92992 65720 92996
rect 65736 93052 65800 93056
rect 65736 92996 65740 93052
rect 65740 92996 65796 93052
rect 65796 92996 65800 93052
rect 65736 92992 65800 92996
rect 65816 93052 65880 93056
rect 65816 92996 65820 93052
rect 65820 92996 65876 93052
rect 65876 92996 65880 93052
rect 65816 92992 65880 92996
rect 65896 93052 65960 93056
rect 65896 92996 65900 93052
rect 65900 92996 65956 93052
rect 65956 92996 65960 93052
rect 65896 92992 65960 92996
rect 96376 93052 96440 93056
rect 96376 92996 96380 93052
rect 96380 92996 96436 93052
rect 96436 92996 96440 93052
rect 96376 92992 96440 92996
rect 96456 93052 96520 93056
rect 96456 92996 96460 93052
rect 96460 92996 96516 93052
rect 96516 92996 96520 93052
rect 96456 92992 96520 92996
rect 96536 93052 96600 93056
rect 96536 92996 96540 93052
rect 96540 92996 96596 93052
rect 96596 92996 96600 93052
rect 96536 92992 96600 92996
rect 96616 93052 96680 93056
rect 96616 92996 96620 93052
rect 96620 92996 96676 93052
rect 96676 92996 96680 93052
rect 96616 92992 96680 92996
rect 56916 92924 56980 92988
rect 44588 92788 44652 92852
rect 51948 92788 52012 92852
rect 39620 92652 39684 92716
rect 38148 92516 38212 92580
rect 45876 92516 45940 92580
rect 61884 92652 61948 92716
rect 48268 92516 48332 92580
rect 64276 92516 64340 92580
rect 69244 92576 69308 92580
rect 69244 92520 69258 92576
rect 69258 92520 69308 92576
rect 69244 92516 69308 92520
rect 70716 92516 70780 92580
rect 4876 92508 4940 92512
rect 4876 92452 4880 92508
rect 4880 92452 4936 92508
rect 4936 92452 4940 92508
rect 4876 92448 4940 92452
rect 4956 92508 5020 92512
rect 4956 92452 4960 92508
rect 4960 92452 5016 92508
rect 5016 92452 5020 92508
rect 4956 92448 5020 92452
rect 5036 92508 5100 92512
rect 5036 92452 5040 92508
rect 5040 92452 5096 92508
rect 5096 92452 5100 92508
rect 5036 92448 5100 92452
rect 5116 92508 5180 92512
rect 5116 92452 5120 92508
rect 5120 92452 5176 92508
rect 5176 92452 5180 92508
rect 5116 92448 5180 92452
rect 35596 92508 35660 92512
rect 35596 92452 35600 92508
rect 35600 92452 35656 92508
rect 35656 92452 35660 92508
rect 35596 92448 35660 92452
rect 35676 92508 35740 92512
rect 35676 92452 35680 92508
rect 35680 92452 35736 92508
rect 35736 92452 35740 92508
rect 35676 92448 35740 92452
rect 35756 92508 35820 92512
rect 35756 92452 35760 92508
rect 35760 92452 35816 92508
rect 35816 92452 35820 92508
rect 35756 92448 35820 92452
rect 35836 92508 35900 92512
rect 35836 92452 35840 92508
rect 35840 92452 35896 92508
rect 35896 92452 35900 92508
rect 35836 92448 35900 92452
rect 66316 92508 66380 92512
rect 66316 92452 66320 92508
rect 66320 92452 66376 92508
rect 66376 92452 66380 92508
rect 66316 92448 66380 92452
rect 66396 92508 66460 92512
rect 66396 92452 66400 92508
rect 66400 92452 66456 92508
rect 66456 92452 66460 92508
rect 66396 92448 66460 92452
rect 66476 92508 66540 92512
rect 66476 92452 66480 92508
rect 66480 92452 66536 92508
rect 66536 92452 66540 92508
rect 66476 92448 66540 92452
rect 66556 92508 66620 92512
rect 66556 92452 66560 92508
rect 66560 92452 66616 92508
rect 66616 92452 66620 92508
rect 66556 92448 66620 92452
rect 97036 92508 97100 92512
rect 97036 92452 97040 92508
rect 97040 92452 97096 92508
rect 97096 92452 97100 92508
rect 97036 92448 97100 92452
rect 97116 92508 97180 92512
rect 97116 92452 97120 92508
rect 97120 92452 97176 92508
rect 97176 92452 97180 92508
rect 97116 92448 97180 92452
rect 97196 92508 97260 92512
rect 97196 92452 97200 92508
rect 97200 92452 97256 92508
rect 97256 92452 97260 92508
rect 97196 92448 97260 92452
rect 97276 92508 97340 92512
rect 97276 92452 97280 92508
rect 97280 92452 97336 92508
rect 97336 92452 97340 92508
rect 97276 92448 97340 92452
rect 113652 92508 113716 92512
rect 113652 92452 113656 92508
rect 113656 92452 113712 92508
rect 113712 92452 113716 92508
rect 113652 92448 113716 92452
rect 113732 92508 113796 92512
rect 113732 92452 113736 92508
rect 113736 92452 113792 92508
rect 113792 92452 113796 92508
rect 113732 92448 113796 92452
rect 113812 92508 113876 92512
rect 113812 92452 113816 92508
rect 113816 92452 113872 92508
rect 113872 92452 113876 92508
rect 113812 92448 113876 92452
rect 113892 92508 113956 92512
rect 113892 92452 113896 92508
rect 113896 92452 113952 92508
rect 113952 92452 113956 92508
rect 113892 92448 113956 92452
rect 43300 92108 43364 92172
rect 50660 92108 50724 92172
rect 53236 92108 53300 92172
rect 46796 91972 46860 92036
rect 4216 91964 4280 91968
rect 4216 91908 4220 91964
rect 4220 91908 4276 91964
rect 4276 91908 4280 91964
rect 4216 91904 4280 91908
rect 4296 91964 4360 91968
rect 4296 91908 4300 91964
rect 4300 91908 4356 91964
rect 4356 91908 4360 91964
rect 4296 91904 4360 91908
rect 4376 91964 4440 91968
rect 4376 91908 4380 91964
rect 4380 91908 4436 91964
rect 4436 91908 4440 91964
rect 4376 91904 4440 91908
rect 4456 91964 4520 91968
rect 4456 91908 4460 91964
rect 4460 91908 4516 91964
rect 4516 91908 4520 91964
rect 4456 91904 4520 91908
rect 34936 91964 35000 91968
rect 34936 91908 34940 91964
rect 34940 91908 34996 91964
rect 34996 91908 35000 91964
rect 34936 91904 35000 91908
rect 35016 91964 35080 91968
rect 35016 91908 35020 91964
rect 35020 91908 35076 91964
rect 35076 91908 35080 91964
rect 35016 91904 35080 91908
rect 35096 91964 35160 91968
rect 35096 91908 35100 91964
rect 35100 91908 35156 91964
rect 35156 91908 35160 91964
rect 35096 91904 35160 91908
rect 35176 91964 35240 91968
rect 35176 91908 35180 91964
rect 35180 91908 35236 91964
rect 35236 91908 35240 91964
rect 35176 91904 35240 91908
rect 65656 91964 65720 91968
rect 65656 91908 65660 91964
rect 65660 91908 65716 91964
rect 65716 91908 65720 91964
rect 65656 91904 65720 91908
rect 65736 91964 65800 91968
rect 65736 91908 65740 91964
rect 65740 91908 65796 91964
rect 65796 91908 65800 91964
rect 65736 91904 65800 91908
rect 65816 91964 65880 91968
rect 65816 91908 65820 91964
rect 65820 91908 65876 91964
rect 65876 91908 65880 91964
rect 65816 91904 65880 91908
rect 65896 91964 65960 91968
rect 65896 91908 65900 91964
rect 65900 91908 65956 91964
rect 65956 91908 65960 91964
rect 65896 91904 65960 91908
rect 96376 91964 96440 91968
rect 96376 91908 96380 91964
rect 96380 91908 96436 91964
rect 96436 91908 96440 91964
rect 96376 91904 96440 91908
rect 96456 91964 96520 91968
rect 96456 91908 96460 91964
rect 96460 91908 96516 91964
rect 96516 91908 96520 91964
rect 96456 91904 96520 91908
rect 96536 91964 96600 91968
rect 96536 91908 96540 91964
rect 96540 91908 96596 91964
rect 96596 91908 96600 91964
rect 96536 91904 96600 91908
rect 96616 91964 96680 91968
rect 96616 91908 96620 91964
rect 96620 91908 96676 91964
rect 96676 91908 96680 91964
rect 96616 91904 96680 91908
rect 112916 91964 112980 91968
rect 112916 91908 112920 91964
rect 112920 91908 112976 91964
rect 112976 91908 112980 91964
rect 112916 91904 112980 91908
rect 112996 91964 113060 91968
rect 112996 91908 113000 91964
rect 113000 91908 113056 91964
rect 113056 91908 113060 91964
rect 112996 91904 113060 91908
rect 113076 91964 113140 91968
rect 113076 91908 113080 91964
rect 113080 91908 113136 91964
rect 113136 91908 113140 91964
rect 113076 91904 113140 91908
rect 113156 91964 113220 91968
rect 113156 91908 113160 91964
rect 113160 91908 113216 91964
rect 113216 91908 113220 91964
rect 113156 91904 113220 91908
rect 4876 91420 4940 91424
rect 4876 91364 4880 91420
rect 4880 91364 4936 91420
rect 4936 91364 4940 91420
rect 4876 91360 4940 91364
rect 4956 91420 5020 91424
rect 4956 91364 4960 91420
rect 4960 91364 5016 91420
rect 5016 91364 5020 91420
rect 4956 91360 5020 91364
rect 5036 91420 5100 91424
rect 5036 91364 5040 91420
rect 5040 91364 5096 91420
rect 5096 91364 5100 91420
rect 5036 91360 5100 91364
rect 5116 91420 5180 91424
rect 5116 91364 5120 91420
rect 5120 91364 5176 91420
rect 5176 91364 5180 91420
rect 5116 91360 5180 91364
rect 113652 91420 113716 91424
rect 113652 91364 113656 91420
rect 113656 91364 113712 91420
rect 113712 91364 113716 91420
rect 113652 91360 113716 91364
rect 113732 91420 113796 91424
rect 113732 91364 113736 91420
rect 113736 91364 113792 91420
rect 113792 91364 113796 91420
rect 113732 91360 113796 91364
rect 113812 91420 113876 91424
rect 113812 91364 113816 91420
rect 113816 91364 113872 91420
rect 113872 91364 113876 91420
rect 113812 91360 113876 91364
rect 113892 91420 113956 91424
rect 113892 91364 113896 91420
rect 113896 91364 113952 91420
rect 113952 91364 113956 91420
rect 113892 91360 113956 91364
rect 99972 91216 100036 91220
rect 99972 91160 100022 91216
rect 100022 91160 100036 91216
rect 99972 91156 100036 91160
rect 62988 91020 63052 91084
rect 73292 91080 73356 91084
rect 73292 91024 73306 91080
rect 73306 91024 73356 91080
rect 73292 91020 73356 91024
rect 74212 91080 74276 91084
rect 74212 91024 74226 91080
rect 74226 91024 74276 91080
rect 74212 91020 74276 91024
rect 4216 90876 4280 90880
rect 4216 90820 4220 90876
rect 4220 90820 4276 90876
rect 4276 90820 4280 90876
rect 4216 90816 4280 90820
rect 4296 90876 4360 90880
rect 4296 90820 4300 90876
rect 4300 90820 4356 90876
rect 4356 90820 4360 90876
rect 4296 90816 4360 90820
rect 4376 90876 4440 90880
rect 4376 90820 4380 90876
rect 4380 90820 4436 90876
rect 4436 90820 4440 90876
rect 4376 90816 4440 90820
rect 4456 90876 4520 90880
rect 4456 90820 4460 90876
rect 4460 90820 4516 90876
rect 4516 90820 4520 90876
rect 4456 90816 4520 90820
rect 112916 90876 112980 90880
rect 112916 90820 112920 90876
rect 112920 90820 112976 90876
rect 112976 90820 112980 90876
rect 112916 90816 112980 90820
rect 112996 90876 113060 90880
rect 112996 90820 113000 90876
rect 113000 90820 113056 90876
rect 113056 90820 113060 90876
rect 112996 90816 113060 90820
rect 113076 90876 113140 90880
rect 113076 90820 113080 90876
rect 113080 90820 113136 90876
rect 113136 90820 113140 90876
rect 113076 90816 113140 90820
rect 113156 90876 113220 90880
rect 113156 90820 113160 90876
rect 113160 90820 113216 90876
rect 113216 90820 113220 90876
rect 113156 90816 113220 90820
rect 4876 90332 4940 90336
rect 4876 90276 4880 90332
rect 4880 90276 4936 90332
rect 4936 90276 4940 90332
rect 4876 90272 4940 90276
rect 4956 90332 5020 90336
rect 4956 90276 4960 90332
rect 4960 90276 5016 90332
rect 5016 90276 5020 90332
rect 4956 90272 5020 90276
rect 5036 90332 5100 90336
rect 5036 90276 5040 90332
rect 5040 90276 5096 90332
rect 5096 90276 5100 90332
rect 5036 90272 5100 90276
rect 5116 90332 5180 90336
rect 5116 90276 5120 90332
rect 5120 90276 5176 90332
rect 5176 90276 5180 90332
rect 5116 90272 5180 90276
rect 113652 90332 113716 90336
rect 113652 90276 113656 90332
rect 113656 90276 113712 90332
rect 113712 90276 113716 90332
rect 113652 90272 113716 90276
rect 113732 90332 113796 90336
rect 113732 90276 113736 90332
rect 113736 90276 113792 90332
rect 113792 90276 113796 90332
rect 113732 90272 113796 90276
rect 113812 90332 113876 90336
rect 113812 90276 113816 90332
rect 113816 90276 113872 90332
rect 113872 90276 113876 90332
rect 113812 90272 113876 90276
rect 113892 90332 113956 90336
rect 113892 90276 113896 90332
rect 113896 90276 113952 90332
rect 113952 90276 113956 90332
rect 113892 90272 113956 90276
rect 58150 89992 58214 89996
rect 58150 89936 58162 89992
rect 58162 89936 58214 89992
rect 58150 89932 58214 89936
rect 59510 89932 59574 89996
rect 55566 89796 55630 89860
rect 4216 89788 4280 89792
rect 4216 89732 4220 89788
rect 4220 89732 4276 89788
rect 4276 89732 4280 89788
rect 4216 89728 4280 89732
rect 4296 89788 4360 89792
rect 4296 89732 4300 89788
rect 4300 89732 4356 89788
rect 4356 89732 4360 89788
rect 4296 89728 4360 89732
rect 4376 89788 4440 89792
rect 4376 89732 4380 89788
rect 4380 89732 4436 89788
rect 4436 89732 4440 89788
rect 4376 89728 4440 89732
rect 4456 89788 4520 89792
rect 4456 89732 4460 89788
rect 4460 89732 4516 89788
rect 4516 89732 4520 89788
rect 4456 89728 4520 89732
rect 112916 89788 112980 89792
rect 112916 89732 112920 89788
rect 112920 89732 112976 89788
rect 112976 89732 112980 89788
rect 112916 89728 112980 89732
rect 112996 89788 113060 89792
rect 112996 89732 113000 89788
rect 113000 89732 113056 89788
rect 113056 89732 113060 89788
rect 112996 89728 113060 89732
rect 113076 89788 113140 89792
rect 113076 89732 113080 89788
rect 113080 89732 113136 89788
rect 113136 89732 113140 89788
rect 113076 89728 113140 89732
rect 113156 89788 113220 89792
rect 113156 89732 113160 89788
rect 113160 89732 113216 89788
rect 113216 89732 113220 89788
rect 113156 89728 113220 89732
rect 40606 89660 40670 89724
rect 54342 89660 54406 89724
rect 60598 89660 60662 89724
rect 65630 89660 65694 89724
rect 66854 89720 66918 89724
rect 66854 89664 66866 89720
rect 66866 89664 66918 89720
rect 66854 89660 66918 89664
rect 68214 89660 68278 89724
rect 71886 89720 71950 89724
rect 71886 89664 71926 89720
rect 71926 89664 71950 89720
rect 71886 89660 71950 89664
rect 75558 89660 75622 89724
rect 76918 89660 76982 89724
rect 89430 89720 89494 89724
rect 89430 89664 89442 89720
rect 89442 89664 89494 89720
rect 89430 89660 89494 89664
rect 4876 89244 4940 89248
rect 4876 89188 4880 89244
rect 4880 89188 4936 89244
rect 4936 89188 4940 89244
rect 4876 89184 4940 89188
rect 4956 89244 5020 89248
rect 4956 89188 4960 89244
rect 4960 89188 5016 89244
rect 5016 89188 5020 89244
rect 4956 89184 5020 89188
rect 5036 89244 5100 89248
rect 5036 89188 5040 89244
rect 5040 89188 5096 89244
rect 5096 89188 5100 89244
rect 5036 89184 5100 89188
rect 5116 89244 5180 89248
rect 5116 89188 5120 89244
rect 5120 89188 5176 89244
rect 5176 89188 5180 89244
rect 5116 89184 5180 89188
rect 113652 89244 113716 89248
rect 113652 89188 113656 89244
rect 113656 89188 113712 89244
rect 113712 89188 113716 89244
rect 113652 89184 113716 89188
rect 113732 89244 113796 89248
rect 113732 89188 113736 89244
rect 113736 89188 113792 89244
rect 113792 89188 113796 89244
rect 113732 89184 113796 89188
rect 113812 89244 113876 89248
rect 113812 89188 113816 89244
rect 113816 89188 113872 89244
rect 113872 89188 113876 89244
rect 113812 89184 113876 89188
rect 113892 89244 113956 89248
rect 113892 89188 113896 89244
rect 113896 89188 113952 89244
rect 113952 89188 113956 89244
rect 113892 89184 113956 89188
rect 4216 88700 4280 88704
rect 4216 88644 4220 88700
rect 4220 88644 4276 88700
rect 4276 88644 4280 88700
rect 4216 88640 4280 88644
rect 4296 88700 4360 88704
rect 4296 88644 4300 88700
rect 4300 88644 4356 88700
rect 4356 88644 4360 88700
rect 4296 88640 4360 88644
rect 4376 88700 4440 88704
rect 4376 88644 4380 88700
rect 4380 88644 4436 88700
rect 4436 88644 4440 88700
rect 4376 88640 4440 88644
rect 4456 88700 4520 88704
rect 4456 88644 4460 88700
rect 4460 88644 4516 88700
rect 4516 88644 4520 88700
rect 4456 88640 4520 88644
rect 112916 88700 112980 88704
rect 112916 88644 112920 88700
rect 112920 88644 112976 88700
rect 112976 88644 112980 88700
rect 112916 88640 112980 88644
rect 112996 88700 113060 88704
rect 112996 88644 113000 88700
rect 113000 88644 113056 88700
rect 113056 88644 113060 88700
rect 112996 88640 113060 88644
rect 113076 88700 113140 88704
rect 113076 88644 113080 88700
rect 113080 88644 113136 88700
rect 113136 88644 113140 88700
rect 113076 88640 113140 88644
rect 113156 88700 113220 88704
rect 113156 88644 113160 88700
rect 113160 88644 113216 88700
rect 113216 88644 113220 88700
rect 113156 88640 113220 88644
rect 4876 88156 4940 88160
rect 4876 88100 4880 88156
rect 4880 88100 4936 88156
rect 4936 88100 4940 88156
rect 4876 88096 4940 88100
rect 4956 88156 5020 88160
rect 4956 88100 4960 88156
rect 4960 88100 5016 88156
rect 5016 88100 5020 88156
rect 4956 88096 5020 88100
rect 5036 88156 5100 88160
rect 5036 88100 5040 88156
rect 5040 88100 5096 88156
rect 5096 88100 5100 88156
rect 5036 88096 5100 88100
rect 5116 88156 5180 88160
rect 5116 88100 5120 88156
rect 5120 88100 5176 88156
rect 5176 88100 5180 88156
rect 5116 88096 5180 88100
rect 113652 88156 113716 88160
rect 113652 88100 113656 88156
rect 113656 88100 113712 88156
rect 113712 88100 113716 88156
rect 113652 88096 113716 88100
rect 113732 88156 113796 88160
rect 113732 88100 113736 88156
rect 113736 88100 113792 88156
rect 113792 88100 113796 88156
rect 113732 88096 113796 88100
rect 113812 88156 113876 88160
rect 113812 88100 113816 88156
rect 113816 88100 113872 88156
rect 113872 88100 113876 88156
rect 113812 88096 113876 88100
rect 113892 88156 113956 88160
rect 113892 88100 113896 88156
rect 113896 88100 113952 88156
rect 113952 88100 113956 88156
rect 113892 88096 113956 88100
rect 4216 87612 4280 87616
rect 4216 87556 4220 87612
rect 4220 87556 4276 87612
rect 4276 87556 4280 87612
rect 4216 87552 4280 87556
rect 4296 87612 4360 87616
rect 4296 87556 4300 87612
rect 4300 87556 4356 87612
rect 4356 87556 4360 87612
rect 4296 87552 4360 87556
rect 4376 87612 4440 87616
rect 4376 87556 4380 87612
rect 4380 87556 4436 87612
rect 4436 87556 4440 87612
rect 4376 87552 4440 87556
rect 4456 87612 4520 87616
rect 4456 87556 4460 87612
rect 4460 87556 4516 87612
rect 4516 87556 4520 87612
rect 4456 87552 4520 87556
rect 112916 87612 112980 87616
rect 112916 87556 112920 87612
rect 112920 87556 112976 87612
rect 112976 87556 112980 87612
rect 112916 87552 112980 87556
rect 112996 87612 113060 87616
rect 112996 87556 113000 87612
rect 113000 87556 113056 87612
rect 113056 87556 113060 87612
rect 112996 87552 113060 87556
rect 113076 87612 113140 87616
rect 113076 87556 113080 87612
rect 113080 87556 113136 87612
rect 113136 87556 113140 87612
rect 113076 87552 113140 87556
rect 113156 87612 113220 87616
rect 113156 87556 113160 87612
rect 113160 87556 113216 87612
rect 113216 87556 113220 87612
rect 113156 87552 113220 87556
rect 4876 87068 4940 87072
rect 4876 87012 4880 87068
rect 4880 87012 4936 87068
rect 4936 87012 4940 87068
rect 4876 87008 4940 87012
rect 4956 87068 5020 87072
rect 4956 87012 4960 87068
rect 4960 87012 5016 87068
rect 5016 87012 5020 87068
rect 4956 87008 5020 87012
rect 5036 87068 5100 87072
rect 5036 87012 5040 87068
rect 5040 87012 5096 87068
rect 5096 87012 5100 87068
rect 5036 87008 5100 87012
rect 5116 87068 5180 87072
rect 5116 87012 5120 87068
rect 5120 87012 5176 87068
rect 5176 87012 5180 87068
rect 5116 87008 5180 87012
rect 113652 87068 113716 87072
rect 113652 87012 113656 87068
rect 113656 87012 113712 87068
rect 113712 87012 113716 87068
rect 113652 87008 113716 87012
rect 113732 87068 113796 87072
rect 113732 87012 113736 87068
rect 113736 87012 113792 87068
rect 113792 87012 113796 87068
rect 113732 87008 113796 87012
rect 113812 87068 113876 87072
rect 113812 87012 113816 87068
rect 113816 87012 113872 87068
rect 113872 87012 113876 87068
rect 113812 87008 113876 87012
rect 113892 87068 113956 87072
rect 113892 87012 113896 87068
rect 113896 87012 113952 87068
rect 113952 87012 113956 87068
rect 113892 87008 113956 87012
rect 4216 86524 4280 86528
rect 4216 86468 4220 86524
rect 4220 86468 4276 86524
rect 4276 86468 4280 86524
rect 4216 86464 4280 86468
rect 4296 86524 4360 86528
rect 4296 86468 4300 86524
rect 4300 86468 4356 86524
rect 4356 86468 4360 86524
rect 4296 86464 4360 86468
rect 4376 86524 4440 86528
rect 4376 86468 4380 86524
rect 4380 86468 4436 86524
rect 4436 86468 4440 86524
rect 4376 86464 4440 86468
rect 4456 86524 4520 86528
rect 4456 86468 4460 86524
rect 4460 86468 4516 86524
rect 4516 86468 4520 86524
rect 4456 86464 4520 86468
rect 112916 86524 112980 86528
rect 112916 86468 112920 86524
rect 112920 86468 112976 86524
rect 112976 86468 112980 86524
rect 112916 86464 112980 86468
rect 112996 86524 113060 86528
rect 112996 86468 113000 86524
rect 113000 86468 113056 86524
rect 113056 86468 113060 86524
rect 112996 86464 113060 86468
rect 113076 86524 113140 86528
rect 113076 86468 113080 86524
rect 113080 86468 113136 86524
rect 113136 86468 113140 86524
rect 113076 86464 113140 86468
rect 113156 86524 113220 86528
rect 113156 86468 113160 86524
rect 113160 86468 113216 86524
rect 113216 86468 113220 86524
rect 113156 86464 113220 86468
rect 4876 85980 4940 85984
rect 4876 85924 4880 85980
rect 4880 85924 4936 85980
rect 4936 85924 4940 85980
rect 4876 85920 4940 85924
rect 4956 85980 5020 85984
rect 4956 85924 4960 85980
rect 4960 85924 5016 85980
rect 5016 85924 5020 85980
rect 4956 85920 5020 85924
rect 5036 85980 5100 85984
rect 5036 85924 5040 85980
rect 5040 85924 5096 85980
rect 5096 85924 5100 85980
rect 5036 85920 5100 85924
rect 5116 85980 5180 85984
rect 5116 85924 5120 85980
rect 5120 85924 5176 85980
rect 5176 85924 5180 85980
rect 5116 85920 5180 85924
rect 113652 85980 113716 85984
rect 113652 85924 113656 85980
rect 113656 85924 113712 85980
rect 113712 85924 113716 85980
rect 113652 85920 113716 85924
rect 113732 85980 113796 85984
rect 113732 85924 113736 85980
rect 113736 85924 113792 85980
rect 113792 85924 113796 85980
rect 113732 85920 113796 85924
rect 113812 85980 113876 85984
rect 113812 85924 113816 85980
rect 113816 85924 113872 85980
rect 113872 85924 113876 85980
rect 113812 85920 113876 85924
rect 113892 85980 113956 85984
rect 113892 85924 113896 85980
rect 113896 85924 113952 85980
rect 113952 85924 113956 85980
rect 113892 85920 113956 85924
rect 4216 85436 4280 85440
rect 4216 85380 4220 85436
rect 4220 85380 4276 85436
rect 4276 85380 4280 85436
rect 4216 85376 4280 85380
rect 4296 85436 4360 85440
rect 4296 85380 4300 85436
rect 4300 85380 4356 85436
rect 4356 85380 4360 85436
rect 4296 85376 4360 85380
rect 4376 85436 4440 85440
rect 4376 85380 4380 85436
rect 4380 85380 4436 85436
rect 4436 85380 4440 85436
rect 4376 85376 4440 85380
rect 4456 85436 4520 85440
rect 4456 85380 4460 85436
rect 4460 85380 4516 85436
rect 4516 85380 4520 85436
rect 4456 85376 4520 85380
rect 112916 85436 112980 85440
rect 112916 85380 112920 85436
rect 112920 85380 112976 85436
rect 112976 85380 112980 85436
rect 112916 85376 112980 85380
rect 112996 85436 113060 85440
rect 112996 85380 113000 85436
rect 113000 85380 113056 85436
rect 113056 85380 113060 85436
rect 112996 85376 113060 85380
rect 113076 85436 113140 85440
rect 113076 85380 113080 85436
rect 113080 85380 113136 85436
rect 113136 85380 113140 85436
rect 113076 85376 113140 85380
rect 113156 85436 113220 85440
rect 113156 85380 113160 85436
rect 113160 85380 113216 85436
rect 113216 85380 113220 85436
rect 113156 85376 113220 85380
rect 4876 84892 4940 84896
rect 4876 84836 4880 84892
rect 4880 84836 4936 84892
rect 4936 84836 4940 84892
rect 4876 84832 4940 84836
rect 4956 84892 5020 84896
rect 4956 84836 4960 84892
rect 4960 84836 5016 84892
rect 5016 84836 5020 84892
rect 4956 84832 5020 84836
rect 5036 84892 5100 84896
rect 5036 84836 5040 84892
rect 5040 84836 5096 84892
rect 5096 84836 5100 84892
rect 5036 84832 5100 84836
rect 5116 84892 5180 84896
rect 5116 84836 5120 84892
rect 5120 84836 5176 84892
rect 5176 84836 5180 84892
rect 5116 84832 5180 84836
rect 113652 84892 113716 84896
rect 113652 84836 113656 84892
rect 113656 84836 113712 84892
rect 113712 84836 113716 84892
rect 113652 84832 113716 84836
rect 113732 84892 113796 84896
rect 113732 84836 113736 84892
rect 113736 84836 113792 84892
rect 113792 84836 113796 84892
rect 113732 84832 113796 84836
rect 113812 84892 113876 84896
rect 113812 84836 113816 84892
rect 113816 84836 113872 84892
rect 113872 84836 113876 84892
rect 113812 84832 113876 84836
rect 113892 84892 113956 84896
rect 113892 84836 113896 84892
rect 113896 84836 113952 84892
rect 113952 84836 113956 84892
rect 113892 84832 113956 84836
rect 4216 84348 4280 84352
rect 4216 84292 4220 84348
rect 4220 84292 4276 84348
rect 4276 84292 4280 84348
rect 4216 84288 4280 84292
rect 4296 84348 4360 84352
rect 4296 84292 4300 84348
rect 4300 84292 4356 84348
rect 4356 84292 4360 84348
rect 4296 84288 4360 84292
rect 4376 84348 4440 84352
rect 4376 84292 4380 84348
rect 4380 84292 4436 84348
rect 4436 84292 4440 84348
rect 4376 84288 4440 84292
rect 4456 84348 4520 84352
rect 4456 84292 4460 84348
rect 4460 84292 4516 84348
rect 4516 84292 4520 84348
rect 4456 84288 4520 84292
rect 112916 84348 112980 84352
rect 112916 84292 112920 84348
rect 112920 84292 112976 84348
rect 112976 84292 112980 84348
rect 112916 84288 112980 84292
rect 112996 84348 113060 84352
rect 112996 84292 113000 84348
rect 113000 84292 113056 84348
rect 113056 84292 113060 84348
rect 112996 84288 113060 84292
rect 113076 84348 113140 84352
rect 113076 84292 113080 84348
rect 113080 84292 113136 84348
rect 113136 84292 113140 84348
rect 113076 84288 113140 84292
rect 113156 84348 113220 84352
rect 113156 84292 113160 84348
rect 113160 84292 113216 84348
rect 113216 84292 113220 84348
rect 113156 84288 113220 84292
rect 4876 83804 4940 83808
rect 4876 83748 4880 83804
rect 4880 83748 4936 83804
rect 4936 83748 4940 83804
rect 4876 83744 4940 83748
rect 4956 83804 5020 83808
rect 4956 83748 4960 83804
rect 4960 83748 5016 83804
rect 5016 83748 5020 83804
rect 4956 83744 5020 83748
rect 5036 83804 5100 83808
rect 5036 83748 5040 83804
rect 5040 83748 5096 83804
rect 5096 83748 5100 83804
rect 5036 83744 5100 83748
rect 5116 83804 5180 83808
rect 5116 83748 5120 83804
rect 5120 83748 5176 83804
rect 5176 83748 5180 83804
rect 5116 83744 5180 83748
rect 113652 83804 113716 83808
rect 113652 83748 113656 83804
rect 113656 83748 113712 83804
rect 113712 83748 113716 83804
rect 113652 83744 113716 83748
rect 113732 83804 113796 83808
rect 113732 83748 113736 83804
rect 113736 83748 113792 83804
rect 113792 83748 113796 83804
rect 113732 83744 113796 83748
rect 113812 83804 113876 83808
rect 113812 83748 113816 83804
rect 113816 83748 113872 83804
rect 113872 83748 113876 83804
rect 113812 83744 113876 83748
rect 113892 83804 113956 83808
rect 113892 83748 113896 83804
rect 113896 83748 113952 83804
rect 113952 83748 113956 83804
rect 113892 83744 113956 83748
rect 4216 83260 4280 83264
rect 4216 83204 4220 83260
rect 4220 83204 4276 83260
rect 4276 83204 4280 83260
rect 4216 83200 4280 83204
rect 4296 83260 4360 83264
rect 4296 83204 4300 83260
rect 4300 83204 4356 83260
rect 4356 83204 4360 83260
rect 4296 83200 4360 83204
rect 4376 83260 4440 83264
rect 4376 83204 4380 83260
rect 4380 83204 4436 83260
rect 4436 83204 4440 83260
rect 4376 83200 4440 83204
rect 4456 83260 4520 83264
rect 4456 83204 4460 83260
rect 4460 83204 4516 83260
rect 4516 83204 4520 83260
rect 4456 83200 4520 83204
rect 112916 83260 112980 83264
rect 112916 83204 112920 83260
rect 112920 83204 112976 83260
rect 112976 83204 112980 83260
rect 112916 83200 112980 83204
rect 112996 83260 113060 83264
rect 112996 83204 113000 83260
rect 113000 83204 113056 83260
rect 113056 83204 113060 83260
rect 112996 83200 113060 83204
rect 113076 83260 113140 83264
rect 113076 83204 113080 83260
rect 113080 83204 113136 83260
rect 113136 83204 113140 83260
rect 113076 83200 113140 83204
rect 113156 83260 113220 83264
rect 113156 83204 113160 83260
rect 113160 83204 113216 83260
rect 113216 83204 113220 83260
rect 113156 83200 113220 83204
rect 4876 82716 4940 82720
rect 4876 82660 4880 82716
rect 4880 82660 4936 82716
rect 4936 82660 4940 82716
rect 4876 82656 4940 82660
rect 4956 82716 5020 82720
rect 4956 82660 4960 82716
rect 4960 82660 5016 82716
rect 5016 82660 5020 82716
rect 4956 82656 5020 82660
rect 5036 82716 5100 82720
rect 5036 82660 5040 82716
rect 5040 82660 5096 82716
rect 5096 82660 5100 82716
rect 5036 82656 5100 82660
rect 5116 82716 5180 82720
rect 5116 82660 5120 82716
rect 5120 82660 5176 82716
rect 5176 82660 5180 82716
rect 5116 82656 5180 82660
rect 113652 82716 113716 82720
rect 113652 82660 113656 82716
rect 113656 82660 113712 82716
rect 113712 82660 113716 82716
rect 113652 82656 113716 82660
rect 113732 82716 113796 82720
rect 113732 82660 113736 82716
rect 113736 82660 113792 82716
rect 113792 82660 113796 82716
rect 113732 82656 113796 82660
rect 113812 82716 113876 82720
rect 113812 82660 113816 82716
rect 113816 82660 113872 82716
rect 113872 82660 113876 82716
rect 113812 82656 113876 82660
rect 113892 82716 113956 82720
rect 113892 82660 113896 82716
rect 113896 82660 113952 82716
rect 113952 82660 113956 82716
rect 113892 82656 113956 82660
rect 4216 82172 4280 82176
rect 4216 82116 4220 82172
rect 4220 82116 4276 82172
rect 4276 82116 4280 82172
rect 4216 82112 4280 82116
rect 4296 82172 4360 82176
rect 4296 82116 4300 82172
rect 4300 82116 4356 82172
rect 4356 82116 4360 82172
rect 4296 82112 4360 82116
rect 4376 82172 4440 82176
rect 4376 82116 4380 82172
rect 4380 82116 4436 82172
rect 4436 82116 4440 82172
rect 4376 82112 4440 82116
rect 4456 82172 4520 82176
rect 4456 82116 4460 82172
rect 4460 82116 4516 82172
rect 4516 82116 4520 82172
rect 4456 82112 4520 82116
rect 112916 82172 112980 82176
rect 112916 82116 112920 82172
rect 112920 82116 112976 82172
rect 112976 82116 112980 82172
rect 112916 82112 112980 82116
rect 112996 82172 113060 82176
rect 112996 82116 113000 82172
rect 113000 82116 113056 82172
rect 113056 82116 113060 82172
rect 112996 82112 113060 82116
rect 113076 82172 113140 82176
rect 113076 82116 113080 82172
rect 113080 82116 113136 82172
rect 113136 82116 113140 82172
rect 113076 82112 113140 82116
rect 113156 82172 113220 82176
rect 113156 82116 113160 82172
rect 113160 82116 113216 82172
rect 113216 82116 113220 82172
rect 113156 82112 113220 82116
rect 4876 81628 4940 81632
rect 4876 81572 4880 81628
rect 4880 81572 4936 81628
rect 4936 81572 4940 81628
rect 4876 81568 4940 81572
rect 4956 81628 5020 81632
rect 4956 81572 4960 81628
rect 4960 81572 5016 81628
rect 5016 81572 5020 81628
rect 4956 81568 5020 81572
rect 5036 81628 5100 81632
rect 5036 81572 5040 81628
rect 5040 81572 5096 81628
rect 5096 81572 5100 81628
rect 5036 81568 5100 81572
rect 5116 81628 5180 81632
rect 5116 81572 5120 81628
rect 5120 81572 5176 81628
rect 5176 81572 5180 81628
rect 5116 81568 5180 81572
rect 113652 81628 113716 81632
rect 113652 81572 113656 81628
rect 113656 81572 113712 81628
rect 113712 81572 113716 81628
rect 113652 81568 113716 81572
rect 113732 81628 113796 81632
rect 113732 81572 113736 81628
rect 113736 81572 113792 81628
rect 113792 81572 113796 81628
rect 113732 81568 113796 81572
rect 113812 81628 113876 81632
rect 113812 81572 113816 81628
rect 113816 81572 113872 81628
rect 113872 81572 113876 81628
rect 113812 81568 113876 81572
rect 113892 81628 113956 81632
rect 113892 81572 113896 81628
rect 113896 81572 113952 81628
rect 113952 81572 113956 81628
rect 113892 81568 113956 81572
rect 4216 81084 4280 81088
rect 4216 81028 4220 81084
rect 4220 81028 4276 81084
rect 4276 81028 4280 81084
rect 4216 81024 4280 81028
rect 4296 81084 4360 81088
rect 4296 81028 4300 81084
rect 4300 81028 4356 81084
rect 4356 81028 4360 81084
rect 4296 81024 4360 81028
rect 4376 81084 4440 81088
rect 4376 81028 4380 81084
rect 4380 81028 4436 81084
rect 4436 81028 4440 81084
rect 4376 81024 4440 81028
rect 4456 81084 4520 81088
rect 4456 81028 4460 81084
rect 4460 81028 4516 81084
rect 4516 81028 4520 81084
rect 4456 81024 4520 81028
rect 112916 81084 112980 81088
rect 112916 81028 112920 81084
rect 112920 81028 112976 81084
rect 112976 81028 112980 81084
rect 112916 81024 112980 81028
rect 112996 81084 113060 81088
rect 112996 81028 113000 81084
rect 113000 81028 113056 81084
rect 113056 81028 113060 81084
rect 112996 81024 113060 81028
rect 113076 81084 113140 81088
rect 113076 81028 113080 81084
rect 113080 81028 113136 81084
rect 113136 81028 113140 81084
rect 113076 81024 113140 81028
rect 113156 81084 113220 81088
rect 113156 81028 113160 81084
rect 113160 81028 113216 81084
rect 113216 81028 113220 81084
rect 113156 81024 113220 81028
rect 4876 80540 4940 80544
rect 4876 80484 4880 80540
rect 4880 80484 4936 80540
rect 4936 80484 4940 80540
rect 4876 80480 4940 80484
rect 4956 80540 5020 80544
rect 4956 80484 4960 80540
rect 4960 80484 5016 80540
rect 5016 80484 5020 80540
rect 4956 80480 5020 80484
rect 5036 80540 5100 80544
rect 5036 80484 5040 80540
rect 5040 80484 5096 80540
rect 5096 80484 5100 80540
rect 5036 80480 5100 80484
rect 5116 80540 5180 80544
rect 5116 80484 5120 80540
rect 5120 80484 5176 80540
rect 5176 80484 5180 80540
rect 5116 80480 5180 80484
rect 113652 80540 113716 80544
rect 113652 80484 113656 80540
rect 113656 80484 113712 80540
rect 113712 80484 113716 80540
rect 113652 80480 113716 80484
rect 113732 80540 113796 80544
rect 113732 80484 113736 80540
rect 113736 80484 113792 80540
rect 113792 80484 113796 80540
rect 113732 80480 113796 80484
rect 113812 80540 113876 80544
rect 113812 80484 113816 80540
rect 113816 80484 113872 80540
rect 113872 80484 113876 80540
rect 113812 80480 113876 80484
rect 113892 80540 113956 80544
rect 113892 80484 113896 80540
rect 113896 80484 113952 80540
rect 113952 80484 113956 80540
rect 113892 80480 113956 80484
rect 4216 79996 4280 80000
rect 4216 79940 4220 79996
rect 4220 79940 4276 79996
rect 4276 79940 4280 79996
rect 4216 79936 4280 79940
rect 4296 79996 4360 80000
rect 4296 79940 4300 79996
rect 4300 79940 4356 79996
rect 4356 79940 4360 79996
rect 4296 79936 4360 79940
rect 4376 79996 4440 80000
rect 4376 79940 4380 79996
rect 4380 79940 4436 79996
rect 4436 79940 4440 79996
rect 4376 79936 4440 79940
rect 4456 79996 4520 80000
rect 4456 79940 4460 79996
rect 4460 79940 4516 79996
rect 4516 79940 4520 79996
rect 4456 79936 4520 79940
rect 112916 79996 112980 80000
rect 112916 79940 112920 79996
rect 112920 79940 112976 79996
rect 112976 79940 112980 79996
rect 112916 79936 112980 79940
rect 112996 79996 113060 80000
rect 112996 79940 113000 79996
rect 113000 79940 113056 79996
rect 113056 79940 113060 79996
rect 112996 79936 113060 79940
rect 113076 79996 113140 80000
rect 113076 79940 113080 79996
rect 113080 79940 113136 79996
rect 113136 79940 113140 79996
rect 113076 79936 113140 79940
rect 113156 79996 113220 80000
rect 113156 79940 113160 79996
rect 113160 79940 113216 79996
rect 113216 79940 113220 79996
rect 113156 79936 113220 79940
rect 4876 79452 4940 79456
rect 4876 79396 4880 79452
rect 4880 79396 4936 79452
rect 4936 79396 4940 79452
rect 4876 79392 4940 79396
rect 4956 79452 5020 79456
rect 4956 79396 4960 79452
rect 4960 79396 5016 79452
rect 5016 79396 5020 79452
rect 4956 79392 5020 79396
rect 5036 79452 5100 79456
rect 5036 79396 5040 79452
rect 5040 79396 5096 79452
rect 5096 79396 5100 79452
rect 5036 79392 5100 79396
rect 5116 79452 5180 79456
rect 5116 79396 5120 79452
rect 5120 79396 5176 79452
rect 5176 79396 5180 79452
rect 5116 79392 5180 79396
rect 113652 79452 113716 79456
rect 113652 79396 113656 79452
rect 113656 79396 113712 79452
rect 113712 79396 113716 79452
rect 113652 79392 113716 79396
rect 113732 79452 113796 79456
rect 113732 79396 113736 79452
rect 113736 79396 113792 79452
rect 113792 79396 113796 79452
rect 113732 79392 113796 79396
rect 113812 79452 113876 79456
rect 113812 79396 113816 79452
rect 113816 79396 113872 79452
rect 113872 79396 113876 79452
rect 113812 79392 113876 79396
rect 113892 79452 113956 79456
rect 113892 79396 113896 79452
rect 113896 79396 113952 79452
rect 113952 79396 113956 79452
rect 113892 79392 113956 79396
rect 4216 78908 4280 78912
rect 4216 78852 4220 78908
rect 4220 78852 4276 78908
rect 4276 78852 4280 78908
rect 4216 78848 4280 78852
rect 4296 78908 4360 78912
rect 4296 78852 4300 78908
rect 4300 78852 4356 78908
rect 4356 78852 4360 78908
rect 4296 78848 4360 78852
rect 4376 78908 4440 78912
rect 4376 78852 4380 78908
rect 4380 78852 4436 78908
rect 4436 78852 4440 78908
rect 4376 78848 4440 78852
rect 4456 78908 4520 78912
rect 4456 78852 4460 78908
rect 4460 78852 4516 78908
rect 4516 78852 4520 78908
rect 4456 78848 4520 78852
rect 112916 78908 112980 78912
rect 112916 78852 112920 78908
rect 112920 78852 112976 78908
rect 112976 78852 112980 78908
rect 112916 78848 112980 78852
rect 112996 78908 113060 78912
rect 112996 78852 113000 78908
rect 113000 78852 113056 78908
rect 113056 78852 113060 78908
rect 112996 78848 113060 78852
rect 113076 78908 113140 78912
rect 113076 78852 113080 78908
rect 113080 78852 113136 78908
rect 113136 78852 113140 78908
rect 113076 78848 113140 78852
rect 113156 78908 113220 78912
rect 113156 78852 113160 78908
rect 113160 78852 113216 78908
rect 113216 78852 113220 78908
rect 113156 78848 113220 78852
rect 4876 78364 4940 78368
rect 4876 78308 4880 78364
rect 4880 78308 4936 78364
rect 4936 78308 4940 78364
rect 4876 78304 4940 78308
rect 4956 78364 5020 78368
rect 4956 78308 4960 78364
rect 4960 78308 5016 78364
rect 5016 78308 5020 78364
rect 4956 78304 5020 78308
rect 5036 78364 5100 78368
rect 5036 78308 5040 78364
rect 5040 78308 5096 78364
rect 5096 78308 5100 78364
rect 5036 78304 5100 78308
rect 5116 78364 5180 78368
rect 5116 78308 5120 78364
rect 5120 78308 5176 78364
rect 5176 78308 5180 78364
rect 5116 78304 5180 78308
rect 113652 78364 113716 78368
rect 113652 78308 113656 78364
rect 113656 78308 113712 78364
rect 113712 78308 113716 78364
rect 113652 78304 113716 78308
rect 113732 78364 113796 78368
rect 113732 78308 113736 78364
rect 113736 78308 113792 78364
rect 113792 78308 113796 78364
rect 113732 78304 113796 78308
rect 113812 78364 113876 78368
rect 113812 78308 113816 78364
rect 113816 78308 113872 78364
rect 113872 78308 113876 78364
rect 113812 78304 113876 78308
rect 113892 78364 113956 78368
rect 113892 78308 113896 78364
rect 113896 78308 113952 78364
rect 113952 78308 113956 78364
rect 113892 78304 113956 78308
rect 4216 77820 4280 77824
rect 4216 77764 4220 77820
rect 4220 77764 4276 77820
rect 4276 77764 4280 77820
rect 4216 77760 4280 77764
rect 4296 77820 4360 77824
rect 4296 77764 4300 77820
rect 4300 77764 4356 77820
rect 4356 77764 4360 77820
rect 4296 77760 4360 77764
rect 4376 77820 4440 77824
rect 4376 77764 4380 77820
rect 4380 77764 4436 77820
rect 4436 77764 4440 77820
rect 4376 77760 4440 77764
rect 4456 77820 4520 77824
rect 4456 77764 4460 77820
rect 4460 77764 4516 77820
rect 4516 77764 4520 77820
rect 4456 77760 4520 77764
rect 112916 77820 112980 77824
rect 112916 77764 112920 77820
rect 112920 77764 112976 77820
rect 112976 77764 112980 77820
rect 112916 77760 112980 77764
rect 112996 77820 113060 77824
rect 112996 77764 113000 77820
rect 113000 77764 113056 77820
rect 113056 77764 113060 77820
rect 112996 77760 113060 77764
rect 113076 77820 113140 77824
rect 113076 77764 113080 77820
rect 113080 77764 113136 77820
rect 113136 77764 113140 77820
rect 113076 77760 113140 77764
rect 113156 77820 113220 77824
rect 113156 77764 113160 77820
rect 113160 77764 113216 77820
rect 113216 77764 113220 77820
rect 113156 77760 113220 77764
rect 4876 77276 4940 77280
rect 4876 77220 4880 77276
rect 4880 77220 4936 77276
rect 4936 77220 4940 77276
rect 4876 77216 4940 77220
rect 4956 77276 5020 77280
rect 4956 77220 4960 77276
rect 4960 77220 5016 77276
rect 5016 77220 5020 77276
rect 4956 77216 5020 77220
rect 5036 77276 5100 77280
rect 5036 77220 5040 77276
rect 5040 77220 5096 77276
rect 5096 77220 5100 77276
rect 5036 77216 5100 77220
rect 5116 77276 5180 77280
rect 5116 77220 5120 77276
rect 5120 77220 5176 77276
rect 5176 77220 5180 77276
rect 5116 77216 5180 77220
rect 113652 77276 113716 77280
rect 113652 77220 113656 77276
rect 113656 77220 113712 77276
rect 113712 77220 113716 77276
rect 113652 77216 113716 77220
rect 113732 77276 113796 77280
rect 113732 77220 113736 77276
rect 113736 77220 113792 77276
rect 113792 77220 113796 77276
rect 113732 77216 113796 77220
rect 113812 77276 113876 77280
rect 113812 77220 113816 77276
rect 113816 77220 113872 77276
rect 113872 77220 113876 77276
rect 113812 77216 113876 77220
rect 113892 77276 113956 77280
rect 113892 77220 113896 77276
rect 113896 77220 113952 77276
rect 113952 77220 113956 77276
rect 113892 77216 113956 77220
rect 4216 76732 4280 76736
rect 4216 76676 4220 76732
rect 4220 76676 4276 76732
rect 4276 76676 4280 76732
rect 4216 76672 4280 76676
rect 4296 76732 4360 76736
rect 4296 76676 4300 76732
rect 4300 76676 4356 76732
rect 4356 76676 4360 76732
rect 4296 76672 4360 76676
rect 4376 76732 4440 76736
rect 4376 76676 4380 76732
rect 4380 76676 4436 76732
rect 4436 76676 4440 76732
rect 4376 76672 4440 76676
rect 4456 76732 4520 76736
rect 4456 76676 4460 76732
rect 4460 76676 4516 76732
rect 4516 76676 4520 76732
rect 4456 76672 4520 76676
rect 112916 76732 112980 76736
rect 112916 76676 112920 76732
rect 112920 76676 112976 76732
rect 112976 76676 112980 76732
rect 112916 76672 112980 76676
rect 112996 76732 113060 76736
rect 112996 76676 113000 76732
rect 113000 76676 113056 76732
rect 113056 76676 113060 76732
rect 112996 76672 113060 76676
rect 113076 76732 113140 76736
rect 113076 76676 113080 76732
rect 113080 76676 113136 76732
rect 113136 76676 113140 76732
rect 113076 76672 113140 76676
rect 113156 76732 113220 76736
rect 113156 76676 113160 76732
rect 113160 76676 113216 76732
rect 113216 76676 113220 76732
rect 113156 76672 113220 76676
rect 4876 76188 4940 76192
rect 4876 76132 4880 76188
rect 4880 76132 4936 76188
rect 4936 76132 4940 76188
rect 4876 76128 4940 76132
rect 4956 76188 5020 76192
rect 4956 76132 4960 76188
rect 4960 76132 5016 76188
rect 5016 76132 5020 76188
rect 4956 76128 5020 76132
rect 5036 76188 5100 76192
rect 5036 76132 5040 76188
rect 5040 76132 5096 76188
rect 5096 76132 5100 76188
rect 5036 76128 5100 76132
rect 5116 76188 5180 76192
rect 5116 76132 5120 76188
rect 5120 76132 5176 76188
rect 5176 76132 5180 76188
rect 5116 76128 5180 76132
rect 113652 76188 113716 76192
rect 113652 76132 113656 76188
rect 113656 76132 113712 76188
rect 113712 76132 113716 76188
rect 113652 76128 113716 76132
rect 113732 76188 113796 76192
rect 113732 76132 113736 76188
rect 113736 76132 113792 76188
rect 113792 76132 113796 76188
rect 113732 76128 113796 76132
rect 113812 76188 113876 76192
rect 113812 76132 113816 76188
rect 113816 76132 113872 76188
rect 113872 76132 113876 76188
rect 113812 76128 113876 76132
rect 113892 76188 113956 76192
rect 113892 76132 113896 76188
rect 113896 76132 113952 76188
rect 113952 76132 113956 76188
rect 113892 76128 113956 76132
rect 4216 75644 4280 75648
rect 4216 75588 4220 75644
rect 4220 75588 4276 75644
rect 4276 75588 4280 75644
rect 4216 75584 4280 75588
rect 4296 75644 4360 75648
rect 4296 75588 4300 75644
rect 4300 75588 4356 75644
rect 4356 75588 4360 75644
rect 4296 75584 4360 75588
rect 4376 75644 4440 75648
rect 4376 75588 4380 75644
rect 4380 75588 4436 75644
rect 4436 75588 4440 75644
rect 4376 75584 4440 75588
rect 4456 75644 4520 75648
rect 4456 75588 4460 75644
rect 4460 75588 4516 75644
rect 4516 75588 4520 75644
rect 4456 75584 4520 75588
rect 112916 75644 112980 75648
rect 112916 75588 112920 75644
rect 112920 75588 112976 75644
rect 112976 75588 112980 75644
rect 112916 75584 112980 75588
rect 112996 75644 113060 75648
rect 112996 75588 113000 75644
rect 113000 75588 113056 75644
rect 113056 75588 113060 75644
rect 112996 75584 113060 75588
rect 113076 75644 113140 75648
rect 113076 75588 113080 75644
rect 113080 75588 113136 75644
rect 113136 75588 113140 75644
rect 113076 75584 113140 75588
rect 113156 75644 113220 75648
rect 113156 75588 113160 75644
rect 113160 75588 113216 75644
rect 113216 75588 113220 75644
rect 113156 75584 113220 75588
rect 4876 75100 4940 75104
rect 4876 75044 4880 75100
rect 4880 75044 4936 75100
rect 4936 75044 4940 75100
rect 4876 75040 4940 75044
rect 4956 75100 5020 75104
rect 4956 75044 4960 75100
rect 4960 75044 5016 75100
rect 5016 75044 5020 75100
rect 4956 75040 5020 75044
rect 5036 75100 5100 75104
rect 5036 75044 5040 75100
rect 5040 75044 5096 75100
rect 5096 75044 5100 75100
rect 5036 75040 5100 75044
rect 5116 75100 5180 75104
rect 5116 75044 5120 75100
rect 5120 75044 5176 75100
rect 5176 75044 5180 75100
rect 5116 75040 5180 75044
rect 113652 75100 113716 75104
rect 113652 75044 113656 75100
rect 113656 75044 113712 75100
rect 113712 75044 113716 75100
rect 113652 75040 113716 75044
rect 113732 75100 113796 75104
rect 113732 75044 113736 75100
rect 113736 75044 113792 75100
rect 113792 75044 113796 75100
rect 113732 75040 113796 75044
rect 113812 75100 113876 75104
rect 113812 75044 113816 75100
rect 113816 75044 113872 75100
rect 113872 75044 113876 75100
rect 113812 75040 113876 75044
rect 113892 75100 113956 75104
rect 113892 75044 113896 75100
rect 113896 75044 113952 75100
rect 113952 75044 113956 75100
rect 113892 75040 113956 75044
rect 4216 74556 4280 74560
rect 4216 74500 4220 74556
rect 4220 74500 4276 74556
rect 4276 74500 4280 74556
rect 4216 74496 4280 74500
rect 4296 74556 4360 74560
rect 4296 74500 4300 74556
rect 4300 74500 4356 74556
rect 4356 74500 4360 74556
rect 4296 74496 4360 74500
rect 4376 74556 4440 74560
rect 4376 74500 4380 74556
rect 4380 74500 4436 74556
rect 4436 74500 4440 74556
rect 4376 74496 4440 74500
rect 4456 74556 4520 74560
rect 4456 74500 4460 74556
rect 4460 74500 4516 74556
rect 4516 74500 4520 74556
rect 4456 74496 4520 74500
rect 112916 74556 112980 74560
rect 112916 74500 112920 74556
rect 112920 74500 112976 74556
rect 112976 74500 112980 74556
rect 112916 74496 112980 74500
rect 112996 74556 113060 74560
rect 112996 74500 113000 74556
rect 113000 74500 113056 74556
rect 113056 74500 113060 74556
rect 112996 74496 113060 74500
rect 113076 74556 113140 74560
rect 113076 74500 113080 74556
rect 113080 74500 113136 74556
rect 113136 74500 113140 74556
rect 113076 74496 113140 74500
rect 113156 74556 113220 74560
rect 113156 74500 113160 74556
rect 113160 74500 113216 74556
rect 113216 74500 113220 74556
rect 113156 74496 113220 74500
rect 4876 74012 4940 74016
rect 4876 73956 4880 74012
rect 4880 73956 4936 74012
rect 4936 73956 4940 74012
rect 4876 73952 4940 73956
rect 4956 74012 5020 74016
rect 4956 73956 4960 74012
rect 4960 73956 5016 74012
rect 5016 73956 5020 74012
rect 4956 73952 5020 73956
rect 5036 74012 5100 74016
rect 5036 73956 5040 74012
rect 5040 73956 5096 74012
rect 5096 73956 5100 74012
rect 5036 73952 5100 73956
rect 5116 74012 5180 74016
rect 5116 73956 5120 74012
rect 5120 73956 5176 74012
rect 5176 73956 5180 74012
rect 5116 73952 5180 73956
rect 113652 74012 113716 74016
rect 113652 73956 113656 74012
rect 113656 73956 113712 74012
rect 113712 73956 113716 74012
rect 113652 73952 113716 73956
rect 113732 74012 113796 74016
rect 113732 73956 113736 74012
rect 113736 73956 113792 74012
rect 113792 73956 113796 74012
rect 113732 73952 113796 73956
rect 113812 74012 113876 74016
rect 113812 73956 113816 74012
rect 113816 73956 113872 74012
rect 113872 73956 113876 74012
rect 113812 73952 113876 73956
rect 113892 74012 113956 74016
rect 113892 73956 113896 74012
rect 113896 73956 113952 74012
rect 113952 73956 113956 74012
rect 113892 73952 113956 73956
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 112916 73468 112980 73472
rect 112916 73412 112920 73468
rect 112920 73412 112976 73468
rect 112976 73412 112980 73468
rect 112916 73408 112980 73412
rect 112996 73468 113060 73472
rect 112996 73412 113000 73468
rect 113000 73412 113056 73468
rect 113056 73412 113060 73468
rect 112996 73408 113060 73412
rect 113076 73468 113140 73472
rect 113076 73412 113080 73468
rect 113080 73412 113136 73468
rect 113136 73412 113140 73468
rect 113076 73408 113140 73412
rect 113156 73468 113220 73472
rect 113156 73412 113160 73468
rect 113160 73412 113216 73468
rect 113216 73412 113220 73468
rect 113156 73408 113220 73412
rect 4876 72924 4940 72928
rect 4876 72868 4880 72924
rect 4880 72868 4936 72924
rect 4936 72868 4940 72924
rect 4876 72864 4940 72868
rect 4956 72924 5020 72928
rect 4956 72868 4960 72924
rect 4960 72868 5016 72924
rect 5016 72868 5020 72924
rect 4956 72864 5020 72868
rect 5036 72924 5100 72928
rect 5036 72868 5040 72924
rect 5040 72868 5096 72924
rect 5096 72868 5100 72924
rect 5036 72864 5100 72868
rect 5116 72924 5180 72928
rect 5116 72868 5120 72924
rect 5120 72868 5176 72924
rect 5176 72868 5180 72924
rect 5116 72864 5180 72868
rect 113652 72924 113716 72928
rect 113652 72868 113656 72924
rect 113656 72868 113712 72924
rect 113712 72868 113716 72924
rect 113652 72864 113716 72868
rect 113732 72924 113796 72928
rect 113732 72868 113736 72924
rect 113736 72868 113792 72924
rect 113792 72868 113796 72924
rect 113732 72864 113796 72868
rect 113812 72924 113876 72928
rect 113812 72868 113816 72924
rect 113816 72868 113872 72924
rect 113872 72868 113876 72924
rect 113812 72864 113876 72868
rect 113892 72924 113956 72928
rect 113892 72868 113896 72924
rect 113896 72868 113952 72924
rect 113952 72868 113956 72924
rect 113892 72864 113956 72868
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 112916 72380 112980 72384
rect 112916 72324 112920 72380
rect 112920 72324 112976 72380
rect 112976 72324 112980 72380
rect 112916 72320 112980 72324
rect 112996 72380 113060 72384
rect 112996 72324 113000 72380
rect 113000 72324 113056 72380
rect 113056 72324 113060 72380
rect 112996 72320 113060 72324
rect 113076 72380 113140 72384
rect 113076 72324 113080 72380
rect 113080 72324 113136 72380
rect 113136 72324 113140 72380
rect 113076 72320 113140 72324
rect 113156 72380 113220 72384
rect 113156 72324 113160 72380
rect 113160 72324 113216 72380
rect 113216 72324 113220 72380
rect 113156 72320 113220 72324
rect 4876 71836 4940 71840
rect 4876 71780 4880 71836
rect 4880 71780 4936 71836
rect 4936 71780 4940 71836
rect 4876 71776 4940 71780
rect 4956 71836 5020 71840
rect 4956 71780 4960 71836
rect 4960 71780 5016 71836
rect 5016 71780 5020 71836
rect 4956 71776 5020 71780
rect 5036 71836 5100 71840
rect 5036 71780 5040 71836
rect 5040 71780 5096 71836
rect 5096 71780 5100 71836
rect 5036 71776 5100 71780
rect 5116 71836 5180 71840
rect 5116 71780 5120 71836
rect 5120 71780 5176 71836
rect 5176 71780 5180 71836
rect 5116 71776 5180 71780
rect 113652 71836 113716 71840
rect 113652 71780 113656 71836
rect 113656 71780 113712 71836
rect 113712 71780 113716 71836
rect 113652 71776 113716 71780
rect 113732 71836 113796 71840
rect 113732 71780 113736 71836
rect 113736 71780 113792 71836
rect 113792 71780 113796 71836
rect 113732 71776 113796 71780
rect 113812 71836 113876 71840
rect 113812 71780 113816 71836
rect 113816 71780 113872 71836
rect 113872 71780 113876 71836
rect 113812 71776 113876 71780
rect 113892 71836 113956 71840
rect 113892 71780 113896 71836
rect 113896 71780 113952 71836
rect 113952 71780 113956 71836
rect 113892 71776 113956 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 112916 71292 112980 71296
rect 112916 71236 112920 71292
rect 112920 71236 112976 71292
rect 112976 71236 112980 71292
rect 112916 71232 112980 71236
rect 112996 71292 113060 71296
rect 112996 71236 113000 71292
rect 113000 71236 113056 71292
rect 113056 71236 113060 71292
rect 112996 71232 113060 71236
rect 113076 71292 113140 71296
rect 113076 71236 113080 71292
rect 113080 71236 113136 71292
rect 113136 71236 113140 71292
rect 113076 71232 113140 71236
rect 113156 71292 113220 71296
rect 113156 71236 113160 71292
rect 113160 71236 113216 71292
rect 113216 71236 113220 71292
rect 113156 71232 113220 71236
rect 4876 70748 4940 70752
rect 4876 70692 4880 70748
rect 4880 70692 4936 70748
rect 4936 70692 4940 70748
rect 4876 70688 4940 70692
rect 4956 70748 5020 70752
rect 4956 70692 4960 70748
rect 4960 70692 5016 70748
rect 5016 70692 5020 70748
rect 4956 70688 5020 70692
rect 5036 70748 5100 70752
rect 5036 70692 5040 70748
rect 5040 70692 5096 70748
rect 5096 70692 5100 70748
rect 5036 70688 5100 70692
rect 5116 70748 5180 70752
rect 5116 70692 5120 70748
rect 5120 70692 5176 70748
rect 5176 70692 5180 70748
rect 5116 70688 5180 70692
rect 113652 70748 113716 70752
rect 113652 70692 113656 70748
rect 113656 70692 113712 70748
rect 113712 70692 113716 70748
rect 113652 70688 113716 70692
rect 113732 70748 113796 70752
rect 113732 70692 113736 70748
rect 113736 70692 113792 70748
rect 113792 70692 113796 70748
rect 113732 70688 113796 70692
rect 113812 70748 113876 70752
rect 113812 70692 113816 70748
rect 113816 70692 113872 70748
rect 113872 70692 113876 70748
rect 113812 70688 113876 70692
rect 113892 70748 113956 70752
rect 113892 70692 113896 70748
rect 113896 70692 113952 70748
rect 113952 70692 113956 70748
rect 113892 70688 113956 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 112916 70204 112980 70208
rect 112916 70148 112920 70204
rect 112920 70148 112976 70204
rect 112976 70148 112980 70204
rect 112916 70144 112980 70148
rect 112996 70204 113060 70208
rect 112996 70148 113000 70204
rect 113000 70148 113056 70204
rect 113056 70148 113060 70204
rect 112996 70144 113060 70148
rect 113076 70204 113140 70208
rect 113076 70148 113080 70204
rect 113080 70148 113136 70204
rect 113136 70148 113140 70204
rect 113076 70144 113140 70148
rect 113156 70204 113220 70208
rect 113156 70148 113160 70204
rect 113160 70148 113216 70204
rect 113216 70148 113220 70204
rect 113156 70144 113220 70148
rect 4876 69660 4940 69664
rect 4876 69604 4880 69660
rect 4880 69604 4936 69660
rect 4936 69604 4940 69660
rect 4876 69600 4940 69604
rect 4956 69660 5020 69664
rect 4956 69604 4960 69660
rect 4960 69604 5016 69660
rect 5016 69604 5020 69660
rect 4956 69600 5020 69604
rect 5036 69660 5100 69664
rect 5036 69604 5040 69660
rect 5040 69604 5096 69660
rect 5096 69604 5100 69660
rect 5036 69600 5100 69604
rect 5116 69660 5180 69664
rect 5116 69604 5120 69660
rect 5120 69604 5176 69660
rect 5176 69604 5180 69660
rect 5116 69600 5180 69604
rect 113652 69660 113716 69664
rect 113652 69604 113656 69660
rect 113656 69604 113712 69660
rect 113712 69604 113716 69660
rect 113652 69600 113716 69604
rect 113732 69660 113796 69664
rect 113732 69604 113736 69660
rect 113736 69604 113792 69660
rect 113792 69604 113796 69660
rect 113732 69600 113796 69604
rect 113812 69660 113876 69664
rect 113812 69604 113816 69660
rect 113816 69604 113872 69660
rect 113872 69604 113876 69660
rect 113812 69600 113876 69604
rect 113892 69660 113956 69664
rect 113892 69604 113896 69660
rect 113896 69604 113952 69660
rect 113952 69604 113956 69660
rect 113892 69600 113956 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 112916 69116 112980 69120
rect 112916 69060 112920 69116
rect 112920 69060 112976 69116
rect 112976 69060 112980 69116
rect 112916 69056 112980 69060
rect 112996 69116 113060 69120
rect 112996 69060 113000 69116
rect 113000 69060 113056 69116
rect 113056 69060 113060 69116
rect 112996 69056 113060 69060
rect 113076 69116 113140 69120
rect 113076 69060 113080 69116
rect 113080 69060 113136 69116
rect 113136 69060 113140 69116
rect 113076 69056 113140 69060
rect 113156 69116 113220 69120
rect 113156 69060 113160 69116
rect 113160 69060 113216 69116
rect 113216 69060 113220 69116
rect 113156 69056 113220 69060
rect 4876 68572 4940 68576
rect 4876 68516 4880 68572
rect 4880 68516 4936 68572
rect 4936 68516 4940 68572
rect 4876 68512 4940 68516
rect 4956 68572 5020 68576
rect 4956 68516 4960 68572
rect 4960 68516 5016 68572
rect 5016 68516 5020 68572
rect 4956 68512 5020 68516
rect 5036 68572 5100 68576
rect 5036 68516 5040 68572
rect 5040 68516 5096 68572
rect 5096 68516 5100 68572
rect 5036 68512 5100 68516
rect 5116 68572 5180 68576
rect 5116 68516 5120 68572
rect 5120 68516 5176 68572
rect 5176 68516 5180 68572
rect 5116 68512 5180 68516
rect 113652 68572 113716 68576
rect 113652 68516 113656 68572
rect 113656 68516 113712 68572
rect 113712 68516 113716 68572
rect 113652 68512 113716 68516
rect 113732 68572 113796 68576
rect 113732 68516 113736 68572
rect 113736 68516 113792 68572
rect 113792 68516 113796 68572
rect 113732 68512 113796 68516
rect 113812 68572 113876 68576
rect 113812 68516 113816 68572
rect 113816 68516 113872 68572
rect 113872 68516 113876 68572
rect 113812 68512 113876 68516
rect 113892 68572 113956 68576
rect 113892 68516 113896 68572
rect 113896 68516 113952 68572
rect 113952 68516 113956 68572
rect 113892 68512 113956 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 112916 68028 112980 68032
rect 112916 67972 112920 68028
rect 112920 67972 112976 68028
rect 112976 67972 112980 68028
rect 112916 67968 112980 67972
rect 112996 68028 113060 68032
rect 112996 67972 113000 68028
rect 113000 67972 113056 68028
rect 113056 67972 113060 68028
rect 112996 67968 113060 67972
rect 113076 68028 113140 68032
rect 113076 67972 113080 68028
rect 113080 67972 113136 68028
rect 113136 67972 113140 68028
rect 113076 67968 113140 67972
rect 113156 68028 113220 68032
rect 113156 67972 113160 68028
rect 113160 67972 113216 68028
rect 113216 67972 113220 68028
rect 113156 67968 113220 67972
rect 4876 67484 4940 67488
rect 4876 67428 4880 67484
rect 4880 67428 4936 67484
rect 4936 67428 4940 67484
rect 4876 67424 4940 67428
rect 4956 67484 5020 67488
rect 4956 67428 4960 67484
rect 4960 67428 5016 67484
rect 5016 67428 5020 67484
rect 4956 67424 5020 67428
rect 5036 67484 5100 67488
rect 5036 67428 5040 67484
rect 5040 67428 5096 67484
rect 5096 67428 5100 67484
rect 5036 67424 5100 67428
rect 5116 67484 5180 67488
rect 5116 67428 5120 67484
rect 5120 67428 5176 67484
rect 5176 67428 5180 67484
rect 5116 67424 5180 67428
rect 113652 67484 113716 67488
rect 113652 67428 113656 67484
rect 113656 67428 113712 67484
rect 113712 67428 113716 67484
rect 113652 67424 113716 67428
rect 113732 67484 113796 67488
rect 113732 67428 113736 67484
rect 113736 67428 113792 67484
rect 113792 67428 113796 67484
rect 113732 67424 113796 67428
rect 113812 67484 113876 67488
rect 113812 67428 113816 67484
rect 113816 67428 113872 67484
rect 113872 67428 113876 67484
rect 113812 67424 113876 67428
rect 113892 67484 113956 67488
rect 113892 67428 113896 67484
rect 113896 67428 113952 67484
rect 113952 67428 113956 67484
rect 113892 67424 113956 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 112916 66940 112980 66944
rect 112916 66884 112920 66940
rect 112920 66884 112976 66940
rect 112976 66884 112980 66940
rect 112916 66880 112980 66884
rect 112996 66940 113060 66944
rect 112996 66884 113000 66940
rect 113000 66884 113056 66940
rect 113056 66884 113060 66940
rect 112996 66880 113060 66884
rect 113076 66940 113140 66944
rect 113076 66884 113080 66940
rect 113080 66884 113136 66940
rect 113136 66884 113140 66940
rect 113076 66880 113140 66884
rect 113156 66940 113220 66944
rect 113156 66884 113160 66940
rect 113160 66884 113216 66940
rect 113216 66884 113220 66940
rect 113156 66880 113220 66884
rect 4876 66396 4940 66400
rect 4876 66340 4880 66396
rect 4880 66340 4936 66396
rect 4936 66340 4940 66396
rect 4876 66336 4940 66340
rect 4956 66396 5020 66400
rect 4956 66340 4960 66396
rect 4960 66340 5016 66396
rect 5016 66340 5020 66396
rect 4956 66336 5020 66340
rect 5036 66396 5100 66400
rect 5036 66340 5040 66396
rect 5040 66340 5096 66396
rect 5096 66340 5100 66396
rect 5036 66336 5100 66340
rect 5116 66396 5180 66400
rect 5116 66340 5120 66396
rect 5120 66340 5176 66396
rect 5176 66340 5180 66396
rect 5116 66336 5180 66340
rect 113652 66396 113716 66400
rect 113652 66340 113656 66396
rect 113656 66340 113712 66396
rect 113712 66340 113716 66396
rect 113652 66336 113716 66340
rect 113732 66396 113796 66400
rect 113732 66340 113736 66396
rect 113736 66340 113792 66396
rect 113792 66340 113796 66396
rect 113732 66336 113796 66340
rect 113812 66396 113876 66400
rect 113812 66340 113816 66396
rect 113816 66340 113872 66396
rect 113872 66340 113876 66396
rect 113812 66336 113876 66340
rect 113892 66396 113956 66400
rect 113892 66340 113896 66396
rect 113896 66340 113952 66396
rect 113952 66340 113956 66396
rect 113892 66336 113956 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 112916 65852 112980 65856
rect 112916 65796 112920 65852
rect 112920 65796 112976 65852
rect 112976 65796 112980 65852
rect 112916 65792 112980 65796
rect 112996 65852 113060 65856
rect 112996 65796 113000 65852
rect 113000 65796 113056 65852
rect 113056 65796 113060 65852
rect 112996 65792 113060 65796
rect 113076 65852 113140 65856
rect 113076 65796 113080 65852
rect 113080 65796 113136 65852
rect 113136 65796 113140 65852
rect 113076 65792 113140 65796
rect 113156 65852 113220 65856
rect 113156 65796 113160 65852
rect 113160 65796 113216 65852
rect 113216 65796 113220 65852
rect 113156 65792 113220 65796
rect 4876 65308 4940 65312
rect 4876 65252 4880 65308
rect 4880 65252 4936 65308
rect 4936 65252 4940 65308
rect 4876 65248 4940 65252
rect 4956 65308 5020 65312
rect 4956 65252 4960 65308
rect 4960 65252 5016 65308
rect 5016 65252 5020 65308
rect 4956 65248 5020 65252
rect 5036 65308 5100 65312
rect 5036 65252 5040 65308
rect 5040 65252 5096 65308
rect 5096 65252 5100 65308
rect 5036 65248 5100 65252
rect 5116 65308 5180 65312
rect 5116 65252 5120 65308
rect 5120 65252 5176 65308
rect 5176 65252 5180 65308
rect 5116 65248 5180 65252
rect 113652 65308 113716 65312
rect 113652 65252 113656 65308
rect 113656 65252 113712 65308
rect 113712 65252 113716 65308
rect 113652 65248 113716 65252
rect 113732 65308 113796 65312
rect 113732 65252 113736 65308
rect 113736 65252 113792 65308
rect 113792 65252 113796 65308
rect 113732 65248 113796 65252
rect 113812 65308 113876 65312
rect 113812 65252 113816 65308
rect 113816 65252 113872 65308
rect 113872 65252 113876 65308
rect 113812 65248 113876 65252
rect 113892 65308 113956 65312
rect 113892 65252 113896 65308
rect 113896 65252 113952 65308
rect 113952 65252 113956 65308
rect 113892 65248 113956 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 112916 64764 112980 64768
rect 112916 64708 112920 64764
rect 112920 64708 112976 64764
rect 112976 64708 112980 64764
rect 112916 64704 112980 64708
rect 112996 64764 113060 64768
rect 112996 64708 113000 64764
rect 113000 64708 113056 64764
rect 113056 64708 113060 64764
rect 112996 64704 113060 64708
rect 113076 64764 113140 64768
rect 113076 64708 113080 64764
rect 113080 64708 113136 64764
rect 113136 64708 113140 64764
rect 113076 64704 113140 64708
rect 113156 64764 113220 64768
rect 113156 64708 113160 64764
rect 113160 64708 113216 64764
rect 113216 64708 113220 64764
rect 113156 64704 113220 64708
rect 4876 64220 4940 64224
rect 4876 64164 4880 64220
rect 4880 64164 4936 64220
rect 4936 64164 4940 64220
rect 4876 64160 4940 64164
rect 4956 64220 5020 64224
rect 4956 64164 4960 64220
rect 4960 64164 5016 64220
rect 5016 64164 5020 64220
rect 4956 64160 5020 64164
rect 5036 64220 5100 64224
rect 5036 64164 5040 64220
rect 5040 64164 5096 64220
rect 5096 64164 5100 64220
rect 5036 64160 5100 64164
rect 5116 64220 5180 64224
rect 5116 64164 5120 64220
rect 5120 64164 5176 64220
rect 5176 64164 5180 64220
rect 5116 64160 5180 64164
rect 113652 64220 113716 64224
rect 113652 64164 113656 64220
rect 113656 64164 113712 64220
rect 113712 64164 113716 64220
rect 113652 64160 113716 64164
rect 113732 64220 113796 64224
rect 113732 64164 113736 64220
rect 113736 64164 113792 64220
rect 113792 64164 113796 64220
rect 113732 64160 113796 64164
rect 113812 64220 113876 64224
rect 113812 64164 113816 64220
rect 113816 64164 113872 64220
rect 113872 64164 113876 64220
rect 113812 64160 113876 64164
rect 113892 64220 113956 64224
rect 113892 64164 113896 64220
rect 113896 64164 113952 64220
rect 113952 64164 113956 64220
rect 113892 64160 113956 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 112916 63676 112980 63680
rect 112916 63620 112920 63676
rect 112920 63620 112976 63676
rect 112976 63620 112980 63676
rect 112916 63616 112980 63620
rect 112996 63676 113060 63680
rect 112996 63620 113000 63676
rect 113000 63620 113056 63676
rect 113056 63620 113060 63676
rect 112996 63616 113060 63620
rect 113076 63676 113140 63680
rect 113076 63620 113080 63676
rect 113080 63620 113136 63676
rect 113136 63620 113140 63676
rect 113076 63616 113140 63620
rect 113156 63676 113220 63680
rect 113156 63620 113160 63676
rect 113160 63620 113216 63676
rect 113216 63620 113220 63676
rect 113156 63616 113220 63620
rect 4876 63132 4940 63136
rect 4876 63076 4880 63132
rect 4880 63076 4936 63132
rect 4936 63076 4940 63132
rect 4876 63072 4940 63076
rect 4956 63132 5020 63136
rect 4956 63076 4960 63132
rect 4960 63076 5016 63132
rect 5016 63076 5020 63132
rect 4956 63072 5020 63076
rect 5036 63132 5100 63136
rect 5036 63076 5040 63132
rect 5040 63076 5096 63132
rect 5096 63076 5100 63132
rect 5036 63072 5100 63076
rect 5116 63132 5180 63136
rect 5116 63076 5120 63132
rect 5120 63076 5176 63132
rect 5176 63076 5180 63132
rect 5116 63072 5180 63076
rect 113652 63132 113716 63136
rect 113652 63076 113656 63132
rect 113656 63076 113712 63132
rect 113712 63076 113716 63132
rect 113652 63072 113716 63076
rect 113732 63132 113796 63136
rect 113732 63076 113736 63132
rect 113736 63076 113792 63132
rect 113792 63076 113796 63132
rect 113732 63072 113796 63076
rect 113812 63132 113876 63136
rect 113812 63076 113816 63132
rect 113816 63076 113872 63132
rect 113872 63076 113876 63132
rect 113812 63072 113876 63076
rect 113892 63132 113956 63136
rect 113892 63076 113896 63132
rect 113896 63076 113952 63132
rect 113952 63076 113956 63132
rect 113892 63072 113956 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 112916 62588 112980 62592
rect 112916 62532 112920 62588
rect 112920 62532 112976 62588
rect 112976 62532 112980 62588
rect 112916 62528 112980 62532
rect 112996 62588 113060 62592
rect 112996 62532 113000 62588
rect 113000 62532 113056 62588
rect 113056 62532 113060 62588
rect 112996 62528 113060 62532
rect 113076 62588 113140 62592
rect 113076 62532 113080 62588
rect 113080 62532 113136 62588
rect 113136 62532 113140 62588
rect 113076 62528 113140 62532
rect 113156 62588 113220 62592
rect 113156 62532 113160 62588
rect 113160 62532 113216 62588
rect 113216 62532 113220 62588
rect 113156 62528 113220 62532
rect 4876 62044 4940 62048
rect 4876 61988 4880 62044
rect 4880 61988 4936 62044
rect 4936 61988 4940 62044
rect 4876 61984 4940 61988
rect 4956 62044 5020 62048
rect 4956 61988 4960 62044
rect 4960 61988 5016 62044
rect 5016 61988 5020 62044
rect 4956 61984 5020 61988
rect 5036 62044 5100 62048
rect 5036 61988 5040 62044
rect 5040 61988 5096 62044
rect 5096 61988 5100 62044
rect 5036 61984 5100 61988
rect 5116 62044 5180 62048
rect 5116 61988 5120 62044
rect 5120 61988 5176 62044
rect 5176 61988 5180 62044
rect 5116 61984 5180 61988
rect 113652 62044 113716 62048
rect 113652 61988 113656 62044
rect 113656 61988 113712 62044
rect 113712 61988 113716 62044
rect 113652 61984 113716 61988
rect 113732 62044 113796 62048
rect 113732 61988 113736 62044
rect 113736 61988 113792 62044
rect 113792 61988 113796 62044
rect 113732 61984 113796 61988
rect 113812 62044 113876 62048
rect 113812 61988 113816 62044
rect 113816 61988 113872 62044
rect 113872 61988 113876 62044
rect 113812 61984 113876 61988
rect 113892 62044 113956 62048
rect 113892 61988 113896 62044
rect 113896 61988 113952 62044
rect 113952 61988 113956 62044
rect 113892 61984 113956 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 112916 61500 112980 61504
rect 112916 61444 112920 61500
rect 112920 61444 112976 61500
rect 112976 61444 112980 61500
rect 112916 61440 112980 61444
rect 112996 61500 113060 61504
rect 112996 61444 113000 61500
rect 113000 61444 113056 61500
rect 113056 61444 113060 61500
rect 112996 61440 113060 61444
rect 113076 61500 113140 61504
rect 113076 61444 113080 61500
rect 113080 61444 113136 61500
rect 113136 61444 113140 61500
rect 113076 61440 113140 61444
rect 113156 61500 113220 61504
rect 113156 61444 113160 61500
rect 113160 61444 113216 61500
rect 113216 61444 113220 61500
rect 113156 61440 113220 61444
rect 4876 60956 4940 60960
rect 4876 60900 4880 60956
rect 4880 60900 4936 60956
rect 4936 60900 4940 60956
rect 4876 60896 4940 60900
rect 4956 60956 5020 60960
rect 4956 60900 4960 60956
rect 4960 60900 5016 60956
rect 5016 60900 5020 60956
rect 4956 60896 5020 60900
rect 5036 60956 5100 60960
rect 5036 60900 5040 60956
rect 5040 60900 5096 60956
rect 5096 60900 5100 60956
rect 5036 60896 5100 60900
rect 5116 60956 5180 60960
rect 5116 60900 5120 60956
rect 5120 60900 5176 60956
rect 5176 60900 5180 60956
rect 5116 60896 5180 60900
rect 113652 60956 113716 60960
rect 113652 60900 113656 60956
rect 113656 60900 113712 60956
rect 113712 60900 113716 60956
rect 113652 60896 113716 60900
rect 113732 60956 113796 60960
rect 113732 60900 113736 60956
rect 113736 60900 113792 60956
rect 113792 60900 113796 60956
rect 113732 60896 113796 60900
rect 113812 60956 113876 60960
rect 113812 60900 113816 60956
rect 113816 60900 113872 60956
rect 113872 60900 113876 60956
rect 113812 60896 113876 60900
rect 113892 60956 113956 60960
rect 113892 60900 113896 60956
rect 113896 60900 113952 60956
rect 113952 60900 113956 60956
rect 113892 60896 113956 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 112916 60412 112980 60416
rect 112916 60356 112920 60412
rect 112920 60356 112976 60412
rect 112976 60356 112980 60412
rect 112916 60352 112980 60356
rect 112996 60412 113060 60416
rect 112996 60356 113000 60412
rect 113000 60356 113056 60412
rect 113056 60356 113060 60412
rect 112996 60352 113060 60356
rect 113076 60412 113140 60416
rect 113076 60356 113080 60412
rect 113080 60356 113136 60412
rect 113136 60356 113140 60412
rect 113076 60352 113140 60356
rect 113156 60412 113220 60416
rect 113156 60356 113160 60412
rect 113160 60356 113216 60412
rect 113216 60356 113220 60412
rect 113156 60352 113220 60356
rect 4876 59868 4940 59872
rect 4876 59812 4880 59868
rect 4880 59812 4936 59868
rect 4936 59812 4940 59868
rect 4876 59808 4940 59812
rect 4956 59868 5020 59872
rect 4956 59812 4960 59868
rect 4960 59812 5016 59868
rect 5016 59812 5020 59868
rect 4956 59808 5020 59812
rect 5036 59868 5100 59872
rect 5036 59812 5040 59868
rect 5040 59812 5096 59868
rect 5096 59812 5100 59868
rect 5036 59808 5100 59812
rect 5116 59868 5180 59872
rect 5116 59812 5120 59868
rect 5120 59812 5176 59868
rect 5176 59812 5180 59868
rect 5116 59808 5180 59812
rect 113652 59868 113716 59872
rect 113652 59812 113656 59868
rect 113656 59812 113712 59868
rect 113712 59812 113716 59868
rect 113652 59808 113716 59812
rect 113732 59868 113796 59872
rect 113732 59812 113736 59868
rect 113736 59812 113792 59868
rect 113792 59812 113796 59868
rect 113732 59808 113796 59812
rect 113812 59868 113876 59872
rect 113812 59812 113816 59868
rect 113816 59812 113872 59868
rect 113872 59812 113876 59868
rect 113812 59808 113876 59812
rect 113892 59868 113956 59872
rect 113892 59812 113896 59868
rect 113896 59812 113952 59868
rect 113952 59812 113956 59868
rect 113892 59808 113956 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 112916 59324 112980 59328
rect 112916 59268 112920 59324
rect 112920 59268 112976 59324
rect 112976 59268 112980 59324
rect 112916 59264 112980 59268
rect 112996 59324 113060 59328
rect 112996 59268 113000 59324
rect 113000 59268 113056 59324
rect 113056 59268 113060 59324
rect 112996 59264 113060 59268
rect 113076 59324 113140 59328
rect 113076 59268 113080 59324
rect 113080 59268 113136 59324
rect 113136 59268 113140 59324
rect 113076 59264 113140 59268
rect 113156 59324 113220 59328
rect 113156 59268 113160 59324
rect 113160 59268 113216 59324
rect 113216 59268 113220 59324
rect 113156 59264 113220 59268
rect 4876 58780 4940 58784
rect 4876 58724 4880 58780
rect 4880 58724 4936 58780
rect 4936 58724 4940 58780
rect 4876 58720 4940 58724
rect 4956 58780 5020 58784
rect 4956 58724 4960 58780
rect 4960 58724 5016 58780
rect 5016 58724 5020 58780
rect 4956 58720 5020 58724
rect 5036 58780 5100 58784
rect 5036 58724 5040 58780
rect 5040 58724 5096 58780
rect 5096 58724 5100 58780
rect 5036 58720 5100 58724
rect 5116 58780 5180 58784
rect 5116 58724 5120 58780
rect 5120 58724 5176 58780
rect 5176 58724 5180 58780
rect 5116 58720 5180 58724
rect 113652 58780 113716 58784
rect 113652 58724 113656 58780
rect 113656 58724 113712 58780
rect 113712 58724 113716 58780
rect 113652 58720 113716 58724
rect 113732 58780 113796 58784
rect 113732 58724 113736 58780
rect 113736 58724 113792 58780
rect 113792 58724 113796 58780
rect 113732 58720 113796 58724
rect 113812 58780 113876 58784
rect 113812 58724 113816 58780
rect 113816 58724 113872 58780
rect 113872 58724 113876 58780
rect 113812 58720 113876 58724
rect 113892 58780 113956 58784
rect 113892 58724 113896 58780
rect 113896 58724 113952 58780
rect 113952 58724 113956 58780
rect 113892 58720 113956 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 112916 58236 112980 58240
rect 112916 58180 112920 58236
rect 112920 58180 112976 58236
rect 112976 58180 112980 58236
rect 112916 58176 112980 58180
rect 112996 58236 113060 58240
rect 112996 58180 113000 58236
rect 113000 58180 113056 58236
rect 113056 58180 113060 58236
rect 112996 58176 113060 58180
rect 113076 58236 113140 58240
rect 113076 58180 113080 58236
rect 113080 58180 113136 58236
rect 113136 58180 113140 58236
rect 113076 58176 113140 58180
rect 113156 58236 113220 58240
rect 113156 58180 113160 58236
rect 113160 58180 113216 58236
rect 113216 58180 113220 58236
rect 113156 58176 113220 58180
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 113652 57692 113716 57696
rect 113652 57636 113656 57692
rect 113656 57636 113712 57692
rect 113712 57636 113716 57692
rect 113652 57632 113716 57636
rect 113732 57692 113796 57696
rect 113732 57636 113736 57692
rect 113736 57636 113792 57692
rect 113792 57636 113796 57692
rect 113732 57632 113796 57636
rect 113812 57692 113876 57696
rect 113812 57636 113816 57692
rect 113816 57636 113872 57692
rect 113872 57636 113876 57692
rect 113812 57632 113876 57636
rect 113892 57692 113956 57696
rect 113892 57636 113896 57692
rect 113896 57636 113952 57692
rect 113952 57636 113956 57692
rect 113892 57632 113956 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 112916 57148 112980 57152
rect 112916 57092 112920 57148
rect 112920 57092 112976 57148
rect 112976 57092 112980 57148
rect 112916 57088 112980 57092
rect 112996 57148 113060 57152
rect 112996 57092 113000 57148
rect 113000 57092 113056 57148
rect 113056 57092 113060 57148
rect 112996 57088 113060 57092
rect 113076 57148 113140 57152
rect 113076 57092 113080 57148
rect 113080 57092 113136 57148
rect 113136 57092 113140 57148
rect 113076 57088 113140 57092
rect 113156 57148 113220 57152
rect 113156 57092 113160 57148
rect 113160 57092 113216 57148
rect 113216 57092 113220 57148
rect 113156 57088 113220 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 113652 56604 113716 56608
rect 113652 56548 113656 56604
rect 113656 56548 113712 56604
rect 113712 56548 113716 56604
rect 113652 56544 113716 56548
rect 113732 56604 113796 56608
rect 113732 56548 113736 56604
rect 113736 56548 113792 56604
rect 113792 56548 113796 56604
rect 113732 56544 113796 56548
rect 113812 56604 113876 56608
rect 113812 56548 113816 56604
rect 113816 56548 113872 56604
rect 113872 56548 113876 56604
rect 113812 56544 113876 56548
rect 113892 56604 113956 56608
rect 113892 56548 113896 56604
rect 113896 56548 113952 56604
rect 113952 56548 113956 56604
rect 113892 56544 113956 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 112916 56060 112980 56064
rect 112916 56004 112920 56060
rect 112920 56004 112976 56060
rect 112976 56004 112980 56060
rect 112916 56000 112980 56004
rect 112996 56060 113060 56064
rect 112996 56004 113000 56060
rect 113000 56004 113056 56060
rect 113056 56004 113060 56060
rect 112996 56000 113060 56004
rect 113076 56060 113140 56064
rect 113076 56004 113080 56060
rect 113080 56004 113136 56060
rect 113136 56004 113140 56060
rect 113076 56000 113140 56004
rect 113156 56060 113220 56064
rect 113156 56004 113160 56060
rect 113160 56004 113216 56060
rect 113216 56004 113220 56060
rect 113156 56000 113220 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 113652 55516 113716 55520
rect 113652 55460 113656 55516
rect 113656 55460 113712 55516
rect 113712 55460 113716 55516
rect 113652 55456 113716 55460
rect 113732 55516 113796 55520
rect 113732 55460 113736 55516
rect 113736 55460 113792 55516
rect 113792 55460 113796 55516
rect 113732 55456 113796 55460
rect 113812 55516 113876 55520
rect 113812 55460 113816 55516
rect 113816 55460 113872 55516
rect 113872 55460 113876 55516
rect 113812 55456 113876 55460
rect 113892 55516 113956 55520
rect 113892 55460 113896 55516
rect 113896 55460 113952 55516
rect 113952 55460 113956 55516
rect 113892 55456 113956 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 112916 54972 112980 54976
rect 112916 54916 112920 54972
rect 112920 54916 112976 54972
rect 112976 54916 112980 54972
rect 112916 54912 112980 54916
rect 112996 54972 113060 54976
rect 112996 54916 113000 54972
rect 113000 54916 113056 54972
rect 113056 54916 113060 54972
rect 112996 54912 113060 54916
rect 113076 54972 113140 54976
rect 113076 54916 113080 54972
rect 113080 54916 113136 54972
rect 113136 54916 113140 54972
rect 113076 54912 113140 54916
rect 113156 54972 113220 54976
rect 113156 54916 113160 54972
rect 113160 54916 113216 54972
rect 113216 54916 113220 54972
rect 113156 54912 113220 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 113652 54428 113716 54432
rect 113652 54372 113656 54428
rect 113656 54372 113712 54428
rect 113712 54372 113716 54428
rect 113652 54368 113716 54372
rect 113732 54428 113796 54432
rect 113732 54372 113736 54428
rect 113736 54372 113792 54428
rect 113792 54372 113796 54428
rect 113732 54368 113796 54372
rect 113812 54428 113876 54432
rect 113812 54372 113816 54428
rect 113816 54372 113872 54428
rect 113872 54372 113876 54428
rect 113812 54368 113876 54372
rect 113892 54428 113956 54432
rect 113892 54372 113896 54428
rect 113896 54372 113952 54428
rect 113952 54372 113956 54428
rect 113892 54368 113956 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 112916 53884 112980 53888
rect 112916 53828 112920 53884
rect 112920 53828 112976 53884
rect 112976 53828 112980 53884
rect 112916 53824 112980 53828
rect 112996 53884 113060 53888
rect 112996 53828 113000 53884
rect 113000 53828 113056 53884
rect 113056 53828 113060 53884
rect 112996 53824 113060 53828
rect 113076 53884 113140 53888
rect 113076 53828 113080 53884
rect 113080 53828 113136 53884
rect 113136 53828 113140 53884
rect 113076 53824 113140 53828
rect 113156 53884 113220 53888
rect 113156 53828 113160 53884
rect 113160 53828 113216 53884
rect 113216 53828 113220 53884
rect 113156 53824 113220 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 113652 53340 113716 53344
rect 113652 53284 113656 53340
rect 113656 53284 113712 53340
rect 113712 53284 113716 53340
rect 113652 53280 113716 53284
rect 113732 53340 113796 53344
rect 113732 53284 113736 53340
rect 113736 53284 113792 53340
rect 113792 53284 113796 53340
rect 113732 53280 113796 53284
rect 113812 53340 113876 53344
rect 113812 53284 113816 53340
rect 113816 53284 113872 53340
rect 113872 53284 113876 53340
rect 113812 53280 113876 53284
rect 113892 53340 113956 53344
rect 113892 53284 113896 53340
rect 113896 53284 113952 53340
rect 113952 53284 113956 53340
rect 113892 53280 113956 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 112916 52796 112980 52800
rect 112916 52740 112920 52796
rect 112920 52740 112976 52796
rect 112976 52740 112980 52796
rect 112916 52736 112980 52740
rect 112996 52796 113060 52800
rect 112996 52740 113000 52796
rect 113000 52740 113056 52796
rect 113056 52740 113060 52796
rect 112996 52736 113060 52740
rect 113076 52796 113140 52800
rect 113076 52740 113080 52796
rect 113080 52740 113136 52796
rect 113136 52740 113140 52796
rect 113076 52736 113140 52740
rect 113156 52796 113220 52800
rect 113156 52740 113160 52796
rect 113160 52740 113216 52796
rect 113216 52740 113220 52796
rect 113156 52736 113220 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 113652 52252 113716 52256
rect 113652 52196 113656 52252
rect 113656 52196 113712 52252
rect 113712 52196 113716 52252
rect 113652 52192 113716 52196
rect 113732 52252 113796 52256
rect 113732 52196 113736 52252
rect 113736 52196 113792 52252
rect 113792 52196 113796 52252
rect 113732 52192 113796 52196
rect 113812 52252 113876 52256
rect 113812 52196 113816 52252
rect 113816 52196 113872 52252
rect 113872 52196 113876 52252
rect 113812 52192 113876 52196
rect 113892 52252 113956 52256
rect 113892 52196 113896 52252
rect 113896 52196 113952 52252
rect 113952 52196 113956 52252
rect 113892 52192 113956 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 112916 51708 112980 51712
rect 112916 51652 112920 51708
rect 112920 51652 112976 51708
rect 112976 51652 112980 51708
rect 112916 51648 112980 51652
rect 112996 51708 113060 51712
rect 112996 51652 113000 51708
rect 113000 51652 113056 51708
rect 113056 51652 113060 51708
rect 112996 51648 113060 51652
rect 113076 51708 113140 51712
rect 113076 51652 113080 51708
rect 113080 51652 113136 51708
rect 113136 51652 113140 51708
rect 113076 51648 113140 51652
rect 113156 51708 113220 51712
rect 113156 51652 113160 51708
rect 113160 51652 113216 51708
rect 113216 51652 113220 51708
rect 113156 51648 113220 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 113652 51164 113716 51168
rect 113652 51108 113656 51164
rect 113656 51108 113712 51164
rect 113712 51108 113716 51164
rect 113652 51104 113716 51108
rect 113732 51164 113796 51168
rect 113732 51108 113736 51164
rect 113736 51108 113792 51164
rect 113792 51108 113796 51164
rect 113732 51104 113796 51108
rect 113812 51164 113876 51168
rect 113812 51108 113816 51164
rect 113816 51108 113872 51164
rect 113872 51108 113876 51164
rect 113812 51104 113876 51108
rect 113892 51164 113956 51168
rect 113892 51108 113896 51164
rect 113896 51108 113952 51164
rect 113952 51108 113956 51164
rect 113892 51104 113956 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 112916 50620 112980 50624
rect 112916 50564 112920 50620
rect 112920 50564 112976 50620
rect 112976 50564 112980 50620
rect 112916 50560 112980 50564
rect 112996 50620 113060 50624
rect 112996 50564 113000 50620
rect 113000 50564 113056 50620
rect 113056 50564 113060 50620
rect 112996 50560 113060 50564
rect 113076 50620 113140 50624
rect 113076 50564 113080 50620
rect 113080 50564 113136 50620
rect 113136 50564 113140 50620
rect 113076 50560 113140 50564
rect 113156 50620 113220 50624
rect 113156 50564 113160 50620
rect 113160 50564 113216 50620
rect 113216 50564 113220 50620
rect 113156 50560 113220 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 113652 50076 113716 50080
rect 113652 50020 113656 50076
rect 113656 50020 113712 50076
rect 113712 50020 113716 50076
rect 113652 50016 113716 50020
rect 113732 50076 113796 50080
rect 113732 50020 113736 50076
rect 113736 50020 113792 50076
rect 113792 50020 113796 50076
rect 113732 50016 113796 50020
rect 113812 50076 113876 50080
rect 113812 50020 113816 50076
rect 113816 50020 113872 50076
rect 113872 50020 113876 50076
rect 113812 50016 113876 50020
rect 113892 50076 113956 50080
rect 113892 50020 113896 50076
rect 113896 50020 113952 50076
rect 113952 50020 113956 50076
rect 113892 50016 113956 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 112916 49532 112980 49536
rect 112916 49476 112920 49532
rect 112920 49476 112976 49532
rect 112976 49476 112980 49532
rect 112916 49472 112980 49476
rect 112996 49532 113060 49536
rect 112996 49476 113000 49532
rect 113000 49476 113056 49532
rect 113056 49476 113060 49532
rect 112996 49472 113060 49476
rect 113076 49532 113140 49536
rect 113076 49476 113080 49532
rect 113080 49476 113136 49532
rect 113136 49476 113140 49532
rect 113076 49472 113140 49476
rect 113156 49532 113220 49536
rect 113156 49476 113160 49532
rect 113160 49476 113216 49532
rect 113216 49476 113220 49532
rect 113156 49472 113220 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 113652 48988 113716 48992
rect 113652 48932 113656 48988
rect 113656 48932 113712 48988
rect 113712 48932 113716 48988
rect 113652 48928 113716 48932
rect 113732 48988 113796 48992
rect 113732 48932 113736 48988
rect 113736 48932 113792 48988
rect 113792 48932 113796 48988
rect 113732 48928 113796 48932
rect 113812 48988 113876 48992
rect 113812 48932 113816 48988
rect 113816 48932 113872 48988
rect 113872 48932 113876 48988
rect 113812 48928 113876 48932
rect 113892 48988 113956 48992
rect 113892 48932 113896 48988
rect 113896 48932 113952 48988
rect 113952 48932 113956 48988
rect 113892 48928 113956 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 112916 48444 112980 48448
rect 112916 48388 112920 48444
rect 112920 48388 112976 48444
rect 112976 48388 112980 48444
rect 112916 48384 112980 48388
rect 112996 48444 113060 48448
rect 112996 48388 113000 48444
rect 113000 48388 113056 48444
rect 113056 48388 113060 48444
rect 112996 48384 113060 48388
rect 113076 48444 113140 48448
rect 113076 48388 113080 48444
rect 113080 48388 113136 48444
rect 113136 48388 113140 48444
rect 113076 48384 113140 48388
rect 113156 48444 113220 48448
rect 113156 48388 113160 48444
rect 113160 48388 113216 48444
rect 113216 48388 113220 48444
rect 113156 48384 113220 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 113652 47900 113716 47904
rect 113652 47844 113656 47900
rect 113656 47844 113712 47900
rect 113712 47844 113716 47900
rect 113652 47840 113716 47844
rect 113732 47900 113796 47904
rect 113732 47844 113736 47900
rect 113736 47844 113792 47900
rect 113792 47844 113796 47900
rect 113732 47840 113796 47844
rect 113812 47900 113876 47904
rect 113812 47844 113816 47900
rect 113816 47844 113872 47900
rect 113872 47844 113876 47900
rect 113812 47840 113876 47844
rect 113892 47900 113956 47904
rect 113892 47844 113896 47900
rect 113896 47844 113952 47900
rect 113952 47844 113956 47900
rect 113892 47840 113956 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 112916 47356 112980 47360
rect 112916 47300 112920 47356
rect 112920 47300 112976 47356
rect 112976 47300 112980 47356
rect 112916 47296 112980 47300
rect 112996 47356 113060 47360
rect 112996 47300 113000 47356
rect 113000 47300 113056 47356
rect 113056 47300 113060 47356
rect 112996 47296 113060 47300
rect 113076 47356 113140 47360
rect 113076 47300 113080 47356
rect 113080 47300 113136 47356
rect 113136 47300 113140 47356
rect 113076 47296 113140 47300
rect 113156 47356 113220 47360
rect 113156 47300 113160 47356
rect 113160 47300 113216 47356
rect 113216 47300 113220 47356
rect 113156 47296 113220 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 113652 46812 113716 46816
rect 113652 46756 113656 46812
rect 113656 46756 113712 46812
rect 113712 46756 113716 46812
rect 113652 46752 113716 46756
rect 113732 46812 113796 46816
rect 113732 46756 113736 46812
rect 113736 46756 113792 46812
rect 113792 46756 113796 46812
rect 113732 46752 113796 46756
rect 113812 46812 113876 46816
rect 113812 46756 113816 46812
rect 113816 46756 113872 46812
rect 113872 46756 113876 46812
rect 113812 46752 113876 46756
rect 113892 46812 113956 46816
rect 113892 46756 113896 46812
rect 113896 46756 113952 46812
rect 113952 46756 113956 46812
rect 113892 46752 113956 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 112916 46268 112980 46272
rect 112916 46212 112920 46268
rect 112920 46212 112976 46268
rect 112976 46212 112980 46268
rect 112916 46208 112980 46212
rect 112996 46268 113060 46272
rect 112996 46212 113000 46268
rect 113000 46212 113056 46268
rect 113056 46212 113060 46268
rect 112996 46208 113060 46212
rect 113076 46268 113140 46272
rect 113076 46212 113080 46268
rect 113080 46212 113136 46268
rect 113136 46212 113140 46268
rect 113076 46208 113140 46212
rect 113156 46268 113220 46272
rect 113156 46212 113160 46268
rect 113160 46212 113216 46268
rect 113216 46212 113220 46268
rect 113156 46208 113220 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 113652 45724 113716 45728
rect 113652 45668 113656 45724
rect 113656 45668 113712 45724
rect 113712 45668 113716 45724
rect 113652 45664 113716 45668
rect 113732 45724 113796 45728
rect 113732 45668 113736 45724
rect 113736 45668 113792 45724
rect 113792 45668 113796 45724
rect 113732 45664 113796 45668
rect 113812 45724 113876 45728
rect 113812 45668 113816 45724
rect 113816 45668 113872 45724
rect 113872 45668 113876 45724
rect 113812 45664 113876 45668
rect 113892 45724 113956 45728
rect 113892 45668 113896 45724
rect 113896 45668 113952 45724
rect 113952 45668 113956 45724
rect 113892 45664 113956 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 112916 45180 112980 45184
rect 112916 45124 112920 45180
rect 112920 45124 112976 45180
rect 112976 45124 112980 45180
rect 112916 45120 112980 45124
rect 112996 45180 113060 45184
rect 112996 45124 113000 45180
rect 113000 45124 113056 45180
rect 113056 45124 113060 45180
rect 112996 45120 113060 45124
rect 113076 45180 113140 45184
rect 113076 45124 113080 45180
rect 113080 45124 113136 45180
rect 113136 45124 113140 45180
rect 113076 45120 113140 45124
rect 113156 45180 113220 45184
rect 113156 45124 113160 45180
rect 113160 45124 113216 45180
rect 113216 45124 113220 45180
rect 113156 45120 113220 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 113652 44636 113716 44640
rect 113652 44580 113656 44636
rect 113656 44580 113712 44636
rect 113712 44580 113716 44636
rect 113652 44576 113716 44580
rect 113732 44636 113796 44640
rect 113732 44580 113736 44636
rect 113736 44580 113792 44636
rect 113792 44580 113796 44636
rect 113732 44576 113796 44580
rect 113812 44636 113876 44640
rect 113812 44580 113816 44636
rect 113816 44580 113872 44636
rect 113872 44580 113876 44636
rect 113812 44576 113876 44580
rect 113892 44636 113956 44640
rect 113892 44580 113896 44636
rect 113896 44580 113952 44636
rect 113952 44580 113956 44636
rect 113892 44576 113956 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 112916 44092 112980 44096
rect 112916 44036 112920 44092
rect 112920 44036 112976 44092
rect 112976 44036 112980 44092
rect 112916 44032 112980 44036
rect 112996 44092 113060 44096
rect 112996 44036 113000 44092
rect 113000 44036 113056 44092
rect 113056 44036 113060 44092
rect 112996 44032 113060 44036
rect 113076 44092 113140 44096
rect 113076 44036 113080 44092
rect 113080 44036 113136 44092
rect 113136 44036 113140 44092
rect 113076 44032 113140 44036
rect 113156 44092 113220 44096
rect 113156 44036 113160 44092
rect 113160 44036 113216 44092
rect 113216 44036 113220 44092
rect 113156 44032 113220 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 113652 43548 113716 43552
rect 113652 43492 113656 43548
rect 113656 43492 113712 43548
rect 113712 43492 113716 43548
rect 113652 43488 113716 43492
rect 113732 43548 113796 43552
rect 113732 43492 113736 43548
rect 113736 43492 113792 43548
rect 113792 43492 113796 43548
rect 113732 43488 113796 43492
rect 113812 43548 113876 43552
rect 113812 43492 113816 43548
rect 113816 43492 113872 43548
rect 113872 43492 113876 43548
rect 113812 43488 113876 43492
rect 113892 43548 113956 43552
rect 113892 43492 113896 43548
rect 113896 43492 113952 43548
rect 113952 43492 113956 43548
rect 113892 43488 113956 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 112916 43004 112980 43008
rect 112916 42948 112920 43004
rect 112920 42948 112976 43004
rect 112976 42948 112980 43004
rect 112916 42944 112980 42948
rect 112996 43004 113060 43008
rect 112996 42948 113000 43004
rect 113000 42948 113056 43004
rect 113056 42948 113060 43004
rect 112996 42944 113060 42948
rect 113076 43004 113140 43008
rect 113076 42948 113080 43004
rect 113080 42948 113136 43004
rect 113136 42948 113140 43004
rect 113076 42944 113140 42948
rect 113156 43004 113220 43008
rect 113156 42948 113160 43004
rect 113160 42948 113216 43004
rect 113216 42948 113220 43004
rect 113156 42944 113220 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 113652 42460 113716 42464
rect 113652 42404 113656 42460
rect 113656 42404 113712 42460
rect 113712 42404 113716 42460
rect 113652 42400 113716 42404
rect 113732 42460 113796 42464
rect 113732 42404 113736 42460
rect 113736 42404 113792 42460
rect 113792 42404 113796 42460
rect 113732 42400 113796 42404
rect 113812 42460 113876 42464
rect 113812 42404 113816 42460
rect 113816 42404 113872 42460
rect 113872 42404 113876 42460
rect 113812 42400 113876 42404
rect 113892 42460 113956 42464
rect 113892 42404 113896 42460
rect 113896 42404 113952 42460
rect 113952 42404 113956 42460
rect 113892 42400 113956 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 112916 41916 112980 41920
rect 112916 41860 112920 41916
rect 112920 41860 112976 41916
rect 112976 41860 112980 41916
rect 112916 41856 112980 41860
rect 112996 41916 113060 41920
rect 112996 41860 113000 41916
rect 113000 41860 113056 41916
rect 113056 41860 113060 41916
rect 112996 41856 113060 41860
rect 113076 41916 113140 41920
rect 113076 41860 113080 41916
rect 113080 41860 113136 41916
rect 113136 41860 113140 41916
rect 113076 41856 113140 41860
rect 113156 41916 113220 41920
rect 113156 41860 113160 41916
rect 113160 41860 113216 41916
rect 113216 41860 113220 41916
rect 113156 41856 113220 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 113652 41372 113716 41376
rect 113652 41316 113656 41372
rect 113656 41316 113712 41372
rect 113712 41316 113716 41372
rect 113652 41312 113716 41316
rect 113732 41372 113796 41376
rect 113732 41316 113736 41372
rect 113736 41316 113792 41372
rect 113792 41316 113796 41372
rect 113732 41312 113796 41316
rect 113812 41372 113876 41376
rect 113812 41316 113816 41372
rect 113816 41316 113872 41372
rect 113872 41316 113876 41372
rect 113812 41312 113876 41316
rect 113892 41372 113956 41376
rect 113892 41316 113896 41372
rect 113896 41316 113952 41372
rect 113952 41316 113956 41372
rect 113892 41312 113956 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 112916 40828 112980 40832
rect 112916 40772 112920 40828
rect 112920 40772 112976 40828
rect 112976 40772 112980 40828
rect 112916 40768 112980 40772
rect 112996 40828 113060 40832
rect 112996 40772 113000 40828
rect 113000 40772 113056 40828
rect 113056 40772 113060 40828
rect 112996 40768 113060 40772
rect 113076 40828 113140 40832
rect 113076 40772 113080 40828
rect 113080 40772 113136 40828
rect 113136 40772 113140 40828
rect 113076 40768 113140 40772
rect 113156 40828 113220 40832
rect 113156 40772 113160 40828
rect 113160 40772 113216 40828
rect 113216 40772 113220 40828
rect 113156 40768 113220 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 113652 40284 113716 40288
rect 113652 40228 113656 40284
rect 113656 40228 113712 40284
rect 113712 40228 113716 40284
rect 113652 40224 113716 40228
rect 113732 40284 113796 40288
rect 113732 40228 113736 40284
rect 113736 40228 113792 40284
rect 113792 40228 113796 40284
rect 113732 40224 113796 40228
rect 113812 40284 113876 40288
rect 113812 40228 113816 40284
rect 113816 40228 113872 40284
rect 113872 40228 113876 40284
rect 113812 40224 113876 40228
rect 113892 40284 113956 40288
rect 113892 40228 113896 40284
rect 113896 40228 113952 40284
rect 113952 40228 113956 40284
rect 113892 40224 113956 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 112916 39740 112980 39744
rect 112916 39684 112920 39740
rect 112920 39684 112976 39740
rect 112976 39684 112980 39740
rect 112916 39680 112980 39684
rect 112996 39740 113060 39744
rect 112996 39684 113000 39740
rect 113000 39684 113056 39740
rect 113056 39684 113060 39740
rect 112996 39680 113060 39684
rect 113076 39740 113140 39744
rect 113076 39684 113080 39740
rect 113080 39684 113136 39740
rect 113136 39684 113140 39740
rect 113076 39680 113140 39684
rect 113156 39740 113220 39744
rect 113156 39684 113160 39740
rect 113160 39684 113216 39740
rect 113216 39684 113220 39740
rect 113156 39680 113220 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 113652 39196 113716 39200
rect 113652 39140 113656 39196
rect 113656 39140 113712 39196
rect 113712 39140 113716 39196
rect 113652 39136 113716 39140
rect 113732 39196 113796 39200
rect 113732 39140 113736 39196
rect 113736 39140 113792 39196
rect 113792 39140 113796 39196
rect 113732 39136 113796 39140
rect 113812 39196 113876 39200
rect 113812 39140 113816 39196
rect 113816 39140 113872 39196
rect 113872 39140 113876 39196
rect 113812 39136 113876 39140
rect 113892 39196 113956 39200
rect 113892 39140 113896 39196
rect 113896 39140 113952 39196
rect 113952 39140 113956 39196
rect 113892 39136 113956 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 112916 38652 112980 38656
rect 112916 38596 112920 38652
rect 112920 38596 112976 38652
rect 112976 38596 112980 38652
rect 112916 38592 112980 38596
rect 112996 38652 113060 38656
rect 112996 38596 113000 38652
rect 113000 38596 113056 38652
rect 113056 38596 113060 38652
rect 112996 38592 113060 38596
rect 113076 38652 113140 38656
rect 113076 38596 113080 38652
rect 113080 38596 113136 38652
rect 113136 38596 113140 38652
rect 113076 38592 113140 38596
rect 113156 38652 113220 38656
rect 113156 38596 113160 38652
rect 113160 38596 113216 38652
rect 113216 38596 113220 38652
rect 113156 38592 113220 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 113652 38108 113716 38112
rect 113652 38052 113656 38108
rect 113656 38052 113712 38108
rect 113712 38052 113716 38108
rect 113652 38048 113716 38052
rect 113732 38108 113796 38112
rect 113732 38052 113736 38108
rect 113736 38052 113792 38108
rect 113792 38052 113796 38108
rect 113732 38048 113796 38052
rect 113812 38108 113876 38112
rect 113812 38052 113816 38108
rect 113816 38052 113872 38108
rect 113872 38052 113876 38108
rect 113812 38048 113876 38052
rect 113892 38108 113956 38112
rect 113892 38052 113896 38108
rect 113896 38052 113952 38108
rect 113952 38052 113956 38108
rect 113892 38048 113956 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 112916 37564 112980 37568
rect 112916 37508 112920 37564
rect 112920 37508 112976 37564
rect 112976 37508 112980 37564
rect 112916 37504 112980 37508
rect 112996 37564 113060 37568
rect 112996 37508 113000 37564
rect 113000 37508 113056 37564
rect 113056 37508 113060 37564
rect 112996 37504 113060 37508
rect 113076 37564 113140 37568
rect 113076 37508 113080 37564
rect 113080 37508 113136 37564
rect 113136 37508 113140 37564
rect 113076 37504 113140 37508
rect 113156 37564 113220 37568
rect 113156 37508 113160 37564
rect 113160 37508 113216 37564
rect 113216 37508 113220 37564
rect 113156 37504 113220 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 113652 37020 113716 37024
rect 113652 36964 113656 37020
rect 113656 36964 113712 37020
rect 113712 36964 113716 37020
rect 113652 36960 113716 36964
rect 113732 37020 113796 37024
rect 113732 36964 113736 37020
rect 113736 36964 113792 37020
rect 113792 36964 113796 37020
rect 113732 36960 113796 36964
rect 113812 37020 113876 37024
rect 113812 36964 113816 37020
rect 113816 36964 113872 37020
rect 113872 36964 113876 37020
rect 113812 36960 113876 36964
rect 113892 37020 113956 37024
rect 113892 36964 113896 37020
rect 113896 36964 113952 37020
rect 113952 36964 113956 37020
rect 113892 36960 113956 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 112916 36476 112980 36480
rect 112916 36420 112920 36476
rect 112920 36420 112976 36476
rect 112976 36420 112980 36476
rect 112916 36416 112980 36420
rect 112996 36476 113060 36480
rect 112996 36420 113000 36476
rect 113000 36420 113056 36476
rect 113056 36420 113060 36476
rect 112996 36416 113060 36420
rect 113076 36476 113140 36480
rect 113076 36420 113080 36476
rect 113080 36420 113136 36476
rect 113136 36420 113140 36476
rect 113076 36416 113140 36420
rect 113156 36476 113220 36480
rect 113156 36420 113160 36476
rect 113160 36420 113216 36476
rect 113216 36420 113220 36476
rect 113156 36416 113220 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 113652 35932 113716 35936
rect 113652 35876 113656 35932
rect 113656 35876 113712 35932
rect 113712 35876 113716 35932
rect 113652 35872 113716 35876
rect 113732 35932 113796 35936
rect 113732 35876 113736 35932
rect 113736 35876 113792 35932
rect 113792 35876 113796 35932
rect 113732 35872 113796 35876
rect 113812 35932 113876 35936
rect 113812 35876 113816 35932
rect 113816 35876 113872 35932
rect 113872 35876 113876 35932
rect 113812 35872 113876 35876
rect 113892 35932 113956 35936
rect 113892 35876 113896 35932
rect 113896 35876 113952 35932
rect 113952 35876 113956 35932
rect 113892 35872 113956 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 112916 35388 112980 35392
rect 112916 35332 112920 35388
rect 112920 35332 112976 35388
rect 112976 35332 112980 35388
rect 112916 35328 112980 35332
rect 112996 35388 113060 35392
rect 112996 35332 113000 35388
rect 113000 35332 113056 35388
rect 113056 35332 113060 35388
rect 112996 35328 113060 35332
rect 113076 35388 113140 35392
rect 113076 35332 113080 35388
rect 113080 35332 113136 35388
rect 113136 35332 113140 35388
rect 113076 35328 113140 35332
rect 113156 35388 113220 35392
rect 113156 35332 113160 35388
rect 113160 35332 113216 35388
rect 113216 35332 113220 35388
rect 113156 35328 113220 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 113652 34844 113716 34848
rect 113652 34788 113656 34844
rect 113656 34788 113712 34844
rect 113712 34788 113716 34844
rect 113652 34784 113716 34788
rect 113732 34844 113796 34848
rect 113732 34788 113736 34844
rect 113736 34788 113792 34844
rect 113792 34788 113796 34844
rect 113732 34784 113796 34788
rect 113812 34844 113876 34848
rect 113812 34788 113816 34844
rect 113816 34788 113872 34844
rect 113872 34788 113876 34844
rect 113812 34784 113876 34788
rect 113892 34844 113956 34848
rect 113892 34788 113896 34844
rect 113896 34788 113952 34844
rect 113952 34788 113956 34844
rect 113892 34784 113956 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 112916 34300 112980 34304
rect 112916 34244 112920 34300
rect 112920 34244 112976 34300
rect 112976 34244 112980 34300
rect 112916 34240 112980 34244
rect 112996 34300 113060 34304
rect 112996 34244 113000 34300
rect 113000 34244 113056 34300
rect 113056 34244 113060 34300
rect 112996 34240 113060 34244
rect 113076 34300 113140 34304
rect 113076 34244 113080 34300
rect 113080 34244 113136 34300
rect 113136 34244 113140 34300
rect 113076 34240 113140 34244
rect 113156 34300 113220 34304
rect 113156 34244 113160 34300
rect 113160 34244 113216 34300
rect 113216 34244 113220 34300
rect 113156 34240 113220 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 113652 33756 113716 33760
rect 113652 33700 113656 33756
rect 113656 33700 113712 33756
rect 113712 33700 113716 33756
rect 113652 33696 113716 33700
rect 113732 33756 113796 33760
rect 113732 33700 113736 33756
rect 113736 33700 113792 33756
rect 113792 33700 113796 33756
rect 113732 33696 113796 33700
rect 113812 33756 113876 33760
rect 113812 33700 113816 33756
rect 113816 33700 113872 33756
rect 113872 33700 113876 33756
rect 113812 33696 113876 33700
rect 113892 33756 113956 33760
rect 113892 33700 113896 33756
rect 113896 33700 113952 33756
rect 113952 33700 113956 33756
rect 113892 33696 113956 33700
rect 109356 33280 109420 33284
rect 109356 33224 109406 33280
rect 109406 33224 109420 33280
rect 109356 33220 109420 33224
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 112916 33212 112980 33216
rect 112916 33156 112920 33212
rect 112920 33156 112976 33212
rect 112976 33156 112980 33212
rect 112916 33152 112980 33156
rect 112996 33212 113060 33216
rect 112996 33156 113000 33212
rect 113000 33156 113056 33212
rect 113056 33156 113060 33212
rect 112996 33152 113060 33156
rect 113076 33212 113140 33216
rect 113076 33156 113080 33212
rect 113080 33156 113136 33212
rect 113136 33156 113140 33212
rect 113076 33152 113140 33156
rect 113156 33212 113220 33216
rect 113156 33156 113160 33212
rect 113160 33156 113216 33212
rect 113216 33156 113220 33212
rect 113156 33152 113220 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 113652 32668 113716 32672
rect 113652 32612 113656 32668
rect 113656 32612 113712 32668
rect 113712 32612 113716 32668
rect 113652 32608 113716 32612
rect 113732 32668 113796 32672
rect 113732 32612 113736 32668
rect 113736 32612 113792 32668
rect 113792 32612 113796 32668
rect 113732 32608 113796 32612
rect 113812 32668 113876 32672
rect 113812 32612 113816 32668
rect 113816 32612 113872 32668
rect 113872 32612 113876 32668
rect 113812 32608 113876 32612
rect 113892 32668 113956 32672
rect 113892 32612 113896 32668
rect 113896 32612 113952 32668
rect 113952 32612 113956 32668
rect 113892 32608 113956 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 112916 32124 112980 32128
rect 112916 32068 112920 32124
rect 112920 32068 112976 32124
rect 112976 32068 112980 32124
rect 112916 32064 112980 32068
rect 112996 32124 113060 32128
rect 112996 32068 113000 32124
rect 113000 32068 113056 32124
rect 113056 32068 113060 32124
rect 112996 32064 113060 32068
rect 113076 32124 113140 32128
rect 113076 32068 113080 32124
rect 113080 32068 113136 32124
rect 113136 32068 113140 32124
rect 113076 32064 113140 32068
rect 113156 32124 113220 32128
rect 113156 32068 113160 32124
rect 113160 32068 113216 32124
rect 113216 32068 113220 32124
rect 113156 32064 113220 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 113652 31580 113716 31584
rect 113652 31524 113656 31580
rect 113656 31524 113712 31580
rect 113712 31524 113716 31580
rect 113652 31520 113716 31524
rect 113732 31580 113796 31584
rect 113732 31524 113736 31580
rect 113736 31524 113792 31580
rect 113792 31524 113796 31580
rect 113732 31520 113796 31524
rect 113812 31580 113876 31584
rect 113812 31524 113816 31580
rect 113816 31524 113872 31580
rect 113872 31524 113876 31580
rect 113812 31520 113876 31524
rect 113892 31580 113956 31584
rect 113892 31524 113896 31580
rect 113896 31524 113952 31580
rect 113952 31524 113956 31580
rect 113892 31520 113956 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 112916 31036 112980 31040
rect 112916 30980 112920 31036
rect 112920 30980 112976 31036
rect 112976 30980 112980 31036
rect 112916 30976 112980 30980
rect 112996 31036 113060 31040
rect 112996 30980 113000 31036
rect 113000 30980 113056 31036
rect 113056 30980 113060 31036
rect 112996 30976 113060 30980
rect 113076 31036 113140 31040
rect 113076 30980 113080 31036
rect 113080 30980 113136 31036
rect 113136 30980 113140 31036
rect 113076 30976 113140 30980
rect 113156 31036 113220 31040
rect 113156 30980 113160 31036
rect 113160 30980 113216 31036
rect 113216 30980 113220 31036
rect 113156 30976 113220 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 113652 30492 113716 30496
rect 113652 30436 113656 30492
rect 113656 30436 113712 30492
rect 113712 30436 113716 30492
rect 113652 30432 113716 30436
rect 113732 30492 113796 30496
rect 113732 30436 113736 30492
rect 113736 30436 113792 30492
rect 113792 30436 113796 30492
rect 113732 30432 113796 30436
rect 113812 30492 113876 30496
rect 113812 30436 113816 30492
rect 113816 30436 113872 30492
rect 113872 30436 113876 30492
rect 113812 30432 113876 30436
rect 113892 30492 113956 30496
rect 113892 30436 113896 30492
rect 113896 30436 113952 30492
rect 113952 30436 113956 30492
rect 113892 30432 113956 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 112916 29948 112980 29952
rect 112916 29892 112920 29948
rect 112920 29892 112976 29948
rect 112976 29892 112980 29948
rect 112916 29888 112980 29892
rect 112996 29948 113060 29952
rect 112996 29892 113000 29948
rect 113000 29892 113056 29948
rect 113056 29892 113060 29948
rect 112996 29888 113060 29892
rect 113076 29948 113140 29952
rect 113076 29892 113080 29948
rect 113080 29892 113136 29948
rect 113136 29892 113140 29948
rect 113076 29888 113140 29892
rect 113156 29948 113220 29952
rect 113156 29892 113160 29948
rect 113160 29892 113216 29948
rect 113216 29892 113220 29948
rect 113156 29888 113220 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 113652 29404 113716 29408
rect 113652 29348 113656 29404
rect 113656 29348 113712 29404
rect 113712 29348 113716 29404
rect 113652 29344 113716 29348
rect 113732 29404 113796 29408
rect 113732 29348 113736 29404
rect 113736 29348 113792 29404
rect 113792 29348 113796 29404
rect 113732 29344 113796 29348
rect 113812 29404 113876 29408
rect 113812 29348 113816 29404
rect 113816 29348 113872 29404
rect 113872 29348 113876 29404
rect 113812 29344 113876 29348
rect 113892 29404 113956 29408
rect 113892 29348 113896 29404
rect 113896 29348 113952 29404
rect 113952 29348 113956 29404
rect 113892 29344 113956 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 112916 28860 112980 28864
rect 112916 28804 112920 28860
rect 112920 28804 112976 28860
rect 112976 28804 112980 28860
rect 112916 28800 112980 28804
rect 112996 28860 113060 28864
rect 112996 28804 113000 28860
rect 113000 28804 113056 28860
rect 113056 28804 113060 28860
rect 112996 28800 113060 28804
rect 113076 28860 113140 28864
rect 113076 28804 113080 28860
rect 113080 28804 113136 28860
rect 113136 28804 113140 28860
rect 113076 28800 113140 28804
rect 113156 28860 113220 28864
rect 113156 28804 113160 28860
rect 113160 28804 113216 28860
rect 113216 28804 113220 28860
rect 113156 28800 113220 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 113652 28316 113716 28320
rect 113652 28260 113656 28316
rect 113656 28260 113712 28316
rect 113712 28260 113716 28316
rect 113652 28256 113716 28260
rect 113732 28316 113796 28320
rect 113732 28260 113736 28316
rect 113736 28260 113792 28316
rect 113792 28260 113796 28316
rect 113732 28256 113796 28260
rect 113812 28316 113876 28320
rect 113812 28260 113816 28316
rect 113816 28260 113872 28316
rect 113872 28260 113876 28316
rect 113812 28256 113876 28260
rect 113892 28316 113956 28320
rect 113892 28260 113896 28316
rect 113896 28260 113952 28316
rect 113952 28260 113956 28316
rect 113892 28256 113956 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 112916 27772 112980 27776
rect 112916 27716 112920 27772
rect 112920 27716 112976 27772
rect 112976 27716 112980 27772
rect 112916 27712 112980 27716
rect 112996 27772 113060 27776
rect 112996 27716 113000 27772
rect 113000 27716 113056 27772
rect 113056 27716 113060 27772
rect 112996 27712 113060 27716
rect 113076 27772 113140 27776
rect 113076 27716 113080 27772
rect 113080 27716 113136 27772
rect 113136 27716 113140 27772
rect 113076 27712 113140 27716
rect 113156 27772 113220 27776
rect 113156 27716 113160 27772
rect 113160 27716 113216 27772
rect 113216 27716 113220 27772
rect 113156 27712 113220 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 113652 27228 113716 27232
rect 113652 27172 113656 27228
rect 113656 27172 113712 27228
rect 113712 27172 113716 27228
rect 113652 27168 113716 27172
rect 113732 27228 113796 27232
rect 113732 27172 113736 27228
rect 113736 27172 113792 27228
rect 113792 27172 113796 27228
rect 113732 27168 113796 27172
rect 113812 27228 113876 27232
rect 113812 27172 113816 27228
rect 113816 27172 113872 27228
rect 113872 27172 113876 27228
rect 113812 27168 113876 27172
rect 113892 27228 113956 27232
rect 113892 27172 113896 27228
rect 113896 27172 113952 27228
rect 113952 27172 113956 27228
rect 113892 27168 113956 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 112916 26684 112980 26688
rect 112916 26628 112920 26684
rect 112920 26628 112976 26684
rect 112976 26628 112980 26684
rect 112916 26624 112980 26628
rect 112996 26684 113060 26688
rect 112996 26628 113000 26684
rect 113000 26628 113056 26684
rect 113056 26628 113060 26684
rect 112996 26624 113060 26628
rect 113076 26684 113140 26688
rect 113076 26628 113080 26684
rect 113080 26628 113136 26684
rect 113136 26628 113140 26684
rect 113076 26624 113140 26628
rect 113156 26684 113220 26688
rect 113156 26628 113160 26684
rect 113160 26628 113216 26684
rect 113216 26628 113220 26684
rect 113156 26624 113220 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 113652 26140 113716 26144
rect 113652 26084 113656 26140
rect 113656 26084 113712 26140
rect 113712 26084 113716 26140
rect 113652 26080 113716 26084
rect 113732 26140 113796 26144
rect 113732 26084 113736 26140
rect 113736 26084 113792 26140
rect 113792 26084 113796 26140
rect 113732 26080 113796 26084
rect 113812 26140 113876 26144
rect 113812 26084 113816 26140
rect 113816 26084 113872 26140
rect 113872 26084 113876 26140
rect 113812 26080 113876 26084
rect 113892 26140 113956 26144
rect 113892 26084 113896 26140
rect 113896 26084 113952 26140
rect 113952 26084 113956 26140
rect 113892 26080 113956 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 112916 25596 112980 25600
rect 112916 25540 112920 25596
rect 112920 25540 112976 25596
rect 112976 25540 112980 25596
rect 112916 25536 112980 25540
rect 112996 25596 113060 25600
rect 112996 25540 113000 25596
rect 113000 25540 113056 25596
rect 113056 25540 113060 25596
rect 112996 25536 113060 25540
rect 113076 25596 113140 25600
rect 113076 25540 113080 25596
rect 113080 25540 113136 25596
rect 113136 25540 113140 25596
rect 113076 25536 113140 25540
rect 113156 25596 113220 25600
rect 113156 25540 113160 25596
rect 113160 25540 113216 25596
rect 113216 25540 113220 25596
rect 113156 25536 113220 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 113652 25052 113716 25056
rect 113652 24996 113656 25052
rect 113656 24996 113712 25052
rect 113712 24996 113716 25052
rect 113652 24992 113716 24996
rect 113732 25052 113796 25056
rect 113732 24996 113736 25052
rect 113736 24996 113792 25052
rect 113792 24996 113796 25052
rect 113732 24992 113796 24996
rect 113812 25052 113876 25056
rect 113812 24996 113816 25052
rect 113816 24996 113872 25052
rect 113872 24996 113876 25052
rect 113812 24992 113876 24996
rect 113892 25052 113956 25056
rect 113892 24996 113896 25052
rect 113896 24996 113952 25052
rect 113952 24996 113956 25052
rect 113892 24992 113956 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 112916 24508 112980 24512
rect 112916 24452 112920 24508
rect 112920 24452 112976 24508
rect 112976 24452 112980 24508
rect 112916 24448 112980 24452
rect 112996 24508 113060 24512
rect 112996 24452 113000 24508
rect 113000 24452 113056 24508
rect 113056 24452 113060 24508
rect 112996 24448 113060 24452
rect 113076 24508 113140 24512
rect 113076 24452 113080 24508
rect 113080 24452 113136 24508
rect 113136 24452 113140 24508
rect 113076 24448 113140 24452
rect 113156 24508 113220 24512
rect 113156 24452 113160 24508
rect 113160 24452 113216 24508
rect 113216 24452 113220 24508
rect 113156 24448 113220 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 113652 23964 113716 23968
rect 113652 23908 113656 23964
rect 113656 23908 113712 23964
rect 113712 23908 113716 23964
rect 113652 23904 113716 23908
rect 113732 23964 113796 23968
rect 113732 23908 113736 23964
rect 113736 23908 113792 23964
rect 113792 23908 113796 23964
rect 113732 23904 113796 23908
rect 113812 23964 113876 23968
rect 113812 23908 113816 23964
rect 113816 23908 113872 23964
rect 113872 23908 113876 23964
rect 113812 23904 113876 23908
rect 113892 23964 113956 23968
rect 113892 23908 113896 23964
rect 113896 23908 113952 23964
rect 113952 23908 113956 23964
rect 113892 23904 113956 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 112916 23420 112980 23424
rect 112916 23364 112920 23420
rect 112920 23364 112976 23420
rect 112976 23364 112980 23420
rect 112916 23360 112980 23364
rect 112996 23420 113060 23424
rect 112996 23364 113000 23420
rect 113000 23364 113056 23420
rect 113056 23364 113060 23420
rect 112996 23360 113060 23364
rect 113076 23420 113140 23424
rect 113076 23364 113080 23420
rect 113080 23364 113136 23420
rect 113136 23364 113140 23420
rect 113076 23360 113140 23364
rect 113156 23420 113220 23424
rect 113156 23364 113160 23420
rect 113160 23364 113216 23420
rect 113216 23364 113220 23420
rect 113156 23360 113220 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 113652 22876 113716 22880
rect 113652 22820 113656 22876
rect 113656 22820 113712 22876
rect 113712 22820 113716 22876
rect 113652 22816 113716 22820
rect 113732 22876 113796 22880
rect 113732 22820 113736 22876
rect 113736 22820 113792 22876
rect 113792 22820 113796 22876
rect 113732 22816 113796 22820
rect 113812 22876 113876 22880
rect 113812 22820 113816 22876
rect 113816 22820 113872 22876
rect 113872 22820 113876 22876
rect 113812 22816 113876 22820
rect 113892 22876 113956 22880
rect 113892 22820 113896 22876
rect 113896 22820 113952 22876
rect 113952 22820 113956 22876
rect 113892 22816 113956 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 112916 22332 112980 22336
rect 112916 22276 112920 22332
rect 112920 22276 112976 22332
rect 112976 22276 112980 22332
rect 112916 22272 112980 22276
rect 112996 22332 113060 22336
rect 112996 22276 113000 22332
rect 113000 22276 113056 22332
rect 113056 22276 113060 22332
rect 112996 22272 113060 22276
rect 113076 22332 113140 22336
rect 113076 22276 113080 22332
rect 113080 22276 113136 22332
rect 113136 22276 113140 22332
rect 113076 22272 113140 22276
rect 113156 22332 113220 22336
rect 113156 22276 113160 22332
rect 113160 22276 113216 22332
rect 113216 22276 113220 22332
rect 113156 22272 113220 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 113652 21788 113716 21792
rect 113652 21732 113656 21788
rect 113656 21732 113712 21788
rect 113712 21732 113716 21788
rect 113652 21728 113716 21732
rect 113732 21788 113796 21792
rect 113732 21732 113736 21788
rect 113736 21732 113792 21788
rect 113792 21732 113796 21788
rect 113732 21728 113796 21732
rect 113812 21788 113876 21792
rect 113812 21732 113816 21788
rect 113816 21732 113872 21788
rect 113872 21732 113876 21788
rect 113812 21728 113876 21732
rect 113892 21788 113956 21792
rect 113892 21732 113896 21788
rect 113896 21732 113952 21788
rect 113952 21732 113956 21788
rect 113892 21728 113956 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 112916 21244 112980 21248
rect 112916 21188 112920 21244
rect 112920 21188 112976 21244
rect 112976 21188 112980 21244
rect 112916 21184 112980 21188
rect 112996 21244 113060 21248
rect 112996 21188 113000 21244
rect 113000 21188 113056 21244
rect 113056 21188 113060 21244
rect 112996 21184 113060 21188
rect 113076 21244 113140 21248
rect 113076 21188 113080 21244
rect 113080 21188 113136 21244
rect 113136 21188 113140 21244
rect 113076 21184 113140 21188
rect 113156 21244 113220 21248
rect 113156 21188 113160 21244
rect 113160 21188 113216 21244
rect 113216 21188 113220 21244
rect 113156 21184 113220 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 113652 20700 113716 20704
rect 113652 20644 113656 20700
rect 113656 20644 113712 20700
rect 113712 20644 113716 20700
rect 113652 20640 113716 20644
rect 113732 20700 113796 20704
rect 113732 20644 113736 20700
rect 113736 20644 113792 20700
rect 113792 20644 113796 20700
rect 113732 20640 113796 20644
rect 113812 20700 113876 20704
rect 113812 20644 113816 20700
rect 113816 20644 113872 20700
rect 113872 20644 113876 20700
rect 113812 20640 113876 20644
rect 113892 20700 113956 20704
rect 113892 20644 113896 20700
rect 113896 20644 113952 20700
rect 113952 20644 113956 20700
rect 113892 20640 113956 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 112916 20156 112980 20160
rect 112916 20100 112920 20156
rect 112920 20100 112976 20156
rect 112976 20100 112980 20156
rect 112916 20096 112980 20100
rect 112996 20156 113060 20160
rect 112996 20100 113000 20156
rect 113000 20100 113056 20156
rect 113056 20100 113060 20156
rect 112996 20096 113060 20100
rect 113076 20156 113140 20160
rect 113076 20100 113080 20156
rect 113080 20100 113136 20156
rect 113136 20100 113140 20156
rect 113076 20096 113140 20100
rect 113156 20156 113220 20160
rect 113156 20100 113160 20156
rect 113160 20100 113216 20156
rect 113216 20100 113220 20156
rect 113156 20096 113220 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 113652 19612 113716 19616
rect 113652 19556 113656 19612
rect 113656 19556 113712 19612
rect 113712 19556 113716 19612
rect 113652 19552 113716 19556
rect 113732 19612 113796 19616
rect 113732 19556 113736 19612
rect 113736 19556 113792 19612
rect 113792 19556 113796 19612
rect 113732 19552 113796 19556
rect 113812 19612 113876 19616
rect 113812 19556 113816 19612
rect 113816 19556 113872 19612
rect 113872 19556 113876 19612
rect 113812 19552 113876 19556
rect 113892 19612 113956 19616
rect 113892 19556 113896 19612
rect 113896 19556 113952 19612
rect 113952 19556 113956 19612
rect 113892 19552 113956 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 112916 19068 112980 19072
rect 112916 19012 112920 19068
rect 112920 19012 112976 19068
rect 112976 19012 112980 19068
rect 112916 19008 112980 19012
rect 112996 19068 113060 19072
rect 112996 19012 113000 19068
rect 113000 19012 113056 19068
rect 113056 19012 113060 19068
rect 112996 19008 113060 19012
rect 113076 19068 113140 19072
rect 113076 19012 113080 19068
rect 113080 19012 113136 19068
rect 113136 19012 113140 19068
rect 113076 19008 113140 19012
rect 113156 19068 113220 19072
rect 113156 19012 113160 19068
rect 113160 19012 113216 19068
rect 113216 19012 113220 19068
rect 113156 19008 113220 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 113652 18524 113716 18528
rect 113652 18468 113656 18524
rect 113656 18468 113712 18524
rect 113712 18468 113716 18524
rect 113652 18464 113716 18468
rect 113732 18524 113796 18528
rect 113732 18468 113736 18524
rect 113736 18468 113792 18524
rect 113792 18468 113796 18524
rect 113732 18464 113796 18468
rect 113812 18524 113876 18528
rect 113812 18468 113816 18524
rect 113816 18468 113872 18524
rect 113872 18468 113876 18524
rect 113812 18464 113876 18468
rect 113892 18524 113956 18528
rect 113892 18468 113896 18524
rect 113896 18468 113952 18524
rect 113952 18468 113956 18524
rect 113892 18464 113956 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 112916 17980 112980 17984
rect 112916 17924 112920 17980
rect 112920 17924 112976 17980
rect 112976 17924 112980 17980
rect 112916 17920 112980 17924
rect 112996 17980 113060 17984
rect 112996 17924 113000 17980
rect 113000 17924 113056 17980
rect 113056 17924 113060 17980
rect 112996 17920 113060 17924
rect 113076 17980 113140 17984
rect 113076 17924 113080 17980
rect 113080 17924 113136 17980
rect 113136 17924 113140 17980
rect 113076 17920 113140 17924
rect 113156 17980 113220 17984
rect 113156 17924 113160 17980
rect 113160 17924 113216 17980
rect 113216 17924 113220 17980
rect 113156 17920 113220 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 113652 17436 113716 17440
rect 113652 17380 113656 17436
rect 113656 17380 113712 17436
rect 113712 17380 113716 17436
rect 113652 17376 113716 17380
rect 113732 17436 113796 17440
rect 113732 17380 113736 17436
rect 113736 17380 113792 17436
rect 113792 17380 113796 17436
rect 113732 17376 113796 17380
rect 113812 17436 113876 17440
rect 113812 17380 113816 17436
rect 113816 17380 113872 17436
rect 113872 17380 113876 17436
rect 113812 17376 113876 17380
rect 113892 17436 113956 17440
rect 113892 17380 113896 17436
rect 113896 17380 113952 17436
rect 113952 17380 113956 17436
rect 113892 17376 113956 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 112916 16892 112980 16896
rect 112916 16836 112920 16892
rect 112920 16836 112976 16892
rect 112976 16836 112980 16892
rect 112916 16832 112980 16836
rect 112996 16892 113060 16896
rect 112996 16836 113000 16892
rect 113000 16836 113056 16892
rect 113056 16836 113060 16892
rect 112996 16832 113060 16836
rect 113076 16892 113140 16896
rect 113076 16836 113080 16892
rect 113080 16836 113136 16892
rect 113136 16836 113140 16892
rect 113076 16832 113140 16836
rect 113156 16892 113220 16896
rect 113156 16836 113160 16892
rect 113160 16836 113216 16892
rect 113216 16836 113220 16892
rect 113156 16832 113220 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 113652 16348 113716 16352
rect 113652 16292 113656 16348
rect 113656 16292 113712 16348
rect 113712 16292 113716 16348
rect 113652 16288 113716 16292
rect 113732 16348 113796 16352
rect 113732 16292 113736 16348
rect 113736 16292 113792 16348
rect 113792 16292 113796 16348
rect 113732 16288 113796 16292
rect 113812 16348 113876 16352
rect 113812 16292 113816 16348
rect 113816 16292 113872 16348
rect 113872 16292 113876 16348
rect 113812 16288 113876 16292
rect 113892 16348 113956 16352
rect 113892 16292 113896 16348
rect 113896 16292 113952 16348
rect 113952 16292 113956 16348
rect 113892 16288 113956 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 112916 15804 112980 15808
rect 112916 15748 112920 15804
rect 112920 15748 112976 15804
rect 112976 15748 112980 15804
rect 112916 15744 112980 15748
rect 112996 15804 113060 15808
rect 112996 15748 113000 15804
rect 113000 15748 113056 15804
rect 113056 15748 113060 15804
rect 112996 15744 113060 15748
rect 113076 15804 113140 15808
rect 113076 15748 113080 15804
rect 113080 15748 113136 15804
rect 113136 15748 113140 15804
rect 113076 15744 113140 15748
rect 113156 15804 113220 15808
rect 113156 15748 113160 15804
rect 113160 15748 113216 15804
rect 113216 15748 113220 15804
rect 113156 15744 113220 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 113652 15260 113716 15264
rect 113652 15204 113656 15260
rect 113656 15204 113712 15260
rect 113712 15204 113716 15260
rect 113652 15200 113716 15204
rect 113732 15260 113796 15264
rect 113732 15204 113736 15260
rect 113736 15204 113792 15260
rect 113792 15204 113796 15260
rect 113732 15200 113796 15204
rect 113812 15260 113876 15264
rect 113812 15204 113816 15260
rect 113816 15204 113872 15260
rect 113872 15204 113876 15260
rect 113812 15200 113876 15204
rect 113892 15260 113956 15264
rect 113892 15204 113896 15260
rect 113896 15204 113952 15260
rect 113952 15204 113956 15260
rect 113892 15200 113956 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 112916 14716 112980 14720
rect 112916 14660 112920 14716
rect 112920 14660 112976 14716
rect 112976 14660 112980 14716
rect 112916 14656 112980 14660
rect 112996 14716 113060 14720
rect 112996 14660 113000 14716
rect 113000 14660 113056 14716
rect 113056 14660 113060 14716
rect 112996 14656 113060 14660
rect 113076 14716 113140 14720
rect 113076 14660 113080 14716
rect 113080 14660 113136 14716
rect 113136 14660 113140 14716
rect 113076 14656 113140 14660
rect 113156 14716 113220 14720
rect 113156 14660 113160 14716
rect 113160 14660 113216 14716
rect 113216 14660 113220 14716
rect 113156 14656 113220 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 113652 14172 113716 14176
rect 113652 14116 113656 14172
rect 113656 14116 113712 14172
rect 113712 14116 113716 14172
rect 113652 14112 113716 14116
rect 113732 14172 113796 14176
rect 113732 14116 113736 14172
rect 113736 14116 113792 14172
rect 113792 14116 113796 14172
rect 113732 14112 113796 14116
rect 113812 14172 113876 14176
rect 113812 14116 113816 14172
rect 113816 14116 113872 14172
rect 113872 14116 113876 14172
rect 113812 14112 113876 14116
rect 113892 14172 113956 14176
rect 113892 14116 113896 14172
rect 113896 14116 113952 14172
rect 113952 14116 113956 14172
rect 113892 14112 113956 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 112916 13628 112980 13632
rect 112916 13572 112920 13628
rect 112920 13572 112976 13628
rect 112976 13572 112980 13628
rect 112916 13568 112980 13572
rect 112996 13628 113060 13632
rect 112996 13572 113000 13628
rect 113000 13572 113056 13628
rect 113056 13572 113060 13628
rect 112996 13568 113060 13572
rect 113076 13628 113140 13632
rect 113076 13572 113080 13628
rect 113080 13572 113136 13628
rect 113136 13572 113140 13628
rect 113076 13568 113140 13572
rect 113156 13628 113220 13632
rect 113156 13572 113160 13628
rect 113160 13572 113216 13628
rect 113216 13572 113220 13628
rect 113156 13568 113220 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 113652 13084 113716 13088
rect 113652 13028 113656 13084
rect 113656 13028 113712 13084
rect 113712 13028 113716 13084
rect 113652 13024 113716 13028
rect 113732 13084 113796 13088
rect 113732 13028 113736 13084
rect 113736 13028 113792 13084
rect 113792 13028 113796 13084
rect 113732 13024 113796 13028
rect 113812 13084 113876 13088
rect 113812 13028 113816 13084
rect 113816 13028 113872 13084
rect 113872 13028 113876 13084
rect 113812 13024 113876 13028
rect 113892 13084 113956 13088
rect 113892 13028 113896 13084
rect 113896 13028 113952 13084
rect 113952 13028 113956 13084
rect 113892 13024 113956 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 112916 12540 112980 12544
rect 112916 12484 112920 12540
rect 112920 12484 112976 12540
rect 112976 12484 112980 12540
rect 112916 12480 112980 12484
rect 112996 12540 113060 12544
rect 112996 12484 113000 12540
rect 113000 12484 113056 12540
rect 113056 12484 113060 12540
rect 112996 12480 113060 12484
rect 113076 12540 113140 12544
rect 113076 12484 113080 12540
rect 113080 12484 113136 12540
rect 113136 12484 113140 12540
rect 113076 12480 113140 12484
rect 113156 12540 113220 12544
rect 113156 12484 113160 12540
rect 113160 12484 113216 12540
rect 113216 12484 113220 12540
rect 113156 12480 113220 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 113652 11996 113716 12000
rect 113652 11940 113656 11996
rect 113656 11940 113712 11996
rect 113712 11940 113716 11996
rect 113652 11936 113716 11940
rect 113732 11996 113796 12000
rect 113732 11940 113736 11996
rect 113736 11940 113792 11996
rect 113792 11940 113796 11996
rect 113732 11936 113796 11940
rect 113812 11996 113876 12000
rect 113812 11940 113816 11996
rect 113816 11940 113872 11996
rect 113872 11940 113876 11996
rect 113812 11936 113876 11940
rect 113892 11996 113956 12000
rect 113892 11940 113896 11996
rect 113896 11940 113952 11996
rect 113952 11940 113956 11996
rect 113892 11936 113956 11940
rect 109356 11868 109420 11932
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 112916 11452 112980 11456
rect 112916 11396 112920 11452
rect 112920 11396 112976 11452
rect 112976 11396 112980 11452
rect 112916 11392 112980 11396
rect 112996 11452 113060 11456
rect 112996 11396 113000 11452
rect 113000 11396 113056 11452
rect 113056 11396 113060 11452
rect 112996 11392 113060 11396
rect 113076 11452 113140 11456
rect 113076 11396 113080 11452
rect 113080 11396 113136 11452
rect 113136 11396 113140 11452
rect 113076 11392 113140 11396
rect 113156 11452 113220 11456
rect 113156 11396 113160 11452
rect 113160 11396 113216 11452
rect 113216 11396 113220 11452
rect 113156 11392 113220 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 113652 10908 113716 10912
rect 113652 10852 113656 10908
rect 113656 10852 113712 10908
rect 113712 10852 113716 10908
rect 113652 10848 113716 10852
rect 113732 10908 113796 10912
rect 113732 10852 113736 10908
rect 113736 10852 113792 10908
rect 113792 10852 113796 10908
rect 113732 10848 113796 10852
rect 113812 10908 113876 10912
rect 113812 10852 113816 10908
rect 113816 10852 113872 10908
rect 113872 10852 113876 10908
rect 113812 10848 113876 10852
rect 113892 10908 113956 10912
rect 113892 10852 113896 10908
rect 113896 10852 113952 10908
rect 113952 10852 113956 10908
rect 113892 10848 113956 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 112916 10364 112980 10368
rect 112916 10308 112920 10364
rect 112920 10308 112976 10364
rect 112976 10308 112980 10364
rect 112916 10304 112980 10308
rect 112996 10364 113060 10368
rect 112996 10308 113000 10364
rect 113000 10308 113056 10364
rect 113056 10308 113060 10364
rect 112996 10304 113060 10308
rect 113076 10364 113140 10368
rect 113076 10308 113080 10364
rect 113080 10308 113136 10364
rect 113136 10308 113140 10364
rect 113076 10304 113140 10308
rect 113156 10364 113220 10368
rect 113156 10308 113160 10364
rect 113160 10308 113216 10364
rect 113216 10308 113220 10364
rect 113156 10304 113220 10308
rect 93348 9964 93412 10028
rect 15854 9888 15918 9892
rect 15854 9832 15898 9888
rect 15898 9832 15918 9888
rect 15854 9828 15918 9832
rect 92694 9888 92758 9892
rect 92694 9832 92754 9888
rect 92754 9832 92758 9888
rect 92694 9828 92758 9832
rect 92966 9828 93030 9892
rect 93102 9828 93166 9892
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 113652 9820 113716 9824
rect 113652 9764 113656 9820
rect 113656 9764 113712 9820
rect 113712 9764 113716 9820
rect 113652 9760 113716 9764
rect 113732 9820 113796 9824
rect 113732 9764 113736 9820
rect 113736 9764 113792 9820
rect 113792 9764 113796 9820
rect 113732 9760 113796 9764
rect 113812 9820 113876 9824
rect 113812 9764 113816 9820
rect 113816 9764 113872 9820
rect 113872 9764 113876 9820
rect 113812 9760 113876 9764
rect 113892 9820 113956 9824
rect 113892 9764 113896 9820
rect 113896 9764 113952 9820
rect 113952 9764 113956 9820
rect 113892 9760 113956 9764
rect 26734 9692 26798 9756
rect 27822 9752 27886 9756
rect 27822 9696 27858 9752
rect 27858 9696 27886 9752
rect 27822 9692 27886 9696
rect 29182 9692 29246 9756
rect 30134 9752 30198 9756
rect 30134 9696 30194 9752
rect 30194 9696 30198 9752
rect 30134 9692 30198 9696
rect 51350 9692 51414 9756
rect 52438 9752 52502 9756
rect 52438 9696 52458 9752
rect 52458 9696 52502 9752
rect 52438 9692 52502 9696
rect 53526 9752 53590 9756
rect 53526 9696 53562 9752
rect 53562 9696 53590 9752
rect 53526 9692 53590 9696
rect 54886 9692 54950 9756
rect 55974 9692 56038 9756
rect 57062 9692 57126 9756
rect 58286 9752 58350 9756
rect 58286 9696 58310 9752
rect 58310 9696 58350 9752
rect 58286 9692 58350 9696
rect 59374 9692 59438 9756
rect 60780 9752 60844 9756
rect 60780 9696 60830 9752
rect 60830 9696 60844 9752
rect 60780 9692 60844 9696
rect 67670 9752 67734 9756
rect 67670 9696 67730 9752
rect 67730 9696 67734 9752
rect 67670 9692 67734 9696
rect 92830 9692 92894 9756
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 112916 9276 112980 9280
rect 112916 9220 112920 9276
rect 112920 9220 112976 9276
rect 112976 9220 112980 9276
rect 112916 9216 112980 9220
rect 112996 9276 113060 9280
rect 112996 9220 113000 9276
rect 113000 9220 113056 9276
rect 113056 9220 113060 9276
rect 112996 9216 113060 9220
rect 113076 9276 113140 9280
rect 113076 9220 113080 9276
rect 113080 9220 113136 9276
rect 113136 9220 113140 9276
rect 113076 9216 113140 9220
rect 113156 9276 113220 9280
rect 113156 9220 113160 9276
rect 113160 9220 113216 9276
rect 113216 9220 113220 9276
rect 113156 9216 113220 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 113652 8732 113716 8736
rect 113652 8676 113656 8732
rect 113656 8676 113712 8732
rect 113712 8676 113716 8732
rect 113652 8672 113716 8676
rect 113732 8732 113796 8736
rect 113732 8676 113736 8732
rect 113736 8676 113792 8732
rect 113792 8676 113796 8732
rect 113732 8672 113796 8676
rect 113812 8732 113876 8736
rect 113812 8676 113816 8732
rect 113816 8676 113872 8732
rect 113872 8676 113876 8732
rect 113812 8672 113876 8676
rect 113892 8732 113956 8736
rect 113892 8676 113896 8732
rect 113896 8676 113952 8732
rect 113952 8676 113956 8732
rect 113892 8672 113956 8676
rect 25452 8196 25516 8260
rect 31340 8196 31404 8260
rect 32628 8196 32692 8260
rect 33732 8256 33796 8260
rect 33732 8200 33782 8256
rect 33782 8200 33796 8256
rect 33732 8196 33796 8200
rect 35020 8196 35084 8260
rect 36124 8256 36188 8260
rect 36124 8200 36174 8256
rect 36174 8200 36188 8256
rect 36124 8196 36188 8200
rect 37228 8196 37292 8260
rect 38332 8256 38396 8260
rect 38332 8200 38346 8256
rect 38346 8200 38396 8256
rect 38332 8196 38396 8200
rect 40724 8196 40788 8260
rect 41828 8196 41892 8260
rect 43116 8196 43180 8260
rect 44220 8196 44284 8260
rect 46612 8256 46676 8260
rect 46612 8200 46662 8256
rect 46662 8200 46676 8256
rect 46612 8196 46676 8200
rect 47716 8256 47780 8260
rect 47716 8200 47766 8256
rect 47766 8200 47780 8256
rect 47716 8196 47780 8200
rect 49004 8256 49068 8260
rect 49004 8200 49054 8256
rect 49054 8200 49068 8256
rect 49004 8196 49068 8200
rect 50292 8256 50356 8260
rect 50292 8200 50342 8256
rect 50342 8200 50356 8256
rect 50292 8196 50356 8200
rect 61884 8256 61948 8260
rect 61884 8200 61934 8256
rect 61934 8200 61948 8256
rect 61884 8196 61948 8200
rect 62988 8196 63052 8260
rect 64092 8256 64156 8260
rect 64092 8200 64106 8256
rect 64106 8200 64156 8256
rect 64092 8196 64156 8200
rect 65196 8196 65260 8260
rect 66668 8256 66732 8260
rect 66668 8200 66718 8256
rect 66718 8200 66732 8256
rect 66668 8196 66732 8200
rect 93348 8196 93412 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 112916 8188 112980 8192
rect 112916 8132 112920 8188
rect 112920 8132 112976 8188
rect 112976 8132 112980 8188
rect 112916 8128 112980 8132
rect 112996 8188 113060 8192
rect 112996 8132 113000 8188
rect 113000 8132 113056 8188
rect 113056 8132 113060 8188
rect 112996 8128 113060 8132
rect 113076 8188 113140 8192
rect 113076 8132 113080 8188
rect 113080 8132 113136 8188
rect 113136 8132 113140 8188
rect 113076 8128 113140 8132
rect 113156 8188 113220 8192
rect 113156 8132 113160 8188
rect 113160 8132 113216 8188
rect 113216 8132 113220 8188
rect 113156 8128 113220 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 66316 7644 66380 7648
rect 66316 7588 66320 7644
rect 66320 7588 66376 7644
rect 66376 7588 66380 7644
rect 66316 7584 66380 7588
rect 66396 7644 66460 7648
rect 66396 7588 66400 7644
rect 66400 7588 66456 7644
rect 66456 7588 66460 7644
rect 66396 7584 66460 7588
rect 66476 7644 66540 7648
rect 66476 7588 66480 7644
rect 66480 7588 66536 7644
rect 66536 7588 66540 7644
rect 66476 7584 66540 7588
rect 66556 7644 66620 7648
rect 66556 7588 66560 7644
rect 66560 7588 66616 7644
rect 66616 7588 66620 7644
rect 66556 7584 66620 7588
rect 97036 7644 97100 7648
rect 97036 7588 97040 7644
rect 97040 7588 97096 7644
rect 97096 7588 97100 7644
rect 97036 7584 97100 7588
rect 97116 7644 97180 7648
rect 97116 7588 97120 7644
rect 97120 7588 97176 7644
rect 97176 7588 97180 7644
rect 97116 7584 97180 7588
rect 97196 7644 97260 7648
rect 97196 7588 97200 7644
rect 97200 7588 97256 7644
rect 97256 7588 97260 7644
rect 97196 7584 97260 7588
rect 97276 7644 97340 7648
rect 97276 7588 97280 7644
rect 97280 7588 97336 7644
rect 97336 7588 97340 7644
rect 97276 7584 97340 7588
rect 113652 7644 113716 7648
rect 113652 7588 113656 7644
rect 113656 7588 113712 7644
rect 113712 7588 113716 7644
rect 113652 7584 113716 7588
rect 113732 7644 113796 7648
rect 113732 7588 113736 7644
rect 113736 7588 113792 7644
rect 113792 7588 113796 7644
rect 113732 7584 113796 7588
rect 113812 7644 113876 7648
rect 113812 7588 113816 7644
rect 113816 7588 113872 7644
rect 113872 7588 113876 7644
rect 113812 7584 113876 7588
rect 113892 7644 113956 7648
rect 113892 7588 113896 7644
rect 113896 7588 113952 7644
rect 113952 7588 113956 7644
rect 113892 7584 113956 7588
rect 45508 7108 45572 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 112916 7100 112980 7104
rect 112916 7044 112920 7100
rect 112920 7044 112976 7100
rect 112976 7044 112980 7100
rect 112916 7040 112980 7044
rect 112996 7100 113060 7104
rect 112996 7044 113000 7100
rect 113000 7044 113056 7100
rect 113056 7044 113060 7100
rect 112996 7040 113060 7044
rect 113076 7100 113140 7104
rect 113076 7044 113080 7100
rect 113080 7044 113136 7100
rect 113136 7044 113140 7100
rect 113076 7040 113140 7044
rect 113156 7100 113220 7104
rect 113156 7044 113160 7100
rect 113160 7044 113216 7100
rect 113216 7044 113220 7100
rect 113156 7040 113220 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 66316 6556 66380 6560
rect 66316 6500 66320 6556
rect 66320 6500 66376 6556
rect 66376 6500 66380 6556
rect 66316 6496 66380 6500
rect 66396 6556 66460 6560
rect 66396 6500 66400 6556
rect 66400 6500 66456 6556
rect 66456 6500 66460 6556
rect 66396 6496 66460 6500
rect 66476 6556 66540 6560
rect 66476 6500 66480 6556
rect 66480 6500 66536 6556
rect 66536 6500 66540 6556
rect 66476 6496 66540 6500
rect 66556 6556 66620 6560
rect 66556 6500 66560 6556
rect 66560 6500 66616 6556
rect 66616 6500 66620 6556
rect 66556 6496 66620 6500
rect 97036 6556 97100 6560
rect 97036 6500 97040 6556
rect 97040 6500 97096 6556
rect 97096 6500 97100 6556
rect 97036 6496 97100 6500
rect 97116 6556 97180 6560
rect 97116 6500 97120 6556
rect 97120 6500 97176 6556
rect 97176 6500 97180 6556
rect 97116 6496 97180 6500
rect 97196 6556 97260 6560
rect 97196 6500 97200 6556
rect 97200 6500 97256 6556
rect 97256 6500 97260 6556
rect 97196 6496 97260 6500
rect 97276 6556 97340 6560
rect 97276 6500 97280 6556
rect 97280 6500 97336 6556
rect 97336 6500 97340 6556
rect 97276 6496 97340 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 66316 5468 66380 5472
rect 66316 5412 66320 5468
rect 66320 5412 66376 5468
rect 66376 5412 66380 5468
rect 66316 5408 66380 5412
rect 66396 5468 66460 5472
rect 66396 5412 66400 5468
rect 66400 5412 66456 5468
rect 66456 5412 66460 5468
rect 66396 5408 66460 5412
rect 66476 5468 66540 5472
rect 66476 5412 66480 5468
rect 66480 5412 66536 5468
rect 66536 5412 66540 5468
rect 66476 5408 66540 5412
rect 66556 5468 66620 5472
rect 66556 5412 66560 5468
rect 66560 5412 66616 5468
rect 66616 5412 66620 5468
rect 66556 5408 66620 5412
rect 97036 5468 97100 5472
rect 97036 5412 97040 5468
rect 97040 5412 97096 5468
rect 97096 5412 97100 5468
rect 97036 5408 97100 5412
rect 97116 5468 97180 5472
rect 97116 5412 97120 5468
rect 97120 5412 97176 5468
rect 97176 5412 97180 5468
rect 97116 5408 97180 5412
rect 97196 5468 97260 5472
rect 97196 5412 97200 5468
rect 97200 5412 97256 5468
rect 97256 5412 97260 5468
rect 97196 5408 97260 5412
rect 97276 5468 97340 5472
rect 97276 5412 97280 5468
rect 97280 5412 97336 5468
rect 97336 5412 97340 5468
rect 97276 5408 97340 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 66316 4380 66380 4384
rect 66316 4324 66320 4380
rect 66320 4324 66376 4380
rect 66376 4324 66380 4380
rect 66316 4320 66380 4324
rect 66396 4380 66460 4384
rect 66396 4324 66400 4380
rect 66400 4324 66456 4380
rect 66456 4324 66460 4380
rect 66396 4320 66460 4324
rect 66476 4380 66540 4384
rect 66476 4324 66480 4380
rect 66480 4324 66536 4380
rect 66536 4324 66540 4380
rect 66476 4320 66540 4324
rect 66556 4380 66620 4384
rect 66556 4324 66560 4380
rect 66560 4324 66616 4380
rect 66616 4324 66620 4380
rect 66556 4320 66620 4324
rect 97036 4380 97100 4384
rect 97036 4324 97040 4380
rect 97040 4324 97096 4380
rect 97096 4324 97100 4380
rect 97036 4320 97100 4324
rect 97116 4380 97180 4384
rect 97116 4324 97120 4380
rect 97120 4324 97176 4380
rect 97176 4324 97180 4380
rect 97116 4320 97180 4324
rect 97196 4380 97260 4384
rect 97196 4324 97200 4380
rect 97200 4324 97256 4380
rect 97256 4324 97260 4380
rect 97196 4320 97260 4324
rect 97276 4380 97340 4384
rect 97276 4324 97280 4380
rect 97280 4324 97336 4380
rect 97336 4324 97340 4380
rect 97276 4320 97340 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 66316 3292 66380 3296
rect 66316 3236 66320 3292
rect 66320 3236 66376 3292
rect 66376 3236 66380 3292
rect 66316 3232 66380 3236
rect 66396 3292 66460 3296
rect 66396 3236 66400 3292
rect 66400 3236 66456 3292
rect 66456 3236 66460 3292
rect 66396 3232 66460 3236
rect 66476 3292 66540 3296
rect 66476 3236 66480 3292
rect 66480 3236 66536 3292
rect 66536 3236 66540 3292
rect 66476 3232 66540 3236
rect 66556 3292 66620 3296
rect 66556 3236 66560 3292
rect 66560 3236 66616 3292
rect 66616 3236 66620 3292
rect 66556 3232 66620 3236
rect 97036 3292 97100 3296
rect 97036 3236 97040 3292
rect 97040 3236 97096 3292
rect 97096 3236 97100 3292
rect 97036 3232 97100 3236
rect 97116 3292 97180 3296
rect 97116 3236 97120 3292
rect 97120 3236 97176 3292
rect 97176 3236 97180 3292
rect 97116 3232 97180 3236
rect 97196 3292 97260 3296
rect 97196 3236 97200 3292
rect 97200 3236 97256 3292
rect 97256 3236 97260 3292
rect 97196 3232 97260 3236
rect 97276 3292 97340 3296
rect 97276 3236 97280 3292
rect 97280 3236 97336 3292
rect 97336 3236 97340 3292
rect 97276 3232 97340 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 39620 2620 39684 2684
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
rect 66316 2204 66380 2208
rect 66316 2148 66320 2204
rect 66320 2148 66376 2204
rect 66376 2148 66380 2204
rect 66316 2144 66380 2148
rect 66396 2204 66460 2208
rect 66396 2148 66400 2204
rect 66400 2148 66456 2204
rect 66456 2148 66460 2204
rect 66396 2144 66460 2148
rect 66476 2204 66540 2208
rect 66476 2148 66480 2204
rect 66480 2148 66536 2204
rect 66536 2148 66540 2204
rect 66476 2144 66540 2148
rect 66556 2204 66620 2208
rect 66556 2148 66560 2204
rect 66560 2148 66616 2204
rect 66616 2148 66620 2204
rect 66556 2144 66620 2148
rect 97036 2204 97100 2208
rect 97036 2148 97040 2204
rect 97040 2148 97096 2204
rect 97096 2148 97100 2204
rect 97036 2144 97100 2148
rect 97116 2204 97180 2208
rect 97116 2148 97120 2204
rect 97120 2148 97176 2204
rect 97176 2148 97180 2204
rect 97116 2144 97180 2148
rect 97196 2204 97260 2208
rect 97196 2148 97200 2204
rect 97200 2148 97256 2204
rect 97256 2148 97260 2204
rect 97196 2144 97260 2148
rect 97276 2204 97340 2208
rect 97276 2148 97280 2204
rect 97280 2148 97336 2204
rect 97336 2148 97340 2204
rect 97276 2144 97340 2148
<< metal4 >>
rect 4208 97408 4528 97424
rect 4208 97344 4216 97408
rect 4280 97344 4296 97408
rect 4360 97344 4376 97408
rect 4440 97344 4456 97408
rect 4520 97344 4528 97408
rect 4208 96320 4528 97344
rect 4208 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4528 96320
rect 4208 95232 4528 96256
rect 4208 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4528 95232
rect 4208 94298 4528 95168
rect 4208 94144 4250 94298
rect 4486 94144 4528 94298
rect 4208 94080 4216 94144
rect 4520 94080 4528 94144
rect 4208 94062 4250 94080
rect 4486 94062 4528 94080
rect 4208 93056 4528 94062
rect 4208 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4528 93056
rect 4208 91968 4528 92992
rect 4208 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4528 91968
rect 4208 90880 4528 91904
rect 4208 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4528 90880
rect 4208 89792 4528 90816
rect 4208 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4528 89792
rect 4208 88704 4528 89728
rect 4208 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4528 88704
rect 4208 87616 4528 88640
rect 4208 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4528 87616
rect 4208 86528 4528 87552
rect 4208 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4528 86528
rect 4208 85440 4528 86464
rect 4208 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4528 85440
rect 4208 84352 4528 85376
rect 4208 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4528 84352
rect 4208 83264 4528 84288
rect 4208 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4528 83264
rect 4208 82176 4528 83200
rect 4208 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4528 82176
rect 4208 81088 4528 82112
rect 4208 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4528 81088
rect 4208 80000 4528 81024
rect 4208 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4528 80000
rect 4208 78912 4528 79936
rect 4208 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4528 78912
rect 4208 77824 4528 78848
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 76736 4528 77760
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 75648 4528 76672
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 4208 74560 4528 75584
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 73472 4528 74496
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66896 4296 66944
rect 4360 66896 4376 66944
rect 4440 66896 4456 66944
rect 4520 66880 4528 66944
rect 4208 66660 4250 66880
rect 4486 66660 4528 66880
rect 4208 65856 4528 66660
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 96864 5188 97424
rect 4868 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5188 96864
rect 4868 95776 5188 96800
rect 4868 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5188 95776
rect 4868 94978 5188 95712
rect 4868 94742 4910 94978
rect 5146 94742 5188 94978
rect 4868 94688 5188 94742
rect 4868 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5188 94688
rect 4868 93600 5188 94624
rect 4868 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5188 93600
rect 4868 92512 5188 93536
rect 4868 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5188 92512
rect 4868 91424 5188 92448
rect 34928 97408 35248 97424
rect 34928 97344 34936 97408
rect 35000 97344 35016 97408
rect 35080 97344 35096 97408
rect 35160 97344 35176 97408
rect 35240 97344 35248 97408
rect 34928 96320 35248 97344
rect 34928 96256 34936 96320
rect 35000 96256 35016 96320
rect 35080 96256 35096 96320
rect 35160 96256 35176 96320
rect 35240 96256 35248 96320
rect 34928 95232 35248 96256
rect 34928 95168 34936 95232
rect 35000 95168 35016 95232
rect 35080 95168 35096 95232
rect 35160 95168 35176 95232
rect 35240 95168 35248 95232
rect 34928 94298 35248 95168
rect 34928 94144 34970 94298
rect 35206 94144 35248 94298
rect 34928 94080 34936 94144
rect 35240 94080 35248 94144
rect 34928 94062 34970 94080
rect 35206 94062 35248 94080
rect 34928 93056 35248 94062
rect 34928 92992 34936 93056
rect 35000 92992 35016 93056
rect 35080 92992 35096 93056
rect 35160 92992 35176 93056
rect 35240 92992 35248 93056
rect 34928 91968 35248 92992
rect 34928 91904 34936 91968
rect 35000 91904 35016 91968
rect 35080 91904 35096 91968
rect 35160 91904 35176 91968
rect 35240 91904 35248 91968
rect 34928 91436 35248 91904
rect 35588 96864 35908 97424
rect 35588 96800 35596 96864
rect 35660 96800 35676 96864
rect 35740 96800 35756 96864
rect 35820 96800 35836 96864
rect 35900 96800 35908 96864
rect 35588 95776 35908 96800
rect 35588 95712 35596 95776
rect 35660 95712 35676 95776
rect 35740 95712 35756 95776
rect 35820 95712 35836 95776
rect 35900 95712 35908 95776
rect 35588 94978 35908 95712
rect 35588 94742 35630 94978
rect 35866 94742 35908 94978
rect 35588 94688 35908 94742
rect 35588 94624 35596 94688
rect 35660 94624 35676 94688
rect 35740 94624 35756 94688
rect 35820 94624 35836 94688
rect 35900 94624 35908 94688
rect 35588 93600 35908 94624
rect 65648 97408 65968 97424
rect 65648 97344 65656 97408
rect 65720 97344 65736 97408
rect 65800 97344 65816 97408
rect 65880 97344 65896 97408
rect 65960 97344 65968 97408
rect 65648 96320 65968 97344
rect 65648 96256 65656 96320
rect 65720 96256 65736 96320
rect 65800 96256 65816 96320
rect 65880 96256 65896 96320
rect 65960 96256 65968 96320
rect 65648 95232 65968 96256
rect 65648 95168 65656 95232
rect 65720 95168 65736 95232
rect 65800 95168 65816 95232
rect 65880 95168 65896 95232
rect 65960 95168 65968 95232
rect 65648 94298 65968 95168
rect 65648 94144 65690 94298
rect 65926 94144 65968 94298
rect 65648 94080 65656 94144
rect 65960 94080 65968 94144
rect 65648 94062 65690 94080
rect 65926 94062 65968 94080
rect 49371 93940 49437 93941
rect 49371 93876 49372 93940
rect 49436 93876 49437 93940
rect 49371 93875 49437 93876
rect 35588 93536 35596 93600
rect 35660 93536 35676 93600
rect 35740 93536 35756 93600
rect 35820 93536 35836 93600
rect 35900 93536 35908 93600
rect 35588 92512 35908 93536
rect 42011 93260 42077 93261
rect 42011 93196 42012 93260
rect 42076 93196 42077 93260
rect 42011 93195 42077 93196
rect 39619 92716 39685 92717
rect 39619 92652 39620 92716
rect 39684 92652 39685 92716
rect 39619 92651 39685 92652
rect 38147 92580 38213 92581
rect 38147 92516 38148 92580
rect 38212 92516 38213 92580
rect 38147 92515 38213 92516
rect 35588 92448 35596 92512
rect 35660 92448 35676 92512
rect 35740 92448 35756 92512
rect 35820 92448 35836 92512
rect 35900 92448 35908 92512
rect 35588 91436 35908 92448
rect 4868 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5188 91424
rect 4868 90336 5188 91360
rect 4868 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5188 90336
rect 4868 89248 5188 90272
rect 38150 90130 38210 92515
rect 39622 90130 39682 92651
rect 42014 90130 42074 93195
rect 44587 92852 44653 92853
rect 44587 92788 44588 92852
rect 44652 92788 44653 92852
rect 44587 92787 44653 92788
rect 43299 92172 43365 92173
rect 43299 92108 43300 92172
rect 43364 92108 43365 92172
rect 43299 92107 43365 92108
rect 43302 90130 43362 92107
rect 44590 90130 44650 92787
rect 45875 92580 45941 92581
rect 45875 92516 45876 92580
rect 45940 92516 45941 92580
rect 45875 92515 45941 92516
rect 48267 92580 48333 92581
rect 48267 92516 48268 92580
rect 48332 92516 48333 92580
rect 48267 92515 48333 92516
rect 38150 90070 38220 90130
rect 38160 89420 38220 90070
rect 39520 90070 39682 90130
rect 41968 90070 42074 90130
rect 43192 90070 43362 90130
rect 44552 90070 44650 90130
rect 39520 89420 39580 90070
rect 40605 89724 40671 89725
rect 40605 89660 40606 89724
rect 40670 89660 40671 89724
rect 40605 89659 40671 89660
rect 40608 89420 40668 89659
rect 41968 89420 42028 90070
rect 43192 89420 43252 90070
rect 44552 89420 44612 90070
rect 45878 89858 45938 92515
rect 46795 92036 46861 92037
rect 46795 91972 46796 92036
rect 46860 91972 46861 92036
rect 46795 91971 46861 91972
rect 45776 89798 45938 89858
rect 46798 89858 46858 91971
rect 48270 89858 48330 92515
rect 49374 89858 49434 93875
rect 65648 93056 65968 94062
rect 65648 92992 65656 93056
rect 65720 92992 65736 93056
rect 65800 92992 65816 93056
rect 65880 92992 65896 93056
rect 65960 92992 65968 93056
rect 56915 92988 56981 92989
rect 56915 92924 56916 92988
rect 56980 92924 56981 92988
rect 56915 92923 56981 92924
rect 51947 92852 52013 92853
rect 51947 92788 51948 92852
rect 52012 92788 52013 92852
rect 51947 92787 52013 92788
rect 50659 92172 50725 92173
rect 50659 92108 50660 92172
rect 50724 92108 50725 92172
rect 50659 92107 50725 92108
rect 46798 89798 46924 89858
rect 45776 89420 45836 89798
rect 46864 89420 46924 89798
rect 48224 89798 48330 89858
rect 49312 89798 49434 89858
rect 50662 89858 50722 92107
rect 51950 89858 52010 92787
rect 53235 92172 53301 92173
rect 53235 92108 53236 92172
rect 53300 92108 53301 92172
rect 53235 92107 53301 92108
rect 50662 89798 50732 89858
rect 48224 89420 48284 89798
rect 49312 89420 49372 89798
rect 50672 89420 50732 89798
rect 51896 89798 52010 89858
rect 53238 89858 53298 92107
rect 56918 90130 56978 92923
rect 61883 92716 61949 92717
rect 61883 92652 61884 92716
rect 61948 92652 61949 92716
rect 61883 92651 61949 92652
rect 56918 90070 56988 90130
rect 55565 89860 55631 89861
rect 53238 89798 53316 89858
rect 51896 89420 51956 89798
rect 53256 89420 53316 89798
rect 55565 89796 55566 89860
rect 55630 89796 55631 89860
rect 55565 89795 55631 89796
rect 54341 89724 54407 89725
rect 54341 89660 54342 89724
rect 54406 89660 54407 89724
rect 54341 89659 54407 89660
rect 54344 89420 54404 89659
rect 55568 89420 55628 89795
rect 56928 89420 56988 90070
rect 58149 89996 58215 89997
rect 58149 89932 58150 89996
rect 58214 89932 58215 89996
rect 58149 89931 58215 89932
rect 59509 89996 59575 89997
rect 59509 89932 59510 89996
rect 59574 89932 59575 89996
rect 59509 89931 59575 89932
rect 58152 89420 58212 89931
rect 59512 89420 59572 89931
rect 61886 89730 61946 92651
rect 64275 92580 64341 92581
rect 64275 92516 64276 92580
rect 64340 92516 64341 92580
rect 64275 92515 64341 92516
rect 62987 91084 63053 91085
rect 62987 91020 62988 91084
rect 63052 91020 63053 91084
rect 62987 91019 63053 91020
rect 62990 89730 63050 91019
rect 64278 89730 64338 92515
rect 65648 91968 65968 92992
rect 65648 91904 65656 91968
rect 65720 91904 65736 91968
rect 65800 91904 65816 91968
rect 65880 91904 65896 91968
rect 65960 91904 65968 91968
rect 65648 91620 65968 91904
rect 66308 96864 66628 97424
rect 66308 96800 66316 96864
rect 66380 96800 66396 96864
rect 66460 96800 66476 96864
rect 66540 96800 66556 96864
rect 66620 96800 66628 96864
rect 66308 95776 66628 96800
rect 66308 95712 66316 95776
rect 66380 95712 66396 95776
rect 66460 95712 66476 95776
rect 66540 95712 66556 95776
rect 66620 95712 66628 95776
rect 66308 94978 66628 95712
rect 66308 94742 66350 94978
rect 66586 94742 66628 94978
rect 66308 94688 66628 94742
rect 66308 94624 66316 94688
rect 66380 94624 66396 94688
rect 66460 94624 66476 94688
rect 66540 94624 66556 94688
rect 66620 94624 66628 94688
rect 66308 93600 66628 94624
rect 66308 93536 66316 93600
rect 66380 93536 66396 93600
rect 66460 93536 66476 93600
rect 66540 93536 66556 93600
rect 66620 93536 66628 93600
rect 66308 92512 66628 93536
rect 96368 97408 96688 97424
rect 96368 97344 96376 97408
rect 96440 97344 96456 97408
rect 96520 97344 96536 97408
rect 96600 97344 96616 97408
rect 96680 97344 96688 97408
rect 96368 96320 96688 97344
rect 96368 96256 96376 96320
rect 96440 96256 96456 96320
rect 96520 96256 96536 96320
rect 96600 96256 96616 96320
rect 96680 96256 96688 96320
rect 96368 95232 96688 96256
rect 96368 95168 96376 95232
rect 96440 95168 96456 95232
rect 96520 95168 96536 95232
rect 96600 95168 96616 95232
rect 96680 95168 96688 95232
rect 96368 94298 96688 95168
rect 96368 94144 96410 94298
rect 96646 94144 96688 94298
rect 96368 94080 96376 94144
rect 96680 94080 96688 94144
rect 96368 94062 96410 94080
rect 96646 94062 96688 94080
rect 96368 93056 96688 94062
rect 96368 92992 96376 93056
rect 96440 92992 96456 93056
rect 96520 92992 96536 93056
rect 96600 92992 96616 93056
rect 96680 92992 96688 93056
rect 69243 92580 69309 92581
rect 69243 92516 69244 92580
rect 69308 92516 69309 92580
rect 69243 92515 69309 92516
rect 70715 92580 70781 92581
rect 70715 92516 70716 92580
rect 70780 92516 70781 92580
rect 70715 92515 70781 92516
rect 66308 92448 66316 92512
rect 66380 92448 66396 92512
rect 66460 92448 66476 92512
rect 66540 92448 66556 92512
rect 66620 92448 66628 92512
rect 66308 91436 66628 92448
rect 60597 89724 60663 89725
rect 60597 89660 60598 89724
rect 60662 89660 60663 89724
rect 61886 89670 62020 89730
rect 62990 89670 63108 89730
rect 60597 89659 60663 89660
rect 60600 89420 60660 89659
rect 61960 89420 62020 89670
rect 63048 89420 63108 89670
rect 64272 89670 64338 89730
rect 69246 89730 69306 92515
rect 70718 89730 70778 92515
rect 96368 91968 96688 92992
rect 96368 91904 96376 91968
rect 96440 91904 96456 91968
rect 96520 91904 96536 91968
rect 96600 91904 96616 91968
rect 96680 91904 96688 91968
rect 96368 91436 96688 91904
rect 97028 96864 97348 97424
rect 97028 96800 97036 96864
rect 97100 96800 97116 96864
rect 97180 96800 97196 96864
rect 97260 96800 97276 96864
rect 97340 96800 97348 96864
rect 97028 95776 97348 96800
rect 97028 95712 97036 95776
rect 97100 95712 97116 95776
rect 97180 95712 97196 95776
rect 97260 95712 97276 95776
rect 97340 95712 97348 95776
rect 97028 94978 97348 95712
rect 97028 94742 97070 94978
rect 97306 94742 97348 94978
rect 97028 94688 97348 94742
rect 97028 94624 97036 94688
rect 97100 94624 97116 94688
rect 97180 94624 97196 94688
rect 97260 94624 97276 94688
rect 97340 94624 97348 94688
rect 97028 93600 97348 94624
rect 97028 93536 97036 93600
rect 97100 93536 97116 93600
rect 97180 93536 97196 93600
rect 97260 93536 97276 93600
rect 97340 93536 97348 93600
rect 97028 92512 97348 93536
rect 97028 92448 97036 92512
rect 97100 92448 97116 92512
rect 97180 92448 97196 92512
rect 97260 92448 97276 92512
rect 97340 92448 97348 92512
rect 97028 91436 97348 92448
rect 112908 91968 113228 92528
rect 112908 91904 112916 91968
rect 112980 91904 112996 91968
rect 113060 91904 113076 91968
rect 113140 91904 113156 91968
rect 113220 91904 113228 91968
rect 99971 91220 100037 91221
rect 99971 91156 99972 91220
rect 100036 91156 100037 91220
rect 99971 91155 100037 91156
rect 73291 91084 73357 91085
rect 73291 91020 73292 91084
rect 73356 91020 73357 91084
rect 73291 91019 73357 91020
rect 74211 91084 74277 91085
rect 74211 91020 74212 91084
rect 74276 91020 74277 91084
rect 74211 91019 74277 91020
rect 73294 89730 73354 91019
rect 65629 89724 65695 89725
rect 64272 89420 64332 89670
rect 65629 89660 65630 89724
rect 65694 89660 65695 89724
rect 65629 89659 65695 89660
rect 66853 89724 66919 89725
rect 66853 89660 66854 89724
rect 66918 89660 66919 89724
rect 66853 89659 66919 89660
rect 68213 89724 68279 89725
rect 68213 89660 68214 89724
rect 68278 89660 68279 89724
rect 69246 89670 69364 89730
rect 68213 89659 68279 89660
rect 65632 89420 65692 89659
rect 66856 89420 66916 89659
rect 68216 89420 68276 89659
rect 69304 89420 69364 89670
rect 70664 89670 70778 89730
rect 71885 89724 71951 89725
rect 70664 89420 70724 89670
rect 71885 89660 71886 89724
rect 71950 89660 71951 89724
rect 71885 89659 71951 89660
rect 73248 89670 73354 89730
rect 74214 89730 74274 91019
rect 99974 90130 100034 91155
rect 112908 90880 113228 91904
rect 112908 90816 112916 90880
rect 112980 90816 112996 90880
rect 113060 90816 113076 90880
rect 113140 90816 113156 90880
rect 113220 90816 113228 90880
rect 99974 90070 100100 90130
rect 74214 89670 74396 89730
rect 71888 89420 71948 89659
rect 73248 89420 73308 89670
rect 74336 89420 74396 89670
rect 75557 89724 75623 89725
rect 75557 89660 75558 89724
rect 75622 89660 75623 89724
rect 75557 89659 75623 89660
rect 76917 89724 76983 89725
rect 76917 89660 76918 89724
rect 76982 89660 76983 89724
rect 76917 89659 76983 89660
rect 89429 89724 89495 89725
rect 89429 89660 89430 89724
rect 89494 89660 89495 89724
rect 89429 89659 89495 89660
rect 75560 89420 75620 89659
rect 76920 89420 76980 89659
rect 89432 89420 89492 89659
rect 100040 89420 100100 90070
rect 112908 89792 113228 90816
rect 112908 89728 112916 89792
rect 112980 89728 112996 89792
rect 113060 89728 113076 89792
rect 113140 89728 113156 89792
rect 113220 89728 113228 89792
rect 4868 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5188 89248
rect 4868 88160 5188 89184
rect 4868 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5188 88160
rect 4868 87072 5188 88096
rect 4868 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5188 87072
rect 4868 85984 5188 87008
rect 4868 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5188 85984
rect 4868 84896 5188 85920
rect 4868 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5188 84896
rect 4868 83808 5188 84832
rect 4868 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5188 83808
rect 4868 82720 5188 83744
rect 4868 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5188 82720
rect 4868 81632 5188 82656
rect 4868 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5188 81632
rect 4868 80544 5188 81568
rect 4868 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5188 80544
rect 4868 79456 5188 80480
rect 4868 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5188 79456
rect 4868 78368 5188 79392
rect 4868 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5188 78368
rect 4868 77280 5188 78304
rect 4868 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5188 77280
rect 4868 76192 5188 77216
rect 4868 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5188 76192
rect 4868 75104 5188 76128
rect 4868 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5188 75104
rect 4868 74016 5188 75040
rect 4868 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5188 74016
rect 4868 72928 5188 73952
rect 4868 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5188 72928
rect 4868 71840 5188 72864
rect 4868 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5188 71840
rect 4868 70752 5188 71776
rect 4868 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5188 70752
rect 4868 69664 5188 70688
rect 4868 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5188 69664
rect 4868 68576 5188 69600
rect 4868 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5188 68576
rect 4868 67556 5188 68512
rect 112908 88704 113228 89728
rect 112908 88640 112916 88704
rect 112980 88640 112996 88704
rect 113060 88640 113076 88704
rect 113140 88640 113156 88704
rect 113220 88640 113228 88704
rect 112908 87616 113228 88640
rect 112908 87552 112916 87616
rect 112980 87552 112996 87616
rect 113060 87552 113076 87616
rect 113140 87552 113156 87616
rect 113220 87552 113228 87616
rect 112908 86528 113228 87552
rect 112908 86464 112916 86528
rect 112980 86464 112996 86528
rect 113060 86464 113076 86528
rect 113140 86464 113156 86528
rect 113220 86464 113228 86528
rect 112908 85440 113228 86464
rect 112908 85376 112916 85440
rect 112980 85376 112996 85440
rect 113060 85376 113076 85440
rect 113140 85376 113156 85440
rect 113220 85376 113228 85440
rect 112908 84352 113228 85376
rect 112908 84288 112916 84352
rect 112980 84288 112996 84352
rect 113060 84288 113076 84352
rect 113140 84288 113156 84352
rect 113220 84288 113228 84352
rect 112908 83264 113228 84288
rect 112908 83200 112916 83264
rect 112980 83200 112996 83264
rect 113060 83200 113076 83264
rect 113140 83200 113156 83264
rect 113220 83200 113228 83264
rect 112908 82176 113228 83200
rect 112908 82112 112916 82176
rect 112980 82112 112996 82176
rect 113060 82112 113076 82176
rect 113140 82112 113156 82176
rect 113220 82112 113228 82176
rect 112908 81088 113228 82112
rect 112908 81024 112916 81088
rect 112980 81024 112996 81088
rect 113060 81024 113076 81088
rect 113140 81024 113156 81088
rect 113220 81024 113228 81088
rect 112908 80000 113228 81024
rect 112908 79936 112916 80000
rect 112980 79936 112996 80000
rect 113060 79936 113076 80000
rect 113140 79936 113156 80000
rect 113220 79936 113228 80000
rect 112908 78912 113228 79936
rect 112908 78848 112916 78912
rect 112980 78848 112996 78912
rect 113060 78848 113076 78912
rect 113140 78848 113156 78912
rect 113220 78848 113228 78912
rect 112908 77824 113228 78848
rect 112908 77760 112916 77824
rect 112980 77760 112996 77824
rect 113060 77760 113076 77824
rect 113140 77760 113156 77824
rect 113220 77760 113228 77824
rect 112908 76736 113228 77760
rect 112908 76672 112916 76736
rect 112980 76672 112996 76736
rect 113060 76672 113076 76736
rect 113140 76672 113156 76736
rect 113220 76672 113228 76736
rect 112908 75648 113228 76672
rect 112908 75584 112916 75648
rect 112980 75584 112996 75648
rect 113060 75584 113076 75648
rect 113140 75584 113156 75648
rect 113220 75584 113228 75648
rect 112908 74560 113228 75584
rect 112908 74496 112916 74560
rect 112980 74496 112996 74560
rect 113060 74496 113076 74560
rect 113140 74496 113156 74560
rect 113220 74496 113228 74560
rect 112908 73472 113228 74496
rect 112908 73408 112916 73472
rect 112980 73408 112996 73472
rect 113060 73408 113076 73472
rect 113140 73408 113156 73472
rect 113220 73408 113228 73472
rect 112908 72384 113228 73408
rect 112908 72320 112916 72384
rect 112980 72320 112996 72384
rect 113060 72320 113076 72384
rect 113140 72320 113156 72384
rect 113220 72320 113228 72384
rect 112908 71296 113228 72320
rect 112908 71232 112916 71296
rect 112980 71232 112996 71296
rect 113060 71232 113076 71296
rect 113140 71232 113156 71296
rect 113220 71232 113228 71296
rect 112908 70208 113228 71232
rect 112908 70144 112916 70208
rect 112980 70144 112996 70208
rect 113060 70144 113076 70208
rect 113140 70144 113156 70208
rect 113220 70144 113228 70208
rect 112908 69120 113228 70144
rect 112908 69056 112916 69120
rect 112980 69056 112996 69120
rect 113060 69056 113076 69120
rect 113140 69056 113156 69120
rect 113220 69056 113228 69120
rect 112908 68032 113228 69056
rect 112908 67968 112916 68032
rect 112980 67968 112996 68032
rect 113060 67968 113076 68032
rect 113140 67968 113156 68032
rect 113220 67968 113228 68032
rect 4868 67488 4910 67556
rect 5146 67488 5188 67556
rect 4868 67424 4876 67488
rect 5180 67424 5188 67488
rect 4868 67320 4910 67424
rect 5146 67320 5188 67424
rect 4868 66400 5188 67320
rect 10272 67556 10620 67598
rect 10272 67320 10328 67556
rect 10564 67320 10620 67556
rect 10272 67278 10620 67320
rect 105336 67556 105684 67598
rect 105336 67320 105392 67556
rect 105628 67320 105684 67556
rect 105336 67278 105684 67320
rect 112908 66944 113228 67968
rect 10952 66896 11300 66938
rect 10952 66660 11008 66896
rect 11244 66660 11300 66896
rect 10952 66618 11300 66660
rect 104656 66896 105004 66938
rect 104656 66660 104712 66896
rect 104948 66660 105004 66896
rect 104656 66618 105004 66660
rect 112908 66880 112916 66944
rect 112980 66896 112996 66944
rect 113060 66896 113076 66944
rect 113140 66896 113156 66944
rect 113220 66880 113228 66944
rect 112908 66660 112950 66880
rect 113186 66660 113228 66880
rect 4868 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5188 66400
rect 4868 65312 5188 66336
rect 4868 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5188 65312
rect 4868 64224 5188 65248
rect 4868 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5188 64224
rect 4868 63136 5188 64160
rect 4868 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5188 63136
rect 4868 62048 5188 63072
rect 4868 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5188 62048
rect 4868 60960 5188 61984
rect 4868 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5188 60960
rect 4868 59872 5188 60896
rect 4868 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5188 59872
rect 4868 58784 5188 59808
rect 4868 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5188 58784
rect 4868 57696 5188 58720
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 112908 65856 113228 66660
rect 112908 65792 112916 65856
rect 112980 65792 112996 65856
rect 113060 65792 113076 65856
rect 113140 65792 113156 65856
rect 113220 65792 113228 65856
rect 112908 64768 113228 65792
rect 112908 64704 112916 64768
rect 112980 64704 112996 64768
rect 113060 64704 113076 64768
rect 113140 64704 113156 64768
rect 113220 64704 113228 64768
rect 112908 63680 113228 64704
rect 112908 63616 112916 63680
rect 112980 63616 112996 63680
rect 113060 63616 113076 63680
rect 113140 63616 113156 63680
rect 113220 63616 113228 63680
rect 112908 62592 113228 63616
rect 112908 62528 112916 62592
rect 112980 62528 112996 62592
rect 113060 62528 113076 62592
rect 113140 62528 113156 62592
rect 113220 62528 113228 62592
rect 112908 61504 113228 62528
rect 112908 61440 112916 61504
rect 112980 61440 112996 61504
rect 113060 61440 113076 61504
rect 113140 61440 113156 61504
rect 113220 61440 113228 61504
rect 112908 60416 113228 61440
rect 112908 60352 112916 60416
rect 112980 60352 112996 60416
rect 113060 60352 113076 60416
rect 113140 60352 113156 60416
rect 113220 60352 113228 60416
rect 112908 59328 113228 60352
rect 112908 59264 112916 59328
rect 112980 59264 112996 59328
rect 113060 59264 113076 59328
rect 113140 59264 113156 59328
rect 113220 59264 113228 59328
rect 112908 58240 113228 59264
rect 112908 58176 112916 58240
rect 112980 58176 112996 58240
rect 113060 58176 113076 58240
rect 113140 58176 113156 58240
rect 113220 58176 113228 58240
rect 112908 57152 113228 58176
rect 112908 57088 112916 57152
rect 112980 57088 112996 57152
rect 113060 57088 113076 57152
rect 113140 57088 113156 57152
rect 113220 57088 113228 57152
rect 112908 56064 113228 57088
rect 112908 56000 112916 56064
rect 112980 56000 112996 56064
rect 113060 56000 113076 56064
rect 113140 56000 113156 56064
rect 113220 56000 113228 56064
rect 112908 54976 113228 56000
rect 112908 54912 112916 54976
rect 112980 54912 112996 54976
rect 113060 54912 113076 54976
rect 113140 54912 113156 54976
rect 113220 54912 113228 54976
rect 112908 53888 113228 54912
rect 112908 53824 112916 53888
rect 112980 53824 112996 53888
rect 113060 53824 113076 53888
rect 113140 53824 113156 53888
rect 113220 53824 113228 53888
rect 112908 52800 113228 53824
rect 112908 52736 112916 52800
rect 112980 52736 112996 52800
rect 113060 52736 113076 52800
rect 113140 52736 113156 52800
rect 113220 52736 113228 52800
rect 112908 51712 113228 52736
rect 112908 51648 112916 51712
rect 112980 51648 112996 51712
rect 113060 51648 113076 51712
rect 113140 51648 113156 51712
rect 113220 51648 113228 51712
rect 112908 50624 113228 51648
rect 112908 50560 112916 50624
rect 112980 50560 112996 50624
rect 113060 50560 113076 50624
rect 113140 50560 113156 50624
rect 113220 50560 113228 50624
rect 112908 49536 113228 50560
rect 112908 49472 112916 49536
rect 112980 49472 112996 49536
rect 113060 49472 113076 49536
rect 113140 49472 113156 49536
rect 113220 49472 113228 49536
rect 112908 48448 113228 49472
rect 112908 48384 112916 48448
rect 112980 48384 112996 48448
rect 113060 48384 113076 48448
rect 113140 48384 113156 48448
rect 113220 48384 113228 48448
rect 112908 47360 113228 48384
rect 112908 47296 112916 47360
rect 112980 47296 112996 47360
rect 113060 47296 113076 47360
rect 113140 47296 113156 47360
rect 113220 47296 113228 47360
rect 112908 46272 113228 47296
rect 112908 46208 112916 46272
rect 112980 46208 112996 46272
rect 113060 46208 113076 46272
rect 113140 46208 113156 46272
rect 113220 46208 113228 46272
rect 112908 45184 113228 46208
rect 112908 45120 112916 45184
rect 112980 45120 112996 45184
rect 113060 45120 113076 45184
rect 113140 45120 113156 45184
rect 113220 45120 113228 45184
rect 112908 44096 113228 45120
rect 112908 44032 112916 44096
rect 112980 44032 112996 44096
rect 113060 44032 113076 44096
rect 113140 44032 113156 44096
rect 113220 44032 113228 44096
rect 112908 43008 113228 44032
rect 112908 42944 112916 43008
rect 112980 42944 112996 43008
rect 113060 42944 113076 43008
rect 113140 42944 113156 43008
rect 113220 42944 113228 43008
rect 112908 41920 113228 42944
rect 112908 41856 112916 41920
rect 112980 41856 112996 41920
rect 113060 41856 113076 41920
rect 113140 41856 113156 41920
rect 113220 41856 113228 41920
rect 112908 40832 113228 41856
rect 112908 40768 112916 40832
rect 112980 40768 112996 40832
rect 113060 40768 113076 40832
rect 113140 40768 113156 40832
rect 113220 40768 113228 40832
rect 112908 39744 113228 40768
rect 112908 39680 112916 39744
rect 112980 39680 112996 39744
rect 113060 39680 113076 39744
rect 113140 39680 113156 39744
rect 113220 39680 113228 39744
rect 112908 38656 113228 39680
rect 112908 38592 112916 38656
rect 112980 38592 112996 38656
rect 113060 38592 113076 38656
rect 113140 38592 113156 38656
rect 113220 38592 113228 38656
rect 112908 37568 113228 38592
rect 112908 37504 112916 37568
rect 112980 37504 112996 37568
rect 113060 37504 113076 37568
rect 113140 37504 113156 37568
rect 113220 37504 113228 37568
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 10272 36920 10620 36962
rect 10272 36684 10328 36920
rect 10564 36684 10620 36920
rect 10272 36642 10620 36684
rect 105336 36920 105684 36962
rect 105336 36684 105392 36920
rect 105628 36684 105684 36920
rect 105336 36642 105684 36684
rect 112908 36480 113228 37504
rect 112908 36416 112916 36480
rect 112980 36416 112996 36480
rect 113060 36416 113076 36480
rect 113140 36416 113156 36480
rect 113220 36416 113228 36480
rect 10952 36260 11300 36302
rect 10952 36024 11008 36260
rect 11244 36024 11300 36260
rect 10952 35982 11300 36024
rect 104656 36260 105004 36302
rect 104656 36024 104712 36260
rect 104948 36024 105004 36260
rect 104656 35982 105004 36024
rect 112908 36260 113228 36416
rect 112908 36024 112950 36260
rect 113186 36024 113228 36260
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 112908 35392 113228 36024
rect 112908 35328 112916 35392
rect 112980 35328 112996 35392
rect 113060 35328 113076 35392
rect 113140 35328 113156 35392
rect 113220 35328 113228 35392
rect 112908 34304 113228 35328
rect 112908 34240 112916 34304
rect 112980 34240 112996 34304
rect 113060 34240 113076 34304
rect 113140 34240 113156 34304
rect 113220 34240 113228 34304
rect 109355 33284 109421 33285
rect 109355 33220 109356 33284
rect 109420 33220 109421 33284
rect 109355 33219 109421 33220
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 109358 11933 109418 33219
rect 112908 33216 113228 34240
rect 112908 33152 112916 33216
rect 112980 33152 112996 33216
rect 113060 33152 113076 33216
rect 113140 33152 113156 33216
rect 113220 33152 113228 33216
rect 112908 32128 113228 33152
rect 112908 32064 112916 32128
rect 112980 32064 112996 32128
rect 113060 32064 113076 32128
rect 113140 32064 113156 32128
rect 113220 32064 113228 32128
rect 112908 31040 113228 32064
rect 112908 30976 112916 31040
rect 112980 30976 112996 31040
rect 113060 30976 113076 31040
rect 113140 30976 113156 31040
rect 113220 30976 113228 31040
rect 112908 29952 113228 30976
rect 112908 29888 112916 29952
rect 112980 29888 112996 29952
rect 113060 29888 113076 29952
rect 113140 29888 113156 29952
rect 113220 29888 113228 29952
rect 112908 28864 113228 29888
rect 112908 28800 112916 28864
rect 112980 28800 112996 28864
rect 113060 28800 113076 28864
rect 113140 28800 113156 28864
rect 113220 28800 113228 28864
rect 112908 27776 113228 28800
rect 112908 27712 112916 27776
rect 112980 27712 112996 27776
rect 113060 27712 113076 27776
rect 113140 27712 113156 27776
rect 113220 27712 113228 27776
rect 112908 26688 113228 27712
rect 112908 26624 112916 26688
rect 112980 26624 112996 26688
rect 113060 26624 113076 26688
rect 113140 26624 113156 26688
rect 113220 26624 113228 26688
rect 112908 25600 113228 26624
rect 112908 25536 112916 25600
rect 112980 25536 112996 25600
rect 113060 25536 113076 25600
rect 113140 25536 113156 25600
rect 113220 25536 113228 25600
rect 112908 24512 113228 25536
rect 112908 24448 112916 24512
rect 112980 24448 112996 24512
rect 113060 24448 113076 24512
rect 113140 24448 113156 24512
rect 113220 24448 113228 24512
rect 112908 23424 113228 24448
rect 112908 23360 112916 23424
rect 112980 23360 112996 23424
rect 113060 23360 113076 23424
rect 113140 23360 113156 23424
rect 113220 23360 113228 23424
rect 112908 22336 113228 23360
rect 112908 22272 112916 22336
rect 112980 22272 112996 22336
rect 113060 22272 113076 22336
rect 113140 22272 113156 22336
rect 113220 22272 113228 22336
rect 112908 21248 113228 22272
rect 112908 21184 112916 21248
rect 112980 21184 112996 21248
rect 113060 21184 113076 21248
rect 113140 21184 113156 21248
rect 113220 21184 113228 21248
rect 112908 20160 113228 21184
rect 112908 20096 112916 20160
rect 112980 20096 112996 20160
rect 113060 20096 113076 20160
rect 113140 20096 113156 20160
rect 113220 20096 113228 20160
rect 112908 19072 113228 20096
rect 112908 19008 112916 19072
rect 112980 19008 112996 19072
rect 113060 19008 113076 19072
rect 113140 19008 113156 19072
rect 113220 19008 113228 19072
rect 112908 17984 113228 19008
rect 112908 17920 112916 17984
rect 112980 17920 112996 17984
rect 113060 17920 113076 17984
rect 113140 17920 113156 17984
rect 113220 17920 113228 17984
rect 112908 16896 113228 17920
rect 112908 16832 112916 16896
rect 112980 16832 112996 16896
rect 113060 16832 113076 16896
rect 113140 16832 113156 16896
rect 113220 16832 113228 16896
rect 112908 15808 113228 16832
rect 112908 15744 112916 15808
rect 112980 15744 112996 15808
rect 113060 15744 113076 15808
rect 113140 15744 113156 15808
rect 113220 15744 113228 15808
rect 112908 14720 113228 15744
rect 112908 14656 112916 14720
rect 112980 14656 112996 14720
rect 113060 14656 113076 14720
rect 113140 14656 113156 14720
rect 113220 14656 113228 14720
rect 112908 13632 113228 14656
rect 112908 13568 112916 13632
rect 112980 13568 112996 13632
rect 113060 13568 113076 13632
rect 113140 13568 113156 13632
rect 113220 13568 113228 13632
rect 112908 12544 113228 13568
rect 112908 12480 112916 12544
rect 112980 12480 112996 12544
rect 113060 12480 113076 12544
rect 113140 12480 113156 12544
rect 113220 12480 113228 12544
rect 109355 11932 109421 11933
rect 109355 11868 109356 11932
rect 109420 11868 109421 11932
rect 109355 11867 109421 11868
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 112908 11456 113228 12480
rect 112908 11392 112916 11456
rect 112980 11392 112996 11456
rect 113060 11392 113076 11456
rect 113140 11392 113156 11456
rect 113220 11392 113228 11456
rect 112908 10368 113228 11392
rect 112908 10304 112916 10368
rect 112980 10304 112996 10368
rect 113060 10304 113076 10368
rect 113140 10304 113156 10368
rect 113220 10304 113228 10368
rect 15856 9893 15916 10106
rect 15853 9892 15919 9893
rect 15853 9828 15854 9892
rect 15918 9828 15919 9892
rect 25512 9890 25572 10106
rect 15853 9827 15919 9828
rect 25454 9830 25572 9890
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 25454 8261 25514 9830
rect 26736 9757 26796 10106
rect 27824 9757 27884 10106
rect 29184 9757 29244 10106
rect 30136 9757 30196 10106
rect 31360 9890 31420 10106
rect 31342 9830 31420 9890
rect 32584 9890 32644 10106
rect 33672 9890 33732 10106
rect 35032 9890 35092 10106
rect 32584 9830 32690 9890
rect 33672 9830 33794 9890
rect 26733 9756 26799 9757
rect 26733 9692 26734 9756
rect 26798 9692 26799 9756
rect 26733 9691 26799 9692
rect 27821 9756 27887 9757
rect 27821 9692 27822 9756
rect 27886 9692 27887 9756
rect 27821 9691 27887 9692
rect 29181 9756 29247 9757
rect 29181 9692 29182 9756
rect 29246 9692 29247 9756
rect 29181 9691 29247 9692
rect 30133 9756 30199 9757
rect 30133 9692 30134 9756
rect 30198 9692 30199 9756
rect 30133 9691 30199 9692
rect 31342 8261 31402 9830
rect 32630 8261 32690 9830
rect 33734 8261 33794 9830
rect 35022 9830 35092 9890
rect 36120 9890 36180 10106
rect 37208 9890 37268 10106
rect 38296 9890 38356 10106
rect 39656 9890 39716 10106
rect 40744 9890 40804 10106
rect 41832 9890 41892 10106
rect 36120 9830 36186 9890
rect 37208 9830 37290 9890
rect 38296 9830 38394 9890
rect 35022 8261 35082 9830
rect 36126 8261 36186 9830
rect 37230 8261 37290 9830
rect 38334 8261 38394 9830
rect 39622 9830 39716 9890
rect 40726 9830 40804 9890
rect 41830 9830 41892 9890
rect 43056 9890 43116 10106
rect 44144 9890 44204 10106
rect 45504 9890 45564 10106
rect 43056 9830 43178 9890
rect 44144 9830 44282 9890
rect 25451 8260 25517 8261
rect 25451 8196 25452 8260
rect 25516 8196 25517 8260
rect 25451 8195 25517 8196
rect 31339 8260 31405 8261
rect 31339 8196 31340 8260
rect 31404 8196 31405 8260
rect 31339 8195 31405 8196
rect 32627 8260 32693 8261
rect 32627 8196 32628 8260
rect 32692 8196 32693 8260
rect 32627 8195 32693 8196
rect 33731 8260 33797 8261
rect 33731 8196 33732 8260
rect 33796 8196 33797 8260
rect 33731 8195 33797 8196
rect 35019 8260 35085 8261
rect 35019 8196 35020 8260
rect 35084 8196 35085 8260
rect 35019 8195 35085 8196
rect 36123 8260 36189 8261
rect 36123 8196 36124 8260
rect 36188 8196 36189 8260
rect 36123 8195 36189 8196
rect 37227 8260 37293 8261
rect 37227 8196 37228 8260
rect 37292 8196 37293 8260
rect 37227 8195 37293 8196
rect 38331 8260 38397 8261
rect 38331 8196 38332 8260
rect 38396 8196 38397 8260
rect 38331 8195 38397 8196
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 7104 35248 7880
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 7648 35908 8064
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 39622 2685 39682 9830
rect 40726 8261 40786 9830
rect 41830 8261 41890 9830
rect 43118 8261 43178 9830
rect 44222 8261 44282 9830
rect 45326 9830 45564 9890
rect 46592 9890 46652 10106
rect 47680 9890 47740 10106
rect 48904 9890 48964 10106
rect 50264 9890 50324 10106
rect 46592 9830 46674 9890
rect 47680 9830 47778 9890
rect 48904 9830 49066 9890
rect 50264 9830 50354 9890
rect 40723 8260 40789 8261
rect 40723 8196 40724 8260
rect 40788 8196 40789 8260
rect 40723 8195 40789 8196
rect 41827 8260 41893 8261
rect 41827 8196 41828 8260
rect 41892 8196 41893 8260
rect 41827 8195 41893 8196
rect 43115 8260 43181 8261
rect 43115 8196 43116 8260
rect 43180 8196 43181 8260
rect 43115 8195 43181 8196
rect 44219 8260 44285 8261
rect 44219 8196 44220 8260
rect 44284 8196 44285 8260
rect 44219 8195 44285 8196
rect 45326 7170 45386 9830
rect 46614 8261 46674 9830
rect 47718 8261 47778 9830
rect 49006 8261 49066 9830
rect 50294 8261 50354 9830
rect 51352 9757 51412 10106
rect 52440 9757 52500 10106
rect 53528 9757 53588 10106
rect 54888 9757 54948 10106
rect 55976 9757 56036 10106
rect 57064 9757 57124 10106
rect 58288 9757 58348 10106
rect 59376 9757 59436 10106
rect 60736 9890 60796 10106
rect 60736 9830 60842 9890
rect 60782 9757 60842 9830
rect 51349 9756 51415 9757
rect 51349 9692 51350 9756
rect 51414 9692 51415 9756
rect 51349 9691 51415 9692
rect 52437 9756 52503 9757
rect 52437 9692 52438 9756
rect 52502 9692 52503 9756
rect 52437 9691 52503 9692
rect 53525 9756 53591 9757
rect 53525 9692 53526 9756
rect 53590 9692 53591 9756
rect 53525 9691 53591 9692
rect 54885 9756 54951 9757
rect 54885 9692 54886 9756
rect 54950 9692 54951 9756
rect 54885 9691 54951 9692
rect 55973 9756 56039 9757
rect 55973 9692 55974 9756
rect 56038 9692 56039 9756
rect 55973 9691 56039 9692
rect 57061 9756 57127 9757
rect 57061 9692 57062 9756
rect 57126 9692 57127 9756
rect 57061 9691 57127 9692
rect 58285 9756 58351 9757
rect 58285 9692 58286 9756
rect 58350 9692 58351 9756
rect 58285 9691 58351 9692
rect 59373 9756 59439 9757
rect 59373 9692 59374 9756
rect 59438 9692 59439 9756
rect 59373 9691 59439 9692
rect 60779 9756 60845 9757
rect 60779 9692 60780 9756
rect 60844 9692 60845 9756
rect 60779 9691 60845 9692
rect 61824 9690 61884 10106
rect 62912 9690 62972 10106
rect 64000 9690 64060 10106
rect 65224 9890 65284 10106
rect 65198 9830 65284 9890
rect 66584 9890 66644 10106
rect 66584 9830 66730 9890
rect 61824 9630 61946 9690
rect 62912 9630 63050 9690
rect 64000 9630 64154 9690
rect 61886 8261 61946 9630
rect 62990 8261 63050 9630
rect 64094 8261 64154 9630
rect 65198 8261 65258 9830
rect 66670 8261 66730 9830
rect 67672 9757 67732 10106
rect 92696 9893 92756 10106
rect 92693 9892 92759 9893
rect 92693 9828 92694 9892
rect 92758 9828 92759 9892
rect 92693 9827 92759 9828
rect 92832 9757 92892 10106
rect 92968 9893 93028 10106
rect 93104 9893 93164 10106
rect 93347 10028 93413 10029
rect 93347 9964 93348 10028
rect 93412 9964 93413 10028
rect 93347 9963 93413 9964
rect 92965 9892 93031 9893
rect 92965 9828 92966 9892
rect 93030 9828 93031 9892
rect 92965 9827 93031 9828
rect 93101 9892 93167 9893
rect 93101 9828 93102 9892
rect 93166 9828 93167 9892
rect 93101 9827 93167 9828
rect 67669 9756 67735 9757
rect 67669 9692 67670 9756
rect 67734 9692 67735 9756
rect 67669 9691 67735 9692
rect 92829 9756 92895 9757
rect 92829 9692 92830 9756
rect 92894 9692 92895 9756
rect 92829 9691 92895 9692
rect 93350 8261 93410 9963
rect 112908 9280 113228 10304
rect 112908 9216 112916 9280
rect 112980 9216 112996 9280
rect 113060 9216 113076 9280
rect 113140 9216 113156 9280
rect 113220 9216 113228 9280
rect 46611 8260 46677 8261
rect 46611 8196 46612 8260
rect 46676 8196 46677 8260
rect 46611 8195 46677 8196
rect 47715 8260 47781 8261
rect 47715 8196 47716 8260
rect 47780 8196 47781 8260
rect 47715 8195 47781 8196
rect 49003 8260 49069 8261
rect 49003 8196 49004 8260
rect 49068 8196 49069 8260
rect 49003 8195 49069 8196
rect 50291 8260 50357 8261
rect 50291 8196 50292 8260
rect 50356 8196 50357 8260
rect 50291 8195 50357 8196
rect 61883 8260 61949 8261
rect 61883 8196 61884 8260
rect 61948 8196 61949 8260
rect 61883 8195 61949 8196
rect 62987 8260 63053 8261
rect 62987 8196 62988 8260
rect 63052 8196 63053 8260
rect 62987 8195 63053 8196
rect 64091 8260 64157 8261
rect 64091 8196 64092 8260
rect 64156 8196 64157 8260
rect 64091 8195 64157 8196
rect 65195 8260 65261 8261
rect 65195 8196 65196 8260
rect 65260 8196 65261 8260
rect 65195 8195 65261 8196
rect 66667 8260 66733 8261
rect 66667 8196 66668 8260
rect 66732 8196 66733 8260
rect 66667 8195 66733 8196
rect 93347 8260 93413 8261
rect 93347 8196 93348 8260
rect 93412 8196 93413 8260
rect 93347 8195 93413 8196
rect 112908 8192 113228 9216
rect 112908 8128 112916 8192
rect 112980 8128 112996 8192
rect 113060 8128 113076 8192
rect 113140 8128 113156 8192
rect 113220 8128 113228 8192
rect 45507 7172 45573 7173
rect 45507 7170 45508 7172
rect 45326 7110 45508 7170
rect 45507 7108 45508 7110
rect 45572 7108 45573 7172
rect 45507 7107 45573 7108
rect 65648 7104 65968 7880
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5624 65968 5952
rect 65648 5388 65690 5624
rect 65926 5388 65968 5624
rect 65648 4928 65968 5388
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 39619 2684 39685 2685
rect 39619 2620 39620 2684
rect 39684 2620 39685 2684
rect 39619 2619 39685 2620
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
rect 65648 2128 65968 2688
rect 66308 7648 66628 7880
rect 66308 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66628 7648
rect 66308 6560 66628 7584
rect 66308 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66628 6560
rect 66308 6284 66628 6496
rect 66308 6048 66350 6284
rect 66586 6048 66628 6284
rect 66308 5472 66628 6048
rect 66308 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66628 5472
rect 66308 4384 66628 5408
rect 66308 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66628 4384
rect 66308 3296 66628 4320
rect 66308 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66628 3296
rect 66308 2208 66628 3232
rect 66308 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66628 2208
rect 66308 2128 66628 2144
rect 96368 7104 96688 8064
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 5624 96688 5952
rect 96368 5388 96410 5624
rect 96646 5388 96688 5624
rect 96368 4928 96688 5388
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2128 96688 2688
rect 97028 7648 97348 8064
rect 97028 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97348 7648
rect 97028 6560 97348 7584
rect 112908 7104 113228 8128
rect 112908 7040 112916 7104
rect 112980 7040 112996 7104
rect 113060 7040 113076 7104
rect 113140 7040 113156 7104
rect 113220 7040 113228 7104
rect 112908 7024 113228 7040
rect 113644 92512 113964 92528
rect 113644 92448 113652 92512
rect 113716 92448 113732 92512
rect 113796 92448 113812 92512
rect 113876 92448 113892 92512
rect 113956 92448 113964 92512
rect 113644 91424 113964 92448
rect 113644 91360 113652 91424
rect 113716 91360 113732 91424
rect 113796 91360 113812 91424
rect 113876 91360 113892 91424
rect 113956 91360 113964 91424
rect 113644 90336 113964 91360
rect 113644 90272 113652 90336
rect 113716 90272 113732 90336
rect 113796 90272 113812 90336
rect 113876 90272 113892 90336
rect 113956 90272 113964 90336
rect 113644 89248 113964 90272
rect 113644 89184 113652 89248
rect 113716 89184 113732 89248
rect 113796 89184 113812 89248
rect 113876 89184 113892 89248
rect 113956 89184 113964 89248
rect 113644 88160 113964 89184
rect 113644 88096 113652 88160
rect 113716 88096 113732 88160
rect 113796 88096 113812 88160
rect 113876 88096 113892 88160
rect 113956 88096 113964 88160
rect 113644 87072 113964 88096
rect 113644 87008 113652 87072
rect 113716 87008 113732 87072
rect 113796 87008 113812 87072
rect 113876 87008 113892 87072
rect 113956 87008 113964 87072
rect 113644 85984 113964 87008
rect 113644 85920 113652 85984
rect 113716 85920 113732 85984
rect 113796 85920 113812 85984
rect 113876 85920 113892 85984
rect 113956 85920 113964 85984
rect 113644 84896 113964 85920
rect 113644 84832 113652 84896
rect 113716 84832 113732 84896
rect 113796 84832 113812 84896
rect 113876 84832 113892 84896
rect 113956 84832 113964 84896
rect 113644 83808 113964 84832
rect 113644 83744 113652 83808
rect 113716 83744 113732 83808
rect 113796 83744 113812 83808
rect 113876 83744 113892 83808
rect 113956 83744 113964 83808
rect 113644 82720 113964 83744
rect 113644 82656 113652 82720
rect 113716 82656 113732 82720
rect 113796 82656 113812 82720
rect 113876 82656 113892 82720
rect 113956 82656 113964 82720
rect 113644 81632 113964 82656
rect 113644 81568 113652 81632
rect 113716 81568 113732 81632
rect 113796 81568 113812 81632
rect 113876 81568 113892 81632
rect 113956 81568 113964 81632
rect 113644 80544 113964 81568
rect 113644 80480 113652 80544
rect 113716 80480 113732 80544
rect 113796 80480 113812 80544
rect 113876 80480 113892 80544
rect 113956 80480 113964 80544
rect 113644 79456 113964 80480
rect 113644 79392 113652 79456
rect 113716 79392 113732 79456
rect 113796 79392 113812 79456
rect 113876 79392 113892 79456
rect 113956 79392 113964 79456
rect 113644 78368 113964 79392
rect 113644 78304 113652 78368
rect 113716 78304 113732 78368
rect 113796 78304 113812 78368
rect 113876 78304 113892 78368
rect 113956 78304 113964 78368
rect 113644 77280 113964 78304
rect 113644 77216 113652 77280
rect 113716 77216 113732 77280
rect 113796 77216 113812 77280
rect 113876 77216 113892 77280
rect 113956 77216 113964 77280
rect 113644 76192 113964 77216
rect 113644 76128 113652 76192
rect 113716 76128 113732 76192
rect 113796 76128 113812 76192
rect 113876 76128 113892 76192
rect 113956 76128 113964 76192
rect 113644 75104 113964 76128
rect 113644 75040 113652 75104
rect 113716 75040 113732 75104
rect 113796 75040 113812 75104
rect 113876 75040 113892 75104
rect 113956 75040 113964 75104
rect 113644 74016 113964 75040
rect 113644 73952 113652 74016
rect 113716 73952 113732 74016
rect 113796 73952 113812 74016
rect 113876 73952 113892 74016
rect 113956 73952 113964 74016
rect 113644 72928 113964 73952
rect 113644 72864 113652 72928
rect 113716 72864 113732 72928
rect 113796 72864 113812 72928
rect 113876 72864 113892 72928
rect 113956 72864 113964 72928
rect 113644 71840 113964 72864
rect 113644 71776 113652 71840
rect 113716 71776 113732 71840
rect 113796 71776 113812 71840
rect 113876 71776 113892 71840
rect 113956 71776 113964 71840
rect 113644 70752 113964 71776
rect 113644 70688 113652 70752
rect 113716 70688 113732 70752
rect 113796 70688 113812 70752
rect 113876 70688 113892 70752
rect 113956 70688 113964 70752
rect 113644 69664 113964 70688
rect 113644 69600 113652 69664
rect 113716 69600 113732 69664
rect 113796 69600 113812 69664
rect 113876 69600 113892 69664
rect 113956 69600 113964 69664
rect 113644 68576 113964 69600
rect 113644 68512 113652 68576
rect 113716 68512 113732 68576
rect 113796 68512 113812 68576
rect 113876 68512 113892 68576
rect 113956 68512 113964 68576
rect 113644 67556 113964 68512
rect 113644 67488 113686 67556
rect 113922 67488 113964 67556
rect 113644 67424 113652 67488
rect 113956 67424 113964 67488
rect 113644 67320 113686 67424
rect 113922 67320 113964 67424
rect 113644 66400 113964 67320
rect 113644 66336 113652 66400
rect 113716 66336 113732 66400
rect 113796 66336 113812 66400
rect 113876 66336 113892 66400
rect 113956 66336 113964 66400
rect 113644 65312 113964 66336
rect 113644 65248 113652 65312
rect 113716 65248 113732 65312
rect 113796 65248 113812 65312
rect 113876 65248 113892 65312
rect 113956 65248 113964 65312
rect 113644 64224 113964 65248
rect 113644 64160 113652 64224
rect 113716 64160 113732 64224
rect 113796 64160 113812 64224
rect 113876 64160 113892 64224
rect 113956 64160 113964 64224
rect 113644 63136 113964 64160
rect 113644 63072 113652 63136
rect 113716 63072 113732 63136
rect 113796 63072 113812 63136
rect 113876 63072 113892 63136
rect 113956 63072 113964 63136
rect 113644 62048 113964 63072
rect 113644 61984 113652 62048
rect 113716 61984 113732 62048
rect 113796 61984 113812 62048
rect 113876 61984 113892 62048
rect 113956 61984 113964 62048
rect 113644 60960 113964 61984
rect 113644 60896 113652 60960
rect 113716 60896 113732 60960
rect 113796 60896 113812 60960
rect 113876 60896 113892 60960
rect 113956 60896 113964 60960
rect 113644 59872 113964 60896
rect 113644 59808 113652 59872
rect 113716 59808 113732 59872
rect 113796 59808 113812 59872
rect 113876 59808 113892 59872
rect 113956 59808 113964 59872
rect 113644 58784 113964 59808
rect 113644 58720 113652 58784
rect 113716 58720 113732 58784
rect 113796 58720 113812 58784
rect 113876 58720 113892 58784
rect 113956 58720 113964 58784
rect 113644 57696 113964 58720
rect 113644 57632 113652 57696
rect 113716 57632 113732 57696
rect 113796 57632 113812 57696
rect 113876 57632 113892 57696
rect 113956 57632 113964 57696
rect 113644 56608 113964 57632
rect 113644 56544 113652 56608
rect 113716 56544 113732 56608
rect 113796 56544 113812 56608
rect 113876 56544 113892 56608
rect 113956 56544 113964 56608
rect 113644 55520 113964 56544
rect 113644 55456 113652 55520
rect 113716 55456 113732 55520
rect 113796 55456 113812 55520
rect 113876 55456 113892 55520
rect 113956 55456 113964 55520
rect 113644 54432 113964 55456
rect 113644 54368 113652 54432
rect 113716 54368 113732 54432
rect 113796 54368 113812 54432
rect 113876 54368 113892 54432
rect 113956 54368 113964 54432
rect 113644 53344 113964 54368
rect 113644 53280 113652 53344
rect 113716 53280 113732 53344
rect 113796 53280 113812 53344
rect 113876 53280 113892 53344
rect 113956 53280 113964 53344
rect 113644 52256 113964 53280
rect 113644 52192 113652 52256
rect 113716 52192 113732 52256
rect 113796 52192 113812 52256
rect 113876 52192 113892 52256
rect 113956 52192 113964 52256
rect 113644 51168 113964 52192
rect 113644 51104 113652 51168
rect 113716 51104 113732 51168
rect 113796 51104 113812 51168
rect 113876 51104 113892 51168
rect 113956 51104 113964 51168
rect 113644 50080 113964 51104
rect 113644 50016 113652 50080
rect 113716 50016 113732 50080
rect 113796 50016 113812 50080
rect 113876 50016 113892 50080
rect 113956 50016 113964 50080
rect 113644 48992 113964 50016
rect 113644 48928 113652 48992
rect 113716 48928 113732 48992
rect 113796 48928 113812 48992
rect 113876 48928 113892 48992
rect 113956 48928 113964 48992
rect 113644 47904 113964 48928
rect 113644 47840 113652 47904
rect 113716 47840 113732 47904
rect 113796 47840 113812 47904
rect 113876 47840 113892 47904
rect 113956 47840 113964 47904
rect 113644 46816 113964 47840
rect 113644 46752 113652 46816
rect 113716 46752 113732 46816
rect 113796 46752 113812 46816
rect 113876 46752 113892 46816
rect 113956 46752 113964 46816
rect 113644 45728 113964 46752
rect 113644 45664 113652 45728
rect 113716 45664 113732 45728
rect 113796 45664 113812 45728
rect 113876 45664 113892 45728
rect 113956 45664 113964 45728
rect 113644 44640 113964 45664
rect 113644 44576 113652 44640
rect 113716 44576 113732 44640
rect 113796 44576 113812 44640
rect 113876 44576 113892 44640
rect 113956 44576 113964 44640
rect 113644 43552 113964 44576
rect 113644 43488 113652 43552
rect 113716 43488 113732 43552
rect 113796 43488 113812 43552
rect 113876 43488 113892 43552
rect 113956 43488 113964 43552
rect 113644 42464 113964 43488
rect 113644 42400 113652 42464
rect 113716 42400 113732 42464
rect 113796 42400 113812 42464
rect 113876 42400 113892 42464
rect 113956 42400 113964 42464
rect 113644 41376 113964 42400
rect 113644 41312 113652 41376
rect 113716 41312 113732 41376
rect 113796 41312 113812 41376
rect 113876 41312 113892 41376
rect 113956 41312 113964 41376
rect 113644 40288 113964 41312
rect 113644 40224 113652 40288
rect 113716 40224 113732 40288
rect 113796 40224 113812 40288
rect 113876 40224 113892 40288
rect 113956 40224 113964 40288
rect 113644 39200 113964 40224
rect 113644 39136 113652 39200
rect 113716 39136 113732 39200
rect 113796 39136 113812 39200
rect 113876 39136 113892 39200
rect 113956 39136 113964 39200
rect 113644 38112 113964 39136
rect 113644 38048 113652 38112
rect 113716 38048 113732 38112
rect 113796 38048 113812 38112
rect 113876 38048 113892 38112
rect 113956 38048 113964 38112
rect 113644 37024 113964 38048
rect 113644 36960 113652 37024
rect 113716 36960 113732 37024
rect 113796 36960 113812 37024
rect 113876 36960 113892 37024
rect 113956 36960 113964 37024
rect 113644 36920 113964 36960
rect 113644 36684 113686 36920
rect 113922 36684 113964 36920
rect 113644 35936 113964 36684
rect 113644 35872 113652 35936
rect 113716 35872 113732 35936
rect 113796 35872 113812 35936
rect 113876 35872 113892 35936
rect 113956 35872 113964 35936
rect 113644 34848 113964 35872
rect 113644 34784 113652 34848
rect 113716 34784 113732 34848
rect 113796 34784 113812 34848
rect 113876 34784 113892 34848
rect 113956 34784 113964 34848
rect 113644 33760 113964 34784
rect 113644 33696 113652 33760
rect 113716 33696 113732 33760
rect 113796 33696 113812 33760
rect 113876 33696 113892 33760
rect 113956 33696 113964 33760
rect 113644 32672 113964 33696
rect 113644 32608 113652 32672
rect 113716 32608 113732 32672
rect 113796 32608 113812 32672
rect 113876 32608 113892 32672
rect 113956 32608 113964 32672
rect 113644 31584 113964 32608
rect 113644 31520 113652 31584
rect 113716 31520 113732 31584
rect 113796 31520 113812 31584
rect 113876 31520 113892 31584
rect 113956 31520 113964 31584
rect 113644 30496 113964 31520
rect 113644 30432 113652 30496
rect 113716 30432 113732 30496
rect 113796 30432 113812 30496
rect 113876 30432 113892 30496
rect 113956 30432 113964 30496
rect 113644 29408 113964 30432
rect 113644 29344 113652 29408
rect 113716 29344 113732 29408
rect 113796 29344 113812 29408
rect 113876 29344 113892 29408
rect 113956 29344 113964 29408
rect 113644 28320 113964 29344
rect 113644 28256 113652 28320
rect 113716 28256 113732 28320
rect 113796 28256 113812 28320
rect 113876 28256 113892 28320
rect 113956 28256 113964 28320
rect 113644 27232 113964 28256
rect 113644 27168 113652 27232
rect 113716 27168 113732 27232
rect 113796 27168 113812 27232
rect 113876 27168 113892 27232
rect 113956 27168 113964 27232
rect 113644 26144 113964 27168
rect 113644 26080 113652 26144
rect 113716 26080 113732 26144
rect 113796 26080 113812 26144
rect 113876 26080 113892 26144
rect 113956 26080 113964 26144
rect 113644 25056 113964 26080
rect 113644 24992 113652 25056
rect 113716 24992 113732 25056
rect 113796 24992 113812 25056
rect 113876 24992 113892 25056
rect 113956 24992 113964 25056
rect 113644 23968 113964 24992
rect 113644 23904 113652 23968
rect 113716 23904 113732 23968
rect 113796 23904 113812 23968
rect 113876 23904 113892 23968
rect 113956 23904 113964 23968
rect 113644 22880 113964 23904
rect 113644 22816 113652 22880
rect 113716 22816 113732 22880
rect 113796 22816 113812 22880
rect 113876 22816 113892 22880
rect 113956 22816 113964 22880
rect 113644 21792 113964 22816
rect 113644 21728 113652 21792
rect 113716 21728 113732 21792
rect 113796 21728 113812 21792
rect 113876 21728 113892 21792
rect 113956 21728 113964 21792
rect 113644 20704 113964 21728
rect 113644 20640 113652 20704
rect 113716 20640 113732 20704
rect 113796 20640 113812 20704
rect 113876 20640 113892 20704
rect 113956 20640 113964 20704
rect 113644 19616 113964 20640
rect 113644 19552 113652 19616
rect 113716 19552 113732 19616
rect 113796 19552 113812 19616
rect 113876 19552 113892 19616
rect 113956 19552 113964 19616
rect 113644 18528 113964 19552
rect 113644 18464 113652 18528
rect 113716 18464 113732 18528
rect 113796 18464 113812 18528
rect 113876 18464 113892 18528
rect 113956 18464 113964 18528
rect 113644 17440 113964 18464
rect 113644 17376 113652 17440
rect 113716 17376 113732 17440
rect 113796 17376 113812 17440
rect 113876 17376 113892 17440
rect 113956 17376 113964 17440
rect 113644 16352 113964 17376
rect 113644 16288 113652 16352
rect 113716 16288 113732 16352
rect 113796 16288 113812 16352
rect 113876 16288 113892 16352
rect 113956 16288 113964 16352
rect 113644 15264 113964 16288
rect 113644 15200 113652 15264
rect 113716 15200 113732 15264
rect 113796 15200 113812 15264
rect 113876 15200 113892 15264
rect 113956 15200 113964 15264
rect 113644 14176 113964 15200
rect 113644 14112 113652 14176
rect 113716 14112 113732 14176
rect 113796 14112 113812 14176
rect 113876 14112 113892 14176
rect 113956 14112 113964 14176
rect 113644 13088 113964 14112
rect 113644 13024 113652 13088
rect 113716 13024 113732 13088
rect 113796 13024 113812 13088
rect 113876 13024 113892 13088
rect 113956 13024 113964 13088
rect 113644 12000 113964 13024
rect 113644 11936 113652 12000
rect 113716 11936 113732 12000
rect 113796 11936 113812 12000
rect 113876 11936 113892 12000
rect 113956 11936 113964 12000
rect 113644 10912 113964 11936
rect 113644 10848 113652 10912
rect 113716 10848 113732 10912
rect 113796 10848 113812 10912
rect 113876 10848 113892 10912
rect 113956 10848 113964 10912
rect 113644 9824 113964 10848
rect 113644 9760 113652 9824
rect 113716 9760 113732 9824
rect 113796 9760 113812 9824
rect 113876 9760 113892 9824
rect 113956 9760 113964 9824
rect 113644 8736 113964 9760
rect 113644 8672 113652 8736
rect 113716 8672 113732 8736
rect 113796 8672 113812 8736
rect 113876 8672 113892 8736
rect 113956 8672 113964 8736
rect 113644 7648 113964 8672
rect 113644 7584 113652 7648
rect 113716 7584 113732 7648
rect 113796 7584 113812 7648
rect 113876 7584 113892 7648
rect 113956 7584 113964 7648
rect 113644 7024 113964 7584
rect 97028 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97348 6560
rect 97028 6284 97348 6496
rect 97028 6048 97070 6284
rect 97306 6048 97348 6284
rect 97028 5472 97348 6048
rect 97028 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97348 5472
rect 97028 4384 97348 5408
rect 97028 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97348 4384
rect 97028 3296 97348 4320
rect 97028 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97348 3296
rect 97028 2208 97348 3232
rect 97028 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97348 2208
rect 97028 2128 97348 2144
<< via4 >>
rect 4250 94144 4486 94298
rect 4250 94080 4280 94144
rect 4280 94080 4296 94144
rect 4296 94080 4360 94144
rect 4360 94080 4376 94144
rect 4376 94080 4440 94144
rect 4440 94080 4456 94144
rect 4456 94080 4486 94144
rect 4250 94062 4486 94080
rect 4250 66880 4280 66896
rect 4280 66880 4296 66896
rect 4296 66880 4360 66896
rect 4360 66880 4376 66896
rect 4376 66880 4440 66896
rect 4440 66880 4456 66896
rect 4456 66880 4486 66896
rect 4250 66660 4486 66880
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 94742 5146 94978
rect 34970 94144 35206 94298
rect 34970 94080 35000 94144
rect 35000 94080 35016 94144
rect 35016 94080 35080 94144
rect 35080 94080 35096 94144
rect 35096 94080 35160 94144
rect 35160 94080 35176 94144
rect 35176 94080 35206 94144
rect 34970 94062 35206 94080
rect 35630 94742 35866 94978
rect 65690 94144 65926 94298
rect 65690 94080 65720 94144
rect 65720 94080 65736 94144
rect 65736 94080 65800 94144
rect 65800 94080 65816 94144
rect 65816 94080 65880 94144
rect 65880 94080 65896 94144
rect 65896 94080 65926 94144
rect 65690 94062 65926 94080
rect 66350 94742 66586 94978
rect 96410 94144 96646 94298
rect 96410 94080 96440 94144
rect 96440 94080 96456 94144
rect 96456 94080 96520 94144
rect 96520 94080 96536 94144
rect 96536 94080 96600 94144
rect 96600 94080 96616 94144
rect 96616 94080 96646 94144
rect 96410 94062 96646 94080
rect 97070 94742 97306 94978
rect 4910 67488 5146 67556
rect 4910 67424 4940 67488
rect 4940 67424 4956 67488
rect 4956 67424 5020 67488
rect 5020 67424 5036 67488
rect 5036 67424 5100 67488
rect 5100 67424 5116 67488
rect 5116 67424 5146 67488
rect 4910 67320 5146 67424
rect 10328 67320 10564 67556
rect 105392 67320 105628 67556
rect 11008 66660 11244 66896
rect 104712 66660 104948 66896
rect 112950 66880 112980 66896
rect 112980 66880 112996 66896
rect 112996 66880 113060 66896
rect 113060 66880 113076 66896
rect 113076 66880 113140 66896
rect 113140 66880 113156 66896
rect 113156 66880 113186 66896
rect 112950 66660 113186 66880
rect 4910 36684 5146 36920
rect 10328 36684 10564 36920
rect 105392 36684 105628 36920
rect 11008 36024 11244 36260
rect 104712 36024 104948 36260
rect 112950 36024 113186 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 6048 35866 6284
rect 65690 5388 65926 5624
rect 66350 6048 66586 6284
rect 96410 5388 96646 5624
rect 113686 67488 113922 67556
rect 113686 67424 113716 67488
rect 113716 67424 113732 67488
rect 113732 67424 113796 67488
rect 113796 67424 113812 67488
rect 113812 67424 113876 67488
rect 113876 67424 113892 67488
rect 113892 67424 113922 67488
rect 113686 67320 113922 67424
rect 113686 36684 113922 36920
rect 97070 6048 97306 6284
<< metal5 >>
rect 4208 94978 118912 95020
rect 4208 94742 4910 94978
rect 5146 94742 35630 94978
rect 35866 94742 66350 94978
rect 66586 94742 97070 94978
rect 97306 94742 118912 94978
rect 4208 94700 118912 94742
rect 4208 94298 118912 94340
rect 4208 94062 4250 94298
rect 4486 94062 34970 94298
rect 35206 94062 65690 94298
rect 65926 94062 96410 94298
rect 96646 94062 118912 94298
rect 4208 94020 118912 94062
rect 1056 67556 118912 67598
rect 1056 67320 4910 67556
rect 5146 67320 10328 67556
rect 10564 67320 105392 67556
rect 105628 67320 113686 67556
rect 113922 67320 118912 67556
rect 1056 67278 118912 67320
rect 1056 66896 118912 66938
rect 1056 66660 4250 66896
rect 4486 66660 11008 66896
rect 11244 66660 104712 66896
rect 104948 66660 112950 66896
rect 113186 66660 118912 66896
rect 1056 66618 118912 66660
rect 1056 36920 118912 36962
rect 1056 36684 4910 36920
rect 5146 36684 10328 36920
rect 10564 36684 105392 36920
rect 105628 36684 113686 36920
rect 113922 36684 118912 36920
rect 1056 36642 118912 36684
rect 1056 36260 118912 36302
rect 1056 36024 4250 36260
rect 4486 36024 11008 36260
rect 11244 36024 104712 36260
rect 104948 36024 112950 36260
rect 113186 36024 118912 36260
rect 1056 35982 118912 36024
rect 1056 6284 118912 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 66350 6284
rect 66586 6048 97070 6284
rect 97306 6048 118912 6284
rect 1056 6006 118912 6048
rect 1056 5624 118912 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 65690 5624
rect 65926 5388 96410 5624
rect 96646 5388 118912 5624
rect 1056 5346 118912 5388
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1
transform 1 0 118036 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1
transform -1 0 118312 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1
transform 1 0 117760 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1
transform 1 0 115368 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1
transform -1 0 114264 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1
transform 1 0 114816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _303_
timestamp 1
transform -1 0 115000 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1
transform -1 0 59524 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _305_
timestamp 1
transform 1 0 117392 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _306_
timestamp 1
transform 1 0 115828 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _307_
timestamp 1
transform -1 0 116564 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _308_
timestamp 1
transform -1 0 116840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _309_
timestamp 1
transform 1 0 116196 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _310_
timestamp 1
transform 1 0 115460 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _311_
timestamp 1
transform -1 0 117300 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _312_
timestamp 1
transform 1 0 116564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _313_
timestamp 1
transform -1 0 115460 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _314_
timestamp 1
transform -1 0 116564 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _315_
timestamp 1
transform -1 0 115184 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _316_
timestamp 1
transform -1 0 117668 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _317_
timestamp 1
transform 1 0 117668 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp 1
transform -1 0 118036 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _319_
timestamp 1
transform 1 0 117484 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _320_
timestamp 1
transform 1 0 117668 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _321_
timestamp 1
transform 1 0 117208 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _322_
timestamp 1
transform 1 0 117208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _323_
timestamp 1
transform -1 0 115736 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _324_
timestamp 1
transform -1 0 116288 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _325_
timestamp 1
transform 1 0 114724 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _326_
timestamp 1
transform 1 0 115092 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _327_
timestamp 1
transform -1 0 116380 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _328_
timestamp 1
transform -1 0 116932 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _329_
timestamp 1
transform -1 0 116932 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _330_
timestamp 1
transform -1 0 118128 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _331_
timestamp 1
transform 1 0 116932 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _332_
timestamp 1
transform -1 0 115092 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _333_
timestamp 1
transform 1 0 112976 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _334_
timestamp 1
transform 1 0 116104 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _335_
timestamp 1
transform -1 0 117024 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _336_
timestamp 1
transform -1 0 115828 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _337_
timestamp 1
transform 1 0 115828 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _338_
timestamp 1
transform -1 0 116196 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _339_
timestamp 1
transform -1 0 115828 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _340_
timestamp 1
transform -1 0 115552 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _341_
timestamp 1
transform -1 0 115368 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _342_
timestamp 1
transform 1 0 114448 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 1
transform -1 0 114448 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1
transform -1 0 112424 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _345_
timestamp 1
transform 1 0 113344 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1
transform 1 0 113436 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _347_
timestamp 1
transform -1 0 112332 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _348_
timestamp 1
transform 1 0 114816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _349_
timestamp 1
transform -1 0 115092 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _350_
timestamp 1
transform 1 0 113620 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _351_
timestamp 1
transform -1 0 112792 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _352_
timestamp 1
transform -1 0 111872 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _353_
timestamp 1
transform 1 0 114448 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _354_
timestamp 1
transform -1 0 114816 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _355_
timestamp 1
transform -1 0 112700 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _356_
timestamp 1
transform 1 0 113252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _357_
timestamp 1
transform -1 0 113252 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _358_
timestamp 1
transform -1 0 112424 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _359_
timestamp 1
transform 1 0 112056 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _360_
timestamp 1
transform 1 0 111780 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _361_
timestamp 1
transform 1 0 110768 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _362_
timestamp 1
transform -1 0 115736 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _363_
timestamp 1
transform -1 0 114172 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _364_
timestamp 1
transform -1 0 110492 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _365_
timestamp 1
transform 1 0 109388 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _366_
timestamp 1
transform 1 0 111228 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _367_
timestamp 1
transform 1 0 111136 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _368_
timestamp 1
transform 1 0 109572 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _369_
timestamp 1
transform 1 0 110216 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _370_
timestamp 1
transform 1 0 110676 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _371_
timestamp 1
transform 1 0 109756 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _372_
timestamp 1
transform -1 0 110216 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _373_
timestamp 1
transform 1 0 110676 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _374_
timestamp 1
transform -1 0 110308 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _375_
timestamp 1
transform -1 0 112332 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _376_
timestamp 1
transform 1 0 110216 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _377_
timestamp 1
transform -1 0 111596 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _378_
timestamp 1
transform 1 0 109664 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _379_
timestamp 1
transform 1 0 109296 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1
transform 1 0 109664 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _381_
timestamp 1
transform -1 0 110492 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _382_
timestamp 1
transform -1 0 111320 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _383_
timestamp 1
transform -1 0 109756 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _384_
timestamp 1
transform 1 0 111596 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _385_
timestamp 1
transform 1 0 111136 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _386_
timestamp 1
transform -1 0 111136 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _387_
timestamp 1
transform -1 0 112332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1
transform 1 0 113160 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _389_
timestamp 1
transform 1 0 109020 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1
transform -1 0 111044 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _391_
timestamp 1
transform 1 0 112792 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _392_
timestamp 1
transform -1 0 111964 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _393_
timestamp 1
transform -1 0 111596 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _394_
timestamp 1
transform 1 0 110952 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _395_
timestamp 1
transform -1 0 111596 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _396_
timestamp 1
transform 1 0 112700 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _397_
timestamp 1
transform -1 0 112148 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _398_
timestamp 1
transform 1 0 112148 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _399_
timestamp 1
transform 1 0 112332 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _400_
timestamp 1
transform 1 0 114356 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _401_
timestamp 1
transform 1 0 113252 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _402_
timestamp 1
transform -1 0 113620 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _403_
timestamp 1
transform 1 0 111688 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1
transform -1 0 112976 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _405_
timestamp 1
transform 1 0 112516 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _406_
timestamp 1
transform 1 0 112792 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _407_
timestamp 1
transform -1 0 114908 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _408_
timestamp 1
transform 1 0 113712 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1
transform 1 0 114540 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _410_
timestamp 1
transform 1 0 113252 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _411_
timestamp 1
transform 1 0 111688 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _412_
timestamp 1
transform 1 0 113804 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _413_
timestamp 1
transform 1 0 111780 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _414_
timestamp 1
transform 1 0 112424 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _415_
timestamp 1
transform -1 0 114264 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _416_
timestamp 1
transform -1 0 116656 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _417_
timestamp 1
transform -1 0 116196 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_2  _418_
timestamp 1
transform 1 0 113436 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _419_
timestamp 1
transform 1 0 112240 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _420_
timestamp 1
transform 1 0 113252 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _421_
timestamp 1
transform -1 0 114540 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _422_
timestamp 1
transform -1 0 116748 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _423_
timestamp 1
transform 1 0 115828 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _424_
timestamp 1
transform 1 0 115460 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _425_
timestamp 1
transform -1 0 117760 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _426_
timestamp 1
transform 1 0 116564 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _427_
timestamp 1
transform 1 0 115184 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _428_
timestamp 1
transform -1 0 117852 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _429_
timestamp 1
transform -1 0 117668 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1
transform -1 0 117484 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _431_
timestamp 1
transform 1 0 117760 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _432_
timestamp 1
transform 1 0 117484 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _433_
timestamp 1
transform -1 0 116472 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1
transform 1 0 115000 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _435_
timestamp 1
transform 1 0 115552 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _436_
timestamp 1
transform -1 0 115644 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _437_
timestamp 1
transform 1 0 117300 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _438_
timestamp 1
transform -1 0 116288 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _439_
timestamp 1
transform -1 0 117300 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _440_
timestamp 1
transform 1 0 118128 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _441_
timestamp 1
transform 1 0 117760 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _442_
timestamp 1
transform -1 0 118312 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1
transform -1 0 117760 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _444_
timestamp 1
transform 1 0 117024 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _445_
timestamp 1
transform 1 0 115460 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _446_
timestamp 1
transform 1 0 116012 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1
transform -1 0 117024 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _448_
timestamp 1
transform 1 0 116288 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _449_
timestamp 1
transform -1 0 116104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _450_
timestamp 1
transform 1 0 114632 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _451_
timestamp 1
transform -1 0 115184 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _452_
timestamp 1
transform 1 0 115184 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _453_
timestamp 1
transform 1 0 114632 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _454_
timestamp 1
transform 1 0 115460 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _455_
timestamp 1
transform 1 0 113528 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _456_
timestamp 1
transform 1 0 113988 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _457_
timestamp 1
transform -1 0 115000 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _458_
timestamp 1
transform 1 0 116932 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _459_
timestamp 1
transform -1 0 117024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _460_
timestamp 1
transform 1 0 117944 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _461_
timestamp 1
transform 1 0 117392 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _462_
timestamp 1
transform -1 0 116104 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _463_
timestamp 1
transform 1 0 116104 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _464_
timestamp 1
transform -1 0 115644 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _465_
timestamp 1
transform 1 0 114172 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1
transform 1 0 114448 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _467_
timestamp 1
transform 1 0 115000 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _468_
timestamp 1
transform 1 0 115000 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _469_
timestamp 1
transform -1 0 113988 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _470_
timestamp 1
transform 1 0 113252 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _471_
timestamp 1
transform 1 0 112884 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _472_
timestamp 1
transform -1 0 115460 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_2  _473_
timestamp 1
transform 1 0 112516 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _474_
timestamp 1
transform 1 0 115644 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 1
transform 1 0 115828 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1
transform -1 0 114632 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _477_
timestamp 1
transform -1 0 115368 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _478_
timestamp 1
transform -1 0 114724 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__a311o_1  _479_
timestamp 1
transform 1 0 113344 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _480_
timestamp 1
transform -1 0 113252 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _481_
timestamp 1
transform 1 0 114080 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _482_
timestamp 1
transform 1 0 113344 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _483_
timestamp 1
transform 1 0 111136 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _484_
timestamp 1
transform 1 0 111320 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp 1
transform -1 0 112884 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _486_
timestamp 1
transform 1 0 112240 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _487_
timestamp 1
transform -1 0 112516 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _488_
timestamp 1
transform 1 0 113436 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _489_
timestamp 1
transform 1 0 113988 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _490_
timestamp 1
transform -1 0 115000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _491_
timestamp 1
transform 1 0 113252 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _492_
timestamp 1
transform -1 0 112148 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _493_
timestamp 1
transform -1 0 112884 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _494_
timestamp 1
transform -1 0 111228 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _495_
timestamp 1
transform -1 0 112056 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _496_
timestamp 1
transform -1 0 111136 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _497_
timestamp 1
transform -1 0 110032 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _498_
timestamp 1
transform 1 0 108652 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _499_
timestamp 1
transform 1 0 111136 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _500_
timestamp 1
transform 1 0 109480 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _501_
timestamp 1
transform -1 0 110584 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _502_
timestamp 1
transform 1 0 108744 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _503_
timestamp 1
transform 1 0 109572 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _504_
timestamp 1
transform 1 0 110216 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _505_
timestamp 1
transform -1 0 111320 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _506_
timestamp 1
transform -1 0 112148 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _507_
timestamp 1
transform 1 0 109756 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _508_
timestamp 1
transform 1 0 112056 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _509_
timestamp 1
transform -1 0 111596 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _510_
timestamp 1
transform -1 0 111320 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _511_
timestamp 1
transform 1 0 110676 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _512_
timestamp 1
transform -1 0 111136 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _513_
timestamp 1
transform 1 0 110584 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _514_
timestamp 1
transform 1 0 110492 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _515_
timestamp 1
transform -1 0 111228 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _516_
timestamp 1
transform -1 0 111228 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _517_
timestamp 1
transform -1 0 111228 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _518_
timestamp 1
transform -1 0 109940 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _519_
timestamp 1
transform 1 0 109940 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _520_
timestamp 1
transform -1 0 110768 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _521_
timestamp 1
transform -1 0 109480 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _522_
timestamp 1
transform 1 0 110400 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _523_
timestamp 1
transform -1 0 109664 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _524_
timestamp 1
transform -1 0 109480 0 -1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _525_
timestamp 1
transform 1 0 109296 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _526_
timestamp 1
transform -1 0 109940 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _527_
timestamp 1
transform 1 0 110032 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _528_
timestamp 1
transform -1 0 109940 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _529_
timestamp 1
transform 1 0 110216 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _530_
timestamp 1
transform -1 0 110032 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _531_
timestamp 1
transform -1 0 110584 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _532_
timestamp 1
transform 1 0 108560 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _533_
timestamp 1
transform -1 0 109756 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _534_
timestamp 1
transform -1 0 109572 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _535_
timestamp 1
transform 1 0 108284 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _536_
timestamp 1
transform -1 0 109388 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _537_
timestamp 1
transform -1 0 108836 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _538_
timestamp 1
transform 1 0 108836 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _539_
timestamp 1
transform -1 0 109020 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _540_
timestamp 1
transform -1 0 109572 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _541_
timestamp 1
transform 1 0 108836 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _542_
timestamp 1
transform 1 0 109112 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _543_
timestamp 1
transform 1 0 108468 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _544_
timestamp 1
transform 1 0 108468 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _545_
timestamp 1
transform 1 0 109112 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _546_
timestamp 1
transform 1 0 109480 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _547_
timestamp 1
transform -1 0 110032 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _548_
timestamp 1
transform -1 0 54556 0 -1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _549_
timestamp 1
transform -1 0 55384 0 -1 94656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _550_
timestamp 1
transform -1 0 56764 0 1 94656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _551_
timestamp 1
transform -1 0 57776 0 -1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _552_
timestamp 1
transform -1 0 58880 0 -1 94656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1
transform -1 0 60076 0 1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _554_
timestamp 1
transform -1 0 61272 0 1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1
transform -1 0 62192 0 1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _556_
timestamp 1
transform -1 0 63020 0 1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1
transform -1 0 64216 0 1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _558_
timestamp 1
transform -1 0 65136 0 1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1
transform -1 0 66424 0 1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _560_
timestamp 1
transform -1 0 67160 0 -1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _561_
timestamp 1
transform -1 0 69000 0 -1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _562_
timestamp 1
transform -1 0 69828 0 -1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _563_
timestamp 1
transform -1 0 70748 0 -1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _564_
timestamp 1
transform -1 0 60352 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _565_
timestamp 1
transform -1 0 61916 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _566_
timestamp 1
transform -1 0 63296 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _567_
timestamp 1
transform -1 0 63388 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _568_
timestamp 1
transform -1 0 65412 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp 1
transform -1 0 65504 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _570_
timestamp 1
transform -1 0 66700 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _571_
timestamp 1
transform -1 0 67252 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _572_
timestamp 1
transform 1 0 68724 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _573_
timestamp 1
transform -1 0 69276 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _574_
timestamp 1
transform -1 0 70104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1
transform -1 0 71024 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _576_
timestamp 1
transform 1 0 72588 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1
transform -1 0 73140 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _578_
timestamp 1
transform -1 0 74888 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _579_
timestamp 1
transform 1 0 108284 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1
transform 1 0 108836 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1
transform 1 0 108284 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1
transform 1 0 108284 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1
transform 1 0 108284 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _584_
timestamp 1
transform 1 0 108284 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _585_
timestamp 1
transform 1 0 108284 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1
transform 1 0 108376 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _587_
timestamp 1
transform 1 0 108284 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _588_
timestamp 1
transform 1 0 55660 0 -1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _589_
timestamp 1
transform 1 0 56764 0 1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _590_
timestamp 1
transform 1 0 57868 0 1 94656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _591_
timestamp 1
transform 1 0 59248 0 -1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _592_
timestamp 1
transform 1 0 59524 0 -1 94656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _593_
timestamp 1
transform 1 0 61088 0 -1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _594_
timestamp 1
transform 1 0 62008 0 1 94656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _595_
timestamp 1
transform 1 0 63204 0 -1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _596_
timestamp 1
transform 1 0 65044 0 -1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _597_
timestamp 1
transform 1 0 65596 0 1 94656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _598_
timestamp 1
transform 1 0 66056 0 1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _599_
timestamp 1
transform 1 0 67436 0 1 94656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _600_
timestamp 1
transform 1 0 68172 0 -1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _601_
timestamp 1
transform 1 0 70012 0 -1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _602_
timestamp 1
transform 1 0 70748 0 1 94656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _603_
timestamp 1
transform 1 0 71668 0 1 95744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _604_
timestamp 1
transform 1 0 108284 0 1 52224
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _605_
timestamp 1
transform -1 0 110400 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _606_
timestamp 1
transform -1 0 110492 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _607_
timestamp 1
transform -1 0 110400 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _608_
timestamp 1
transform 1 0 108284 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _609_
timestamp 1
transform -1 0 110124 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _610_
timestamp 1
transform -1 0 110308 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _611_
timestamp 1
transform -1 0 110400 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _612_
timestamp 1
transform -1 0 110492 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _613_
timestamp 1
transform 1 0 45540 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _614_
timestamp 1
transform 1 0 47012 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _615_
timestamp 1
transform 1 0 48208 0 -1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _616_
timestamp 1
transform 1 0 49496 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _617_
timestamp 1
transform 1 0 50416 0 -1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _618_
timestamp 1
transform 1 0 50784 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _619_
timestamp 1
transform 1 0 52256 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _620_
timestamp 1
transform 1 0 53360 0 -1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _621_
timestamp 1
transform 1 0 53728 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _622_
timestamp 1
transform 1 0 55568 0 -1 94656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _623_
timestamp 1
transform 1 0 56304 0 -1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _624_
timestamp 1
transform 1 0 58144 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _625_
timestamp 1
transform 1 0 58880 0 -1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _626_
timestamp 1
transform 1 0 60720 0 -1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _627_
timestamp 1
transform 1 0 61916 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _628_
timestamp 1
transform 1 0 63572 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _629_
timestamp 1
transform -1 0 57224 0 1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _630_
timestamp 1
transform -1 0 57960 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _631_
timestamp 1
transform -1 0 59248 0 1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _632_
timestamp 1
transform -1 0 59984 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _633_
timestamp 1
transform -1 0 61456 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _634_
timestamp 1
transform -1 0 62928 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _635_
timestamp 1
transform -1 0 64860 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _636_
timestamp 1
transform -1 0 66332 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _637_
timestamp 1
transform -1 0 67068 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _638_
timestamp 1
transform -1 0 68540 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _639_
timestamp 1
transform -1 0 70012 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _640_
timestamp 1
transform -1 0 69736 0 -1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _641_
timestamp 1
transform -1 0 72220 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _642_
timestamp 1
transform -1 0 72220 0 -1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _643_
timestamp 1
transform -1 0 73692 0 1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _644_
timestamp 1
transform -1 0 74796 0 -1 92480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _645_
timestamp 1
transform -1 0 109848 0 -1 67456
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _646_
timestamp 1
transform 1 0 108284 0 1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform -1 0 45540 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 56120 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform -1 0 58144 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform 1 0 58696 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform 1 0 60536 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform -1 0 61916 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform -1 0 63572 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform -1 0 48668 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform 1 0 48024 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform 1 0 49312 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform 1 0 50232 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform -1 0 50784 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform -1 0 55476 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform 1 0 53176 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform -1 0 55660 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform 1 0 55384 0 -1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform 1 0 55568 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__A1
timestamp 1
transform 1 0 110400 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__A
timestamp 1
transform -1 0 110768 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1
transform 1 0 109296 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__A
timestamp 1
transform -1 0 73692 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A
timestamp 1
transform 1 0 74888 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__A
timestamp 1
transform 1 0 108560 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__A
timestamp 1
transform -1 0 109296 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__581__A
timestamp 1
transform 1 0 108560 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__A
timestamp 1
transform 1 0 108284 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A
timestamp 1
transform 1 0 108560 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__A
timestamp 1
transform 1 0 108560 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__585__A
timestamp 1
transform 1 0 108560 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__A
timestamp 1
transform 1 0 108652 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__587__A
timestamp 1
transform 1 0 108560 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__CLK
timestamp 1
transform 1 0 110400 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__CLK
timestamp 1
transform -1 0 110308 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__CLK
timestamp 1
transform -1 0 110860 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__Q
timestamp 1
transform 1 0 110676 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__CLK
timestamp 1
transform 1 0 47012 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__614__CLK
timestamp 1
transform 1 0 46828 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__615__CLK
timestamp 1
transform 1 0 47840 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__CLK
timestamp 1
transform 1 0 49128 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__617__CLK
timestamp 1
transform 1 0 49864 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__CLK
timestamp 1
transform 1 0 72864 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__CLK
timestamp 1
transform -1 0 72404 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__CLK
timestamp 1
transform 1 0 73692 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__CLK
timestamp 1
transform 1 0 74796 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__CLK
timestamp 1
transform 1 0 110032 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__Q
timestamp 1
transform -1 0 110032 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__CLK
timestamp 1
transform 1 0 109940 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__D
timestamp 1
transform -1 0 109940 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1
transform -1 0 65412 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 1
transform 1 0 65044 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_clk_A
timestamp 1
transform 1 0 47012 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_clk_X
timestamp 1
transform 1 0 47196 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_clk_A
timestamp 1
transform 1 0 56488 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_clk_A
timestamp 1
transform -1 0 58420 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_clk_A
timestamp 1
transform -1 0 67712 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_clk_A
timestamp 1
transform -1 0 108468 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_clk_X
timestamp 1
transform 1 0 110124 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_clk_A
timestamp 1
transform -1 0 108468 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_clk_A
timestamp 1
transform 1 0 70840 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_clk_A
timestamp 1
transform 1 0 77280 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_clk_X
timestamp 1
transform 1 0 79304 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 1
transform 1 0 46184 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload3_A
timestamp 1
transform 1 0 108928 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload6_A
timestamp 1
transform 1 0 77832 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout76_A
timestamp 1
transform 1 0 64308 0 -1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout77_A
timestamp 1
transform 1 0 71024 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1
transform -1 0 73508 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1
transform -1 0 75256 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_X
timestamp 1
transform 1 0 75256 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1
transform -1 0 25852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1
transform -1 0 1840 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1
transform -1 0 1840 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1
transform -1 0 1840 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1
transform -1 0 1840 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1
transform -1 0 1840 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1
transform -1 0 1840 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1
transform -1 0 1840 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1
transform -1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1
transform 1 0 118404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1
transform -1 0 118312 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1
transform -1 0 117208 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1
transform -1 0 118588 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1
transform -1 0 43240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1
transform -1 0 44528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1
transform -1 0 45816 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1
transform -1 0 46460 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1
transform -1 0 47748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1
transform -1 0 49036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1
transform -1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1
transform -1 0 33580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1
transform -1 0 34868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1
transform -1 0 36156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1
transform -1 0 37444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1
transform -1 0 38088 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1
transform -1 0 40020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1
transform -1 0 40664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1
transform -1 0 50324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1
transform -1 0 61916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1
transform -1 0 63204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1
transform -1 0 63848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1
transform -1 0 65136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1
transform -1 0 66424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1
transform -1 0 67712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1
transform -1 0 51612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1
transform -1 0 52256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1
transform -1 0 53544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1
transform -1 0 54832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1
transform -1 0 56120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1
transform -1 0 57408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1
transform -1 0 58052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1
transform -1 0 59340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1
transform -1 0 60628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1
transform -1 0 118588 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1
transform -1 0 118312 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1
transform -1 0 118588 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1
transform -1 0 118588 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1
transform -1 0 107640 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_X
timestamp 1
transform -1 0 108192 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew78_X
timestamp 1
transform -1 0 109388 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew80_X
timestamp 1
transform -1 0 109572 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew83_X
timestamp 1
transform -1 0 109204 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew86_X
timestamp 1
transform -1 0 110216 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_load_slew101_X
timestamp 1
transform -1 0 109756 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[0]
timestamp 1
transform -1 0 89608 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[4]
timestamp 1
transform -1 0 93472 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[5]
timestamp 1
transform -1 0 92920 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[6]
timestamp 1
transform -1 0 93104 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[7]
timestamp 1
transform -1 0 93288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_clk0
timestamp 1
transform -1 0 16100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_clk1
timestamp 1
transform -1 0 100280 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 65044 0 -1 92480
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1
transform -1 0 47012 0 -1 92480
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1
transform 1 0 54648 0 -1 93568
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1
transform -1 0 57684 0 1 96832
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1
transform -1 0 70012 0 1 96832
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1
transform 1 0 108284 0 1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1
transform 1 0 108284 0 1 51136
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1
transform -1 0 72864 0 -1 92480
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1
transform 1 0 77464 0 1 92480
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 1
transform -1 0 46184 0 -1 93568
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  clkload1
timestamp 1
transform 1 0 54648 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 1
transform -1 0 56396 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload3
timestamp 1
transform 1 0 108284 0 -1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload4
timestamp 1
transform -1 0 108836 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload5
timestamp 1
transform 1 0 70288 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  clkload6
timestamp 1
transform 1 0 77464 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  clone1
timestamp 1
transform -1 0 110492 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 1
transform -1 0 117392 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout76
timestamp 1
transform -1 0 64308 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout77
timestamp 1
transform -1 0 70656 0 1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout102
timestamp 1
transform -1 0 68724 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout103
timestamp 1
transform -1 0 72588 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout104
timestamp 1
transform 1 0 73784 0 -1 93568
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout105
timestamp 1
transform 1 0 116840 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp 1
transform 1 0 116472 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp 1
transform -1 0 117208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 1
transform 1 0 117116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 1
transform -1 0 116564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout110
timestamp 1
transform -1 0 116840 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout111
timestamp 1
transform -1 0 118404 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout112
timestamp 1
transform -1 0 118036 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_265
timestamp 1
transform 1 0 25484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636968456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_321
timestamp 1
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_329
timestamp 1
transform 1 0 31372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_343
timestamp 1
transform 1 0 32660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_349
timestamp 1
transform 1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_370
timestamp 1
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_378
timestamp 1
transform 1 0 35880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_398
timestamp 1
transform 1 0 37720 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636968456
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_426
timestamp 1
transform 1 0 40296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_433
timestamp 1
transform 1 0 40940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_441
timestamp 1
transform 1 0 41676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_449
timestamp 1
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_455
timestamp 1
transform 1 0 42964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_461
timestamp 1
transform 1 0 43516 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_469
timestamp 1
transform 1 0 44252 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_477
timestamp 1
transform 1 0 44988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_483
timestamp 1
transform 1 0 45540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_489
timestamp 1
transform 1 0 46092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_496
timestamp 1
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_510
timestamp 1
transform 1 0 48024 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_518
timestamp 1
transform 1 0 48760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_524
timestamp 1
transform 1 0 49312 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_538
timestamp 1
transform 1 0 50600 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_546
timestamp 1
transform 1 0 51336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_552
timestamp 1
transform 1 0 51888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_561
timestamp 1
transform 1 0 52716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_567
timestamp 1
transform 1 0 53268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_573
timestamp 1
transform 1 0 53820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_581
timestamp 1
transform 1 0 54556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_589
timestamp 1
transform 1 0 55292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_595
timestamp 1
transform 1 0 55844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_601
timestamp 1
transform 1 0 56396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_609
timestamp 1
transform 1 0 57132 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_622
timestamp 1
transform 1 0 58328 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_630
timestamp 1
transform 1 0 59064 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_636
timestamp 1
transform 1 0 59616 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_650
timestamp 1
transform 1 0 60904 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_658
timestamp 1
transform 1 0 61640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_664
timestamp 1
transform 1 0 62192 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_678
timestamp 1
transform 1 0 63480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_685
timestamp 1
transform 1 0 64124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_693
timestamp 1
transform 1 0 64860 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_701
timestamp 1
transform 1 0 65596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_707
timestamp 1
transform 1 0 66148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_713
timestamp 1
transform 1 0 66700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_721
timestamp 1
transform 1 0 67436 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_727
timestamp 1
transform 1 0 67988 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1636968456
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1636968456
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1636968456
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1636968456
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1636968456
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1636968456
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1636968456
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1636968456
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1636968456
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1636968456
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1636968456
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1636968456
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1636968456
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1636968456
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1636968456
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1636968456
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1636968456
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1636968456
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1636968456
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1636968456
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1636968456
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1636968456
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1636968456
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1636968456
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1636968456
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1636968456
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1636968456
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1636968456
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1636968456
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1636968456
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1636968456
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1161
timestamp 1636968456
transform 1 0 107916 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1173
timestamp 1
transform 1 0 109020 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1177
timestamp 1636968456
transform 1 0 109388 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1189
timestamp 1636968456
transform 1 0 110492 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1201
timestamp 1
transform 1 0 111596 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1205
timestamp 1636968456
transform 1 0 111964 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1217
timestamp 1636968456
transform 1 0 113068 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1229
timestamp 1
transform 1 0 114172 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1233
timestamp 1636968456
transform 1 0 114540 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1245
timestamp 1636968456
transform 1 0 115644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1257
timestamp 1
transform 1 0 116748 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1261
timestamp 1636968456
transform 1 0 117116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1273
timestamp 1
transform 1 0 118220 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636968456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636968456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636968456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636968456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636968456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636968456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636968456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636968456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636968456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636968456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636968456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636968456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636968456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636968456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636968456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636968456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636968456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636968456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636968456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636968456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636968456
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636968456
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636968456
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636968456
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636968456
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636968456
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636968456
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636968456
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636968456
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636968456
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636968456
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636968456
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636968456
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636968456
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636968456
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636968456
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636968456
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636968456
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636968456
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636968456
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1636968456
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1636968456
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1636968456
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1636968456
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1636968456
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1636968456
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1636968456
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1636968456
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1636968456
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1636968456
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1636968456
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1636968456
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1636968456
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1636968456
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1636968456
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1636968456
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1636968456
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1636968456
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1636968456
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1157
timestamp 1636968456
transform 1 0 107548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1
transform 1 0 108652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1177
timestamp 1636968456
transform 1 0 109388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1189
timestamp 1636968456
transform 1 0 110492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1201
timestamp 1636968456
transform 1 0 111596 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1213
timestamp 1636968456
transform 1 0 112700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1225
timestamp 1
transform 1 0 113804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1233
timestamp 1636968456
transform 1 0 114540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1245
timestamp 1636968456
transform 1 0 115644 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1257
timestamp 1636968456
transform 1 0 116748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1269
timestamp 1
transform 1 0 117852 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636968456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636968456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636968456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636968456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636968456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636968456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636968456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636968456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636968456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636968456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636968456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636968456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636968456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636968456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636968456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636968456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636968456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636968456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636968456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636968456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636968456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636968456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636968456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636968456
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636968456
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636968456
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636968456
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636968456
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636968456
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636968456
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636968456
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636968456
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636968456
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636968456
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636968456
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636968456
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636968456
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636968456
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636968456
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636968456
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636968456
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636968456
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636968456
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1636968456
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1636968456
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1636968456
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1636968456
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1636968456
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1636968456
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1636968456
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1636968456
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1636968456
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1636968456
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1636968456
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1636968456
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1636968456
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1636968456
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1636968456
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1636968456
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1636968456
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1636968456
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1636968456
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1636968456
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1185
timestamp 1636968456
transform 1 0 110124 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1197
timestamp 1
transform 1 0 111228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1203
timestamp 1
transform 1 0 111780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1205
timestamp 1636968456
transform 1 0 111964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1217
timestamp 1636968456
transform 1 0 113068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1229
timestamp 1636968456
transform 1 0 114172 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1241
timestamp 1636968456
transform 1 0 115276 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1253
timestamp 1
transform 1 0 116380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1
transform 1 0 116932 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1261
timestamp 1636968456
transform 1 0 117116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1273
timestamp 1
transform 1 0 118220 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636968456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636968456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636968456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636968456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636968456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636968456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636968456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636968456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636968456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636968456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636968456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636968456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636968456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636968456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636968456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636968456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636968456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636968456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636968456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636968456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636968456
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636968456
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636968456
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636968456
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636968456
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636968456
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636968456
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636968456
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636968456
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636968456
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636968456
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636968456
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636968456
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636968456
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636968456
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636968456
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636968456
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636968456
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636968456
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636968456
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1636968456
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1636968456
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1636968456
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1636968456
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1636968456
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1636968456
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1636968456
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1636968456
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1636968456
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1636968456
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1636968456
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1636968456
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1636968456
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1636968456
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1636968456
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1636968456
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1636968456
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1636968456
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1636968456
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1636968456
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1636968456
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1189
timestamp 1636968456
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1201
timestamp 1636968456
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1213
timestamp 1636968456
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1233
timestamp 1636968456
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1245
timestamp 1636968456
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1257
timestamp 1636968456
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1269
timestamp 1
transform 1 0 117852 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636968456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636968456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636968456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636968456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636968456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636968456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636968456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636968456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636968456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636968456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636968456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636968456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636968456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636968456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636968456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636968456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636968456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636968456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636968456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636968456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636968456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636968456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636968456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636968456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636968456
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636968456
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636968456
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636968456
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636968456
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636968456
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636968456
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636968456
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636968456
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636968456
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636968456
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636968456
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636968456
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636968456
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636968456
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1636968456
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1636968456
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636968456
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636968456
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1636968456
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1636968456
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1636968456
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1636968456
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1636968456
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1636968456
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1636968456
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1636968456
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1636968456
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1636968456
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1636968456
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1636968456
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1636968456
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1636968456
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1636968456
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1636968456
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1636968456
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1636968456
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1636968456
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1636968456
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1636968456
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1185
timestamp 1636968456
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1205
timestamp 1636968456
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1217
timestamp 1636968456
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1229
timestamp 1636968456
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1241
timestamp 1636968456
transform 1 0 115276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1253
timestamp 1
transform 1 0 116380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1261
timestamp 1636968456
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1273
timestamp 1
transform 1 0 118220 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636968456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636968456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636968456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636968456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636968456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636968456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636968456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636968456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636968456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636968456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636968456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636968456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636968456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636968456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636968456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636968456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636968456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636968456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636968456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636968456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636968456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636968456
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636968456
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636968456
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636968456
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636968456
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636968456
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636968456
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636968456
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636968456
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636968456
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636968456
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636968456
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636968456
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636968456
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1636968456
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1636968456
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1636968456
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1636968456
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1636968456
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636968456
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1636968456
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1636968456
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1636968456
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1636968456
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1636968456
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1636968456
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1636968456
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1636968456
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1636968456
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1636968456
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1636968456
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1636968456
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1636968456
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1636968456
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1636968456
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1636968456
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1636968456
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1636968456
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1636968456
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1636968456
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1636968456
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1189
timestamp 1636968456
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1201
timestamp 1636968456
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1213
timestamp 1636968456
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1233
timestamp 1636968456
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1245
timestamp 1636968456
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1257
timestamp 1636968456
transform 1 0 116748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1269
timestamp 1
transform 1 0 117852 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636968456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636968456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636968456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636968456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636968456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636968456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636968456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636968456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636968456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636968456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636968456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636968456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636968456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636968456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636968456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1636968456
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1636968456
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636968456
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636968456
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1636968456
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1636968456
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636968456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636968456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1636968456
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1636968456
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636968456
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636968456
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1636968456
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1636968456
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636968456
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636968456
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1636968456
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1636968456
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636968456
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636968456
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1636968456
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1636968456
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1636968456
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1636968456
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1636968456
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1636968456
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1636968456
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1636968456
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1636968456
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1636968456
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1636968456
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1636968456
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1636968456
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1636968456
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1636968456
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1636968456
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1636968456
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1636968456
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1636968456
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1636968456
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1636968456
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1636968456
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1636968456
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1636968456
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1636968456
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1636968456
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1636968456
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1636968456
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1636968456
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1185
timestamp 1636968456
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1205
timestamp 1636968456
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1217
timestamp 1636968456
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1229
timestamp 1636968456
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1241
timestamp 1636968456
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1261
timestamp 1636968456
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1273
timestamp 1
transform 1 0 118220 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636968456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636968456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636968456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636968456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636968456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636968456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636968456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636968456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636968456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636968456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636968456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636968456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636968456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636968456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636968456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636968456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1636968456
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1636968456
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1636968456
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636968456
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636968456
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636968456
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636968456
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1636968456
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1636968456
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1636968456
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1636968456
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1636968456
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1636968456
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1636968456
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1636968456
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1636968456
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1636968456
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1636968456
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1636968456
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1636968456
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1636968456
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1636968456
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1636968456
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1636968456
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1636968456
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1636968456
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1636968456
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1636968456
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1636968456
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1636968456
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1636968456
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1636968456
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1636968456
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1636968456
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1636968456
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1636968456
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1636968456
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1636968456
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1636968456
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1636968456
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1636968456
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1636968456
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1636968456
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1636968456
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1636968456
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1636968456
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1636968456
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1636968456
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1636968456
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1636968456
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1636968456
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1636968456
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1189
timestamp 1636968456
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1201
timestamp 1636968456
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1213
timestamp 1636968456
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1233
timestamp 1636968456
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1245
timestamp 1636968456
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1257
timestamp 1636968456
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1269
timestamp 1
transform 1 0 117852 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636968456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636968456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636968456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636968456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636968456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636968456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636968456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636968456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636968456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636968456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636968456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636968456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636968456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636968456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636968456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636968456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636968456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636968456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636968456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636968456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636968456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636968456
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636968456
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636968456
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636968456
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636968456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636968456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1636968456
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1636968456
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1636968456
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1636968456
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1636968456
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1636968456
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1636968456
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1636968456
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1636968456
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1636968456
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1636968456
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1636968456
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1636968456
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1636968456
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1636968456
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1636968456
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1636968456
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1636968456
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1636968456
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1636968456
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1636968456
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1636968456
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1636968456
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1636968456
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1636968456
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1636968456
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1636968456
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1636968456
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1636968456
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1636968456
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1636968456
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1636968456
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1636968456
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1636968456
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1636968456
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1636968456
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1636968456
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1636968456
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1636968456
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1636968456
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1636968456
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1636968456
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1636968456
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1636968456
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1636968456
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1185
timestamp 1636968456
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1205
timestamp 1636968456
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1217
timestamp 1636968456
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1229
timestamp 1636968456
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1241
timestamp 1636968456
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1261
timestamp 1636968456
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1273
timestamp 1
transform 1 0 118220 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1636968456
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1636968456
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1636968456
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1636968456
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1636968456
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_153
timestamp 1
transform 1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636968456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1636968456
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1636968456
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636968456
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_249
timestamp 1
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_253
timestamp 1636968456
transform 1 0 24380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1636968456
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_284
timestamp 1
transform 1 0 27232 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_290
timestamp 1
transform 1 0 27784 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_294
timestamp 1636968456
transform 1 0 28152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_306
timestamp 1
transform 1 0 29256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_312
timestamp 1
transform 1 0 29808 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_319
timestamp 1636968456
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636968456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636968456
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_365
timestamp 1636968456
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_377
timestamp 1636968456
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636968456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636968456
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_417
timestamp 1
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_421
timestamp 1636968456
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1636968456
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636968456
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636968456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_473
timestamp 1
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1636968456
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1636968456
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636968456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636968456
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_529
timestamp 1
transform 1 0 49772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1636968456
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1636968456
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1636968456
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1636968456
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_585
timestamp 1
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_589
timestamp 1636968456
transform 1 0 55292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_601
timestamp 1636968456
transform 1 0 56396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_613
timestamp 1
transform 1 0 57500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1636968456
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1636968456
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_641
timestamp 1
transform 1 0 60076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_645
timestamp 1636968456
transform 1 0 60444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_657
timestamp 1636968456
transform 1 0 61548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_669
timestamp 1
transform 1 0 62652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1636968456
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1636968456
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_697
timestamp 1
transform 1 0 65228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_701
timestamp 1636968456
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_713
timestamp 1636968456
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_725
timestamp 1
transform 1 0 67804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1636968456
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1636968456
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_753
timestamp 1
transform 1 0 70380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_757
timestamp 1636968456
transform 1 0 70748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_769
timestamp 1636968456
transform 1 0 71852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_781
timestamp 1
transform 1 0 72956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1636968456
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1636968456
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_809
timestamp 1
transform 1 0 75532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_813
timestamp 1636968456
transform 1 0 75900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_825
timestamp 1636968456
transform 1 0 77004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_837
timestamp 1
transform 1 0 78108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1636968456
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1636968456
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_865
timestamp 1
transform 1 0 80684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_869
timestamp 1636968456
transform 1 0 81052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_881
timestamp 1636968456
transform 1 0 82156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_893
timestamp 1
transform 1 0 83260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1636968456
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1636968456
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_925
timestamp 1636968456
transform 1 0 86204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_937
timestamp 1636968456
transform 1 0 87308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_949
timestamp 1
transform 1 0 88412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1636968456
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_965
timestamp 1636968456
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_977
timestamp 1
transform 1 0 90988 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_981
timestamp 1636968456
transform 1 0 91356 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_993
timestamp 1
transform 1 0 92460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1004
timestamp 1
transform 1 0 93472 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1636968456
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1636968456
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1033
timestamp 1
transform 1 0 96140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1636968456
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1049
timestamp 1636968456
transform 1 0 97612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1061
timestamp 1
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1636968456
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1636968456
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1089
timestamp 1
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1093
timestamp 1636968456
transform 1 0 101660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1105
timestamp 1636968456
transform 1 0 102764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1117
timestamp 1
transform 1 0 103868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1636968456
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1636968456
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1145
timestamp 1
transform 1 0 106444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1149
timestamp 1636968456
transform 1 0 106812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1161
timestamp 1636968456
transform 1 0 107916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1173
timestamp 1
transform 1 0 109020 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1636968456
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1189
timestamp 1636968456
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1201
timestamp 1
transform 1 0 111596 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1205
timestamp 1636968456
transform 1 0 111964 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1217
timestamp 1636968456
transform 1 0 113068 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1229
timestamp 1
transform 1 0 114172 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1233
timestamp 1636968456
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1245
timestamp 1636968456
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1257
timestamp 1
transform 1 0 116748 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1261
timestamp 1636968456
transform 1 0 117116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1273
timestamp 1
transform 1 0 118220 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636968456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1165
timestamp 1636968456
transform 1 0 108284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1177
timestamp 1636968456
transform 1 0 109388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1189
timestamp 1
transform 1 0 110492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1191
timestamp 1636968456
transform 1 0 110676 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1203
timestamp 1636968456
transform 1 0 111780 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1215
timestamp 1636968456
transform 1 0 112884 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1227
timestamp 1636968456
transform 1 0 113988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1239
timestamp 1
transform 1 0 115092 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1245
timestamp 1
transform 1 0 115644 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1247
timestamp 1636968456
transform 1 0 115828 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1259
timestamp 1636968456
transform 1 0 116932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1271
timestamp 1
transform 1 0 118036 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636968456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1165
timestamp 1636968456
transform 1 0 108284 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1177
timestamp 1636968456
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1189
timestamp 1636968456
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1201
timestamp 1636968456
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1213
timestamp 1
transform 1 0 112700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1217
timestamp 1
transform 1 0 113068 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1219
timestamp 1636968456
transform 1 0 113252 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1231
timestamp 1636968456
transform 1 0 114356 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1243
timestamp 1636968456
transform 1 0 115460 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1255
timestamp 1636968456
transform 1 0 116564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1267
timestamp 1
transform 1 0 117668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1273
timestamp 1
transform 1 0 118220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1275
timestamp 1
transform 1 0 118404 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636968456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_65
timestamp 1
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1165
timestamp 1636968456
transform 1 0 108284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1177
timestamp 1636968456
transform 1 0 109388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1189
timestamp 1
transform 1 0 110492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1191
timestamp 1636968456
transform 1 0 110676 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1203
timestamp 1636968456
transform 1 0 111780 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1215
timestamp 1636968456
transform 1 0 112884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1227
timestamp 1636968456
transform 1 0 113988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1239
timestamp 1
transform 1 0 115092 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1245
timestamp 1
transform 1 0 115644 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1247
timestamp 1636968456
transform 1 0 115828 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1259
timestamp 1636968456
transform 1 0 116932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1271
timestamp 1
transform 1 0 118036 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp 1
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1165
timestamp 1636968456
transform 1 0 108284 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1177
timestamp 1636968456
transform 1 0 109388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1189
timestamp 1636968456
transform 1 0 110492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1201
timestamp 1636968456
transform 1 0 111596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1213
timestamp 1
transform 1 0 112700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1217
timestamp 1
transform 1 0 113068 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1219
timestamp 1636968456
transform 1 0 113252 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1231
timestamp 1636968456
transform 1 0 114356 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1243
timestamp 1636968456
transform 1 0 115460 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1255
timestamp 1636968456
transform 1 0 116564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1267
timestamp 1
transform 1 0 117668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1273
timestamp 1
transform 1 0 118220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1275
timestamp 1
transform 1 0 118404 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636968456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636968456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1165
timestamp 1636968456
transform 1 0 108284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1177
timestamp 1636968456
transform 1 0 109388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1189
timestamp 1
transform 1 0 110492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1191
timestamp 1636968456
transform 1 0 110676 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1203
timestamp 1636968456
transform 1 0 111780 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1215
timestamp 1636968456
transform 1 0 112884 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1227
timestamp 1636968456
transform 1 0 113988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1239
timestamp 1
transform 1 0 115092 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1245
timestamp 1
transform 1 0 115644 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1247
timestamp 1636968456
transform 1 0 115828 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1259
timestamp 1636968456
transform 1 0 116932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1271
timestamp 1
transform 1 0 118036 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636968456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636968456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636968456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1165
timestamp 1636968456
transform 1 0 108284 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1177
timestamp 1636968456
transform 1 0 109388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1189
timestamp 1636968456
transform 1 0 110492 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1201
timestamp 1636968456
transform 1 0 111596 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1213
timestamp 1
transform 1 0 112700 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1217
timestamp 1
transform 1 0 113068 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1219
timestamp 1636968456
transform 1 0 113252 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1231
timestamp 1636968456
transform 1 0 114356 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1243
timestamp 1636968456
transform 1 0 115460 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1255
timestamp 1636968456
transform 1 0 116564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1267
timestamp 1
transform 1 0 117668 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1273
timestamp 1
transform 1 0 118220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1275
timestamp 1
transform 1 0 118404 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636968456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636968456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_65
timestamp 1
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1165
timestamp 1636968456
transform 1 0 108284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1177
timestamp 1636968456
transform 1 0 109388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1189
timestamp 1
transform 1 0 110492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1191
timestamp 1636968456
transform 1 0 110676 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1203
timestamp 1636968456
transform 1 0 111780 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1215
timestamp 1636968456
transform 1 0 112884 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1227
timestamp 1636968456
transform 1 0 113988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1239
timestamp 1
transform 1 0 115092 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1245
timestamp 1
transform 1 0 115644 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1247
timestamp 1636968456
transform 1 0 115828 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1259
timestamp 1636968456
transform 1 0 116932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1271
timestamp 1
transform 1 0 118036 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636968456
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636968456
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636968456
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1165
timestamp 1636968456
transform 1 0 108284 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1177
timestamp 1636968456
transform 1 0 109388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1189
timestamp 1636968456
transform 1 0 110492 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1201
timestamp 1636968456
transform 1 0 111596 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1213
timestamp 1
transform 1 0 112700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1217
timestamp 1
transform 1 0 113068 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1219
timestamp 1636968456
transform 1 0 113252 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1231
timestamp 1636968456
transform 1 0 114356 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1243
timestamp 1636968456
transform 1 0 115460 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1255
timestamp 1636968456
transform 1 0 116564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1267
timestamp 1
transform 1 0 117668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1273
timestamp 1
transform 1 0 118220 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1275
timestamp 1
transform 1 0 118404 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636968456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636968456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_65
timestamp 1
transform 1 0 7084 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1165
timestamp 1636968456
transform 1 0 108284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1177
timestamp 1636968456
transform 1 0 109388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1189
timestamp 1
transform 1 0 110492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1191
timestamp 1636968456
transform 1 0 110676 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1203
timestamp 1636968456
transform 1 0 111780 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1215
timestamp 1636968456
transform 1 0 112884 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1227
timestamp 1636968456
transform 1 0 113988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1239
timestamp 1
transform 1 0 115092 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1245
timestamp 1
transform 1 0 115644 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1247
timestamp 1636968456
transform 1 0 115828 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1259
timestamp 1636968456
transform 1 0 116932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1271
timestamp 1
transform 1 0 118036 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636968456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636968456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636968456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636968456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1165
timestamp 1636968456
transform 1 0 108284 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1177
timestamp 1636968456
transform 1 0 109388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1189
timestamp 1636968456
transform 1 0 110492 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1201
timestamp 1636968456
transform 1 0 111596 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1213
timestamp 1
transform 1 0 112700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1217
timestamp 1
transform 1 0 113068 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1219
timestamp 1636968456
transform 1 0 113252 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1231
timestamp 1636968456
transform 1 0 114356 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1243
timestamp 1636968456
transform 1 0 115460 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1255
timestamp 1636968456
transform 1 0 116564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1267
timestamp 1
transform 1 0 117668 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1273
timestamp 1
transform 1 0 118220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1275
timestamp 1
transform 1 0 118404 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636968456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636968456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636968456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_65
timestamp 1
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1165
timestamp 1636968456
transform 1 0 108284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1177
timestamp 1636968456
transform 1 0 109388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1189
timestamp 1
transform 1 0 110492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1191
timestamp 1636968456
transform 1 0 110676 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1203
timestamp 1636968456
transform 1 0 111780 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1215
timestamp 1636968456
transform 1 0 112884 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1227
timestamp 1636968456
transform 1 0 113988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1239
timestamp 1
transform 1 0 115092 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1245
timestamp 1
transform 1 0 115644 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1247
timestamp 1636968456
transform 1 0 115828 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1259
timestamp 1636968456
transform 1 0 116932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1271
timestamp 1
transform 1 0 118036 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636968456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636968456
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636968456
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636968456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1165
timestamp 1636968456
transform 1 0 108284 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1177
timestamp 1636968456
transform 1 0 109388 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1189
timestamp 1636968456
transform 1 0 110492 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1201
timestamp 1636968456
transform 1 0 111596 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_1213
timestamp 1
transform 1 0 112700 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1217
timestamp 1
transform 1 0 113068 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1219
timestamp 1636968456
transform 1 0 113252 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1231
timestamp 1636968456
transform 1 0 114356 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1243
timestamp 1636968456
transform 1 0 115460 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1255
timestamp 1636968456
transform 1 0 116564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1267
timestamp 1
transform 1 0 117668 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1273
timestamp 1
transform 1 0 118220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_1275
timestamp 1
transform 1 0 118404 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636968456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1165
timestamp 1636968456
transform 1 0 108284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1177
timestamp 1636968456
transform 1 0 109388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1189
timestamp 1
transform 1 0 110492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1191
timestamp 1636968456
transform 1 0 110676 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1203
timestamp 1636968456
transform 1 0 111780 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1215
timestamp 1636968456
transform 1 0 112884 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1227
timestamp 1636968456
transform 1 0 113988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1239
timestamp 1
transform 1 0 115092 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1245
timestamp 1
transform 1 0 115644 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1247
timestamp 1636968456
transform 1 0 115828 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1259
timestamp 1636968456
transform 1 0 116932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1271
timestamp 1
transform 1 0 118036 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636968456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636968456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1165
timestamp 1636968456
transform 1 0 108284 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1177
timestamp 1636968456
transform 1 0 109388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1189
timestamp 1636968456
transform 1 0 110492 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1201
timestamp 1636968456
transform 1 0 111596 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_1213
timestamp 1
transform 1 0 112700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1217
timestamp 1
transform 1 0 113068 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1219
timestamp 1636968456
transform 1 0 113252 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1231
timestamp 1636968456
transform 1 0 114356 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1243
timestamp 1636968456
transform 1 0 115460 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1255
timestamp 1636968456
transform 1 0 116564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1267
timestamp 1
transform 1 0 117668 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1273
timestamp 1
transform 1 0 118220 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_1275
timestamp 1
transform 1 0 118404 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636968456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_65
timestamp 1
transform 1 0 7084 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1165
timestamp 1636968456
transform 1 0 108284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1177
timestamp 1636968456
transform 1 0 109388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1189
timestamp 1
transform 1 0 110492 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1191
timestamp 1636968456
transform 1 0 110676 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1203
timestamp 1636968456
transform 1 0 111780 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1215
timestamp 1636968456
transform 1 0 112884 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1227
timestamp 1636968456
transform 1 0 113988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1239
timestamp 1
transform 1 0 115092 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1245
timestamp 1
transform 1 0 115644 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1247
timestamp 1636968456
transform 1 0 115828 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1259
timestamp 1636968456
transform 1 0 116932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1271
timestamp 1
transform 1 0 118036 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1636968456
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1636968456
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1636968456
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1636968456
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1165
timestamp 1636968456
transform 1 0 108284 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1177
timestamp 1636968456
transform 1 0 109388 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1189
timestamp 1636968456
transform 1 0 110492 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1201
timestamp 1636968456
transform 1 0 111596 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_1213
timestamp 1
transform 1 0 112700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1217
timestamp 1
transform 1 0 113068 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1219
timestamp 1636968456
transform 1 0 113252 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1231
timestamp 1636968456
transform 1 0 114356 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1243
timestamp 1636968456
transform 1 0 115460 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1255
timestamp 1636968456
transform 1 0 116564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1267
timestamp 1
transform 1 0 117668 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1273
timestamp 1
transform 1 0 118220 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_1275
timestamp 1
transform 1 0 118404 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1165
timestamp 1636968456
transform 1 0 108284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1177
timestamp 1636968456
transform 1 0 109388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1189
timestamp 1
transform 1 0 110492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1191
timestamp 1636968456
transform 1 0 110676 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1203
timestamp 1636968456
transform 1 0 111780 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1215
timestamp 1636968456
transform 1 0 112884 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1227
timestamp 1636968456
transform 1 0 113988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1239
timestamp 1
transform 1 0 115092 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1245
timestamp 1
transform 1 0 115644 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1247
timestamp 1636968456
transform 1 0 115828 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1259
timestamp 1636968456
transform 1 0 116932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1271
timestamp 1
transform 1 0 118036 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636968456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636968456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1165
timestamp 1636968456
transform 1 0 108284 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1177
timestamp 1636968456
transform 1 0 109388 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1189
timestamp 1636968456
transform 1 0 110492 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1201
timestamp 1636968456
transform 1 0 111596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_1213
timestamp 1
transform 1 0 112700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1217
timestamp 1
transform 1 0 113068 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1219
timestamp 1636968456
transform 1 0 113252 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1231
timestamp 1636968456
transform 1 0 114356 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1243
timestamp 1636968456
transform 1 0 115460 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1255
timestamp 1636968456
transform 1 0 116564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1267
timestamp 1
transform 1 0 117668 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1273
timestamp 1
transform 1 0 118220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_1275
timestamp 1
transform 1 0 118404 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636968456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_65
timestamp 1
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1165
timestamp 1636968456
transform 1 0 108284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1177
timestamp 1636968456
transform 1 0 109388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1189
timestamp 1
transform 1 0 110492 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1191
timestamp 1636968456
transform 1 0 110676 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1203
timestamp 1636968456
transform 1 0 111780 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1215
timestamp 1636968456
transform 1 0 112884 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1227
timestamp 1636968456
transform 1 0 113988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1239
timestamp 1
transform 1 0 115092 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1245
timestamp 1
transform 1 0 115644 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1247
timestamp 1636968456
transform 1 0 115828 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1259
timestamp 1636968456
transform 1 0 116932 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1271
timestamp 1
transform 1 0 118036 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636968456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636968456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636968456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1165
timestamp 1636968456
transform 1 0 108284 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1177
timestamp 1636968456
transform 1 0 109388 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1189
timestamp 1636968456
transform 1 0 110492 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1201
timestamp 1636968456
transform 1 0 111596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_1213
timestamp 1
transform 1 0 112700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1217
timestamp 1
transform 1 0 113068 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1219
timestamp 1636968456
transform 1 0 113252 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1231
timestamp 1636968456
transform 1 0 114356 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1243
timestamp 1636968456
transform 1 0 115460 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1255
timestamp 1636968456
transform 1 0 116564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1267
timestamp 1
transform 1 0 117668 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1273
timestamp 1
transform 1 0 118220 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_1275
timestamp 1
transform 1 0 118404 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636968456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636968456
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1165
timestamp 1636968456
transform 1 0 108284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1177
timestamp 1636968456
transform 1 0 109388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1189
timestamp 1
transform 1 0 110492 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1191
timestamp 1636968456
transform 1 0 110676 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1203
timestamp 1636968456
transform 1 0 111780 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1215
timestamp 1636968456
transform 1 0 112884 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1227
timestamp 1636968456
transform 1 0 113988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1239
timestamp 1
transform 1 0 115092 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1245
timestamp 1
transform 1 0 115644 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1247
timestamp 1636968456
transform 1 0 115828 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1259
timestamp 1636968456
transform 1 0 116932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1271
timestamp 1
transform 1 0 118036 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636968456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636968456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636968456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636968456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_69
timestamp 1
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1165
timestamp 1636968456
transform 1 0 108284 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1177
timestamp 1636968456
transform 1 0 109388 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1189
timestamp 1636968456
transform 1 0 110492 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1201
timestamp 1636968456
transform 1 0 111596 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_1213
timestamp 1
transform 1 0 112700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1217
timestamp 1
transform 1 0 113068 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1219
timestamp 1636968456
transform 1 0 113252 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1231
timestamp 1636968456
transform 1 0 114356 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1243
timestamp 1636968456
transform 1 0 115460 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1255
timestamp 1636968456
transform 1 0 116564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1267
timestamp 1
transform 1 0 117668 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1273
timestamp 1
transform 1 0 118220 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1275
timestamp 1
transform 1 0 118404 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636968456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636968456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636968456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636968456
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 1
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1165
timestamp 1636968456
transform 1 0 108284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1177
timestamp 1636968456
transform 1 0 109388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1189
timestamp 1
transform 1 0 110492 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1191
timestamp 1636968456
transform 1 0 110676 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1203
timestamp 1636968456
transform 1 0 111780 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1215
timestamp 1636968456
transform 1 0 112884 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1227
timestamp 1636968456
transform 1 0 113988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1239
timestamp 1
transform 1 0 115092 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1245
timestamp 1
transform 1 0 115644 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1247
timestamp 1636968456
transform 1 0 115828 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1259
timestamp 1636968456
transform 1 0 116932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1271
timestamp 1
transform 1 0 118036 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636968456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636968456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636968456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636968456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1165
timestamp 1636968456
transform 1 0 108284 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1177
timestamp 1636968456
transform 1 0 109388 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1189
timestamp 1636968456
transform 1 0 110492 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1201
timestamp 1636968456
transform 1 0 111596 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_1213
timestamp 1
transform 1 0 112700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1217
timestamp 1
transform 1 0 113068 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1219
timestamp 1636968456
transform 1 0 113252 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1231
timestamp 1636968456
transform 1 0 114356 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1243
timestamp 1636968456
transform 1 0 115460 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1255
timestamp 1636968456
transform 1 0 116564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1267
timestamp 1
transform 1 0 117668 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1273
timestamp 1
transform 1 0 118220 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_1275
timestamp 1
transform 1 0 118404 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636968456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636968456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636968456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636968456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636968456
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_65
timestamp 1
transform 1 0 7084 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1165
timestamp 1636968456
transform 1 0 108284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1177
timestamp 1636968456
transform 1 0 109388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1189
timestamp 1
transform 1 0 110492 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1191
timestamp 1636968456
transform 1 0 110676 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1203
timestamp 1636968456
transform 1 0 111780 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1215
timestamp 1636968456
transform 1 0 112884 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1227
timestamp 1636968456
transform 1 0 113988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1239
timestamp 1
transform 1 0 115092 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1245
timestamp 1
transform 1 0 115644 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1247
timestamp 1636968456
transform 1 0 115828 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1259
timestamp 1636968456
transform 1 0 116932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1271
timestamp 1
transform 1 0 118036 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636968456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636968456
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636968456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636968456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1165
timestamp 1636968456
transform 1 0 108284 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1177
timestamp 1636968456
transform 1 0 109388 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1189
timestamp 1636968456
transform 1 0 110492 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1201
timestamp 1636968456
transform 1 0 111596 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_1213
timestamp 1
transform 1 0 112700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1217
timestamp 1
transform 1 0 113068 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1219
timestamp 1636968456
transform 1 0 113252 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1231
timestamp 1636968456
transform 1 0 114356 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1243
timestamp 1636968456
transform 1 0 115460 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1255
timestamp 1636968456
transform 1 0 116564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1267
timestamp 1
transform 1 0 117668 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1273
timestamp 1
transform 1 0 118220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_1275
timestamp 1
transform 1 0 118404 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636968456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636968456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636968456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636968456
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_65
timestamp 1
transform 1 0 7084 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1165
timestamp 1636968456
transform 1 0 108284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1177
timestamp 1636968456
transform 1 0 109388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1189
timestamp 1
transform 1 0 110492 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1191
timestamp 1636968456
transform 1 0 110676 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1203
timestamp 1636968456
transform 1 0 111780 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1215
timestamp 1636968456
transform 1 0 112884 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1227
timestamp 1636968456
transform 1 0 113988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1239
timestamp 1
transform 1 0 115092 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1245
timestamp 1
transform 1 0 115644 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1247
timestamp 1636968456
transform 1 0 115828 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1259
timestamp 1636968456
transform 1 0 116932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1271
timestamp 1
transform 1 0 118036 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636968456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636968456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636968456
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636968456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1165
timestamp 1636968456
transform 1 0 108284 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1177
timestamp 1636968456
transform 1 0 109388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1189
timestamp 1636968456
transform 1 0 110492 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1201
timestamp 1636968456
transform 1 0 111596 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_1213
timestamp 1
transform 1 0 112700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1217
timestamp 1
transform 1 0 113068 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1219
timestamp 1636968456
transform 1 0 113252 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1231
timestamp 1636968456
transform 1 0 114356 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1243
timestamp 1636968456
transform 1 0 115460 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1255
timestamp 1636968456
transform 1 0 116564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1267
timestamp 1
transform 1 0 117668 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1273
timestamp 1
transform 1 0 118220 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_1275
timestamp 1
transform 1 0 118404 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636968456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636968456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636968456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636968456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1165
timestamp 1636968456
transform 1 0 108284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1177
timestamp 1636968456
transform 1 0 109388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1189
timestamp 1
transform 1 0 110492 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1191
timestamp 1636968456
transform 1 0 110676 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1203
timestamp 1636968456
transform 1 0 111780 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1215
timestamp 1636968456
transform 1 0 112884 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1227
timestamp 1636968456
transform 1 0 113988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1239
timestamp 1
transform 1 0 115092 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1245
timestamp 1
transform 1 0 115644 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1247
timestamp 1636968456
transform 1 0 115828 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1259
timestamp 1636968456
transform 1 0 116932 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1271
timestamp 1
transform 1 0 118036 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636968456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636968456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636968456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636968456
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636968456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_69
timestamp 1
transform 1 0 7452 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1165
timestamp 1636968456
transform 1 0 108284 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1177
timestamp 1636968456
transform 1 0 109388 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1189
timestamp 1636968456
transform 1 0 110492 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1201
timestamp 1636968456
transform 1 0 111596 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_1213
timestamp 1
transform 1 0 112700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1217
timestamp 1
transform 1 0 113068 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1219
timestamp 1636968456
transform 1 0 113252 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1231
timestamp 1636968456
transform 1 0 114356 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1243
timestamp 1636968456
transform 1 0 115460 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1255
timestamp 1636968456
transform 1 0 116564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1267
timestamp 1
transform 1 0 117668 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1273
timestamp 1
transform 1 0 118220 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_1275
timestamp 1
transform 1 0 118404 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636968456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636968456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636968456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_65
timestamp 1
transform 1 0 7084 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1165
timestamp 1636968456
transform 1 0 108284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1177
timestamp 1636968456
transform 1 0 109388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1189
timestamp 1
transform 1 0 110492 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1191
timestamp 1636968456
transform 1 0 110676 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1203
timestamp 1636968456
transform 1 0 111780 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1215
timestamp 1636968456
transform 1 0 112884 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1227
timestamp 1636968456
transform 1 0 113988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1239
timestamp 1
transform 1 0 115092 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1245
timestamp 1
transform 1 0 115644 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1247
timestamp 1636968456
transform 1 0 115828 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1259
timestamp 1636968456
transform 1 0 116932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1271
timestamp 1
transform 1 0 118036 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636968456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636968456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636968456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636968456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1165
timestamp 1636968456
transform 1 0 108284 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1177
timestamp 1636968456
transform 1 0 109388 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1189
timestamp 1636968456
transform 1 0 110492 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1201
timestamp 1636968456
transform 1 0 111596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_1213
timestamp 1
transform 1 0 112700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1217
timestamp 1
transform 1 0 113068 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1219
timestamp 1636968456
transform 1 0 113252 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1231
timestamp 1636968456
transform 1 0 114356 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1243
timestamp 1636968456
transform 1 0 115460 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1255
timestamp 1636968456
transform 1 0 116564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1267
timestamp 1
transform 1 0 117668 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1273
timestamp 1
transform 1 0 118220 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_1275
timestamp 1
transform 1 0 118404 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636968456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636968456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636968456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636968456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1165
timestamp 1636968456
transform 1 0 108284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1177
timestamp 1636968456
transform 1 0 109388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1189
timestamp 1
transform 1 0 110492 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1191
timestamp 1636968456
transform 1 0 110676 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1203
timestamp 1636968456
transform 1 0 111780 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1215
timestamp 1636968456
transform 1 0 112884 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1227
timestamp 1636968456
transform 1 0 113988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1239
timestamp 1
transform 1 0 115092 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1245
timestamp 1
transform 1 0 115644 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1247
timestamp 1636968456
transform 1 0 115828 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1259
timestamp 1636968456
transform 1 0 116932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1271
timestamp 1
transform 1 0 118036 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636968456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636968456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1165
timestamp 1636968456
transform 1 0 108284 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1177
timestamp 1636968456
transform 1 0 109388 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1189
timestamp 1636968456
transform 1 0 110492 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1201
timestamp 1636968456
transform 1 0 111596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_1213
timestamp 1
transform 1 0 112700 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1217
timestamp 1
transform 1 0 113068 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1219
timestamp 1636968456
transform 1 0 113252 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_1231
timestamp 1
transform 1 0 114356 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1235
timestamp 1
transform 1 0 114724 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1240
timestamp 1636968456
transform 1 0 115184 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1252
timestamp 1636968456
transform 1 0 116288 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1264
timestamp 1
transform 1 0 117392 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_1272
timestamp 1
transform 1 0 118128 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_1275
timestamp 1
transform 1 0 118404 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636968456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636968456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_65
timestamp 1
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1165
timestamp 1636968456
transform 1 0 108284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1177
timestamp 1636968456
transform 1 0 109388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1189
timestamp 1
transform 1 0 110492 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_1191
timestamp 1
transform 1 0 110676 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1204
timestamp 1636968456
transform 1 0 111872 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1216
timestamp 1636968456
transform 1 0 112976 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1228
timestamp 1
transform 1 0 114080 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_1244
timestamp 1
transform 1 0 115552 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1247
timestamp 1636968456
transform 1 0 115828 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1259
timestamp 1636968456
transform 1 0 116932 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1271
timestamp 1
transform 1 0 118036 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636968456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636968456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636968456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1165
timestamp 1636968456
transform 1 0 108284 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1177
timestamp 1636968456
transform 1 0 109388 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_1189
timestamp 1
transform 1 0 110492 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_1199
timestamp 1
transform 1 0 111412 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1209
timestamp 1
transform 1 0 112332 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1217
timestamp 1
transform 1 0 113068 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1219
timestamp 1
transform 1 0 113252 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1227
timestamp 1
transform 1 0 113988 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1233
timestamp 1
transform 1 0 114540 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1251
timestamp 1636968456
transform 1 0 116196 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1263
timestamp 1
transform 1 0 117300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_1271
timestamp 1
transform 1 0 118036 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_65
timestamp 1
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1165
timestamp 1636968456
transform 1 0 108284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_1177
timestamp 1
transform 1 0 109388 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1189
timestamp 1
transform 1 0 110492 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_1214
timestamp 1
transform 1 0 112792 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1239
timestamp 1
transform 1 0 115092 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1253
timestamp 1
transform 1 0 116380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1260
timestamp 1
transform 1 0 117024 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1264
timestamp 1
transform 1 0 117392 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_69
timestamp 1
transform 1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1165
timestamp 1636968456
transform 1 0 108284 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_1177
timestamp 1
transform 1 0 109388 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1186
timestamp 1
transform 1 0 110216 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_1194
timestamp 1
transform 1 0 110952 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1205
timestamp 1
transform 1 0 111964 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_1214
timestamp 1
transform 1 0 112792 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_1219
timestamp 1
transform 1 0 113252 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_1239
timestamp 1
transform 1 0 115092 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1243
timestamp 1
transform 1 0 115460 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_1247
timestamp 1
transform 1 0 115828 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_65
timestamp 1
transform 1 0 7084 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1165
timestamp 1636968456
transform 1 0 108284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_1177
timestamp 1
transform 1 0 109388 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_1187
timestamp 1
transform 1 0 110308 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_1196
timestamp 1
transform 1 0 111136 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1204
timestamp 1
transform 1 0 111872 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1213
timestamp 1
transform 1 0 112700 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_1223
timestamp 1
transform 1 0 113620 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_1242
timestamp 1
transform 1 0 115368 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_1252
timestamp 1
transform 1 0 116288 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1270
timestamp 1
transform 1 0 117944 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636968456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636968456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636968456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1636968456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636968456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1
transform 1 0 7452 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1165
timestamp 1636968456
transform 1 0 108284 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_1191
timestamp 1
transform 1 0 110676 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1201
timestamp 1636968456
transform 1 0 111596 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_1213
timestamp 1
transform 1 0 112700 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1217
timestamp 1
transform 1 0 113068 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1219
timestamp 1
transform 1 0 113252 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1229
timestamp 1
transform 1 0 114172 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1266
timestamp 1
transform 1 0 117576 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1273
timestamp 1
transform 1 0 118220 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636968456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_65
timestamp 1
transform 1 0 7084 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1165
timestamp 1
transform 1 0 108284 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_1173
timestamp 1
transform 1 0 109020 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1182
timestamp 1
transform 1 0 109848 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_1187
timestamp 1
transform 1 0 110308 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_1198
timestamp 1
transform 1 0 111320 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_1205
timestamp 1
transform 1 0 111964 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_1223
timestamp 1
transform 1 0 113620 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1230
timestamp 1
transform 1 0 114264 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1236
timestamp 1
transform 1 0 114816 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1240
timestamp 1
transform 1 0 115184 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1265
timestamp 1
transform 1 0 117484 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636968456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636968456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_69
timestamp 1
transform 1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1165
timestamp 1
transform 1 0 108284 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1173
timestamp 1
transform 1 0 109020 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1200
timestamp 1
transform 1 0 111504 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1209
timestamp 1
transform 1 0 112332 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1217
timestamp 1
transform 1 0 113068 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1230
timestamp 1
transform 1 0 114264 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1238
timestamp 1
transform 1 0 115000 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1263
timestamp 1
transform 1 0 117300 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636968456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636968456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_65
timestamp 1
transform 1 0 7084 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_1165
timestamp 1
transform 1 0 108284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1183
timestamp 1
transform 1 0 109940 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1189
timestamp 1
transform 1 0 110492 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_1191
timestamp 1
transform 1 0 110676 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1213
timestamp 1
transform 1 0 112700 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_1237
timestamp 1
transform 1 0 114908 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1245
timestamp 1
transform 1 0 115644 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_1275
timestamp 1
transform 1 0 118404 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636968456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636968456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636968456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1636968456
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_69
timestamp 1
transform 1 0 7452 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_1165
timestamp 1
transform 1 0 108284 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_1177
timestamp 1
transform 1 0 109388 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1185
timestamp 1
transform 1 0 110124 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1195
timestamp 1
transform 1 0 111044 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_1201
timestamp 1
transform 1 0 111596 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1207
timestamp 1
transform 1 0 112148 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_1219
timestamp 1
transform 1 0 113252 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1245
timestamp 1
transform 1 0 115644 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1257
timestamp 1
transform 1 0 116748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_1269
timestamp 1
transform 1 0 117852 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636968456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636968456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636968456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1636968456
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1636968456
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_65
timestamp 1
transform 1 0 7084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1176
timestamp 1
transform 1 0 109296 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1184
timestamp 1
transform 1 0 110032 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_1191
timestamp 1
transform 1 0 110676 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1208
timestamp 1
transform 1 0 112240 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636968456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636968456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1636968456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1636968456
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1636968456
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_69
timestamp 1
transform 1 0 7452 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_1186
timestamp 1
transform 1 0 110216 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1199
timestamp 1
transform 1 0 111412 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1216
timestamp 1
transform 1 0 112976 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1224
timestamp 1
transform 1 0 113712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_1233
timestamp 1
transform 1 0 114540 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1239
timestamp 1
transform 1 0 115092 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1247
timestamp 1
transform 1 0 115828 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1273
timestamp 1
transform 1 0 118220 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1275
timestamp 1
transform 1 0 118404 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636968456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636968456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636968456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636968456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1636968456
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_65
timestamp 1
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_1171
timestamp 1
transform 1 0 108836 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_1176
timestamp 1
transform 1 0 109296 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1191
timestamp 1636968456
transform 1 0 110676 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_1203
timestamp 1
transform 1 0 111780 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_1211
timestamp 1
transform 1 0 112516 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_1216
timestamp 1
transform 1 0 112976 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1221
timestamp 1636968456
transform 1 0 113436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1233
timestamp 1
transform 1 0 114540 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1239
timestamp 1
transform 1 0 115092 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_1274
timestamp 1
transform 1 0 118312 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636968456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636968456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636968456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636968456
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636968456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_69
timestamp 1
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_1183
timestamp 1
transform 1 0 109940 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1217
timestamp 1
transform 1 0 113068 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_1219
timestamp 1
transform 1 0 113252 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_1230
timestamp 1
transform 1 0 114264 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_1250
timestamp 1
transform 1 0 116104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_1256
timestamp 1
transform 1 0 116656 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1268
timestamp 1
transform 1 0 117760 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_1275
timestamp 1
transform 1 0 118404 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636968456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636968456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636968456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636968456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636968456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_65
timestamp 1
transform 1 0 7084 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_1165
timestamp 1
transform 1 0 108284 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1172
timestamp 1
transform 1 0 108928 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_1179
timestamp 1
transform 1 0 109572 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1189
timestamp 1
transform 1 0 110492 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_1191
timestamp 1
transform 1 0 110676 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_1197
timestamp 1
transform 1 0 111228 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1206
timestamp 1636968456
transform 1 0 112056 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_1218
timestamp 1
transform 1 0 113160 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1231
timestamp 1
transform 1 0 114356 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1245
timestamp 1
transform 1 0 115644 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_1252
timestamp 1
transform 1 0 116288 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_1273
timestamp 1
transform 1 0 118220 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636968456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636968456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636968456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636968456
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636968456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_69
timestamp 1
transform 1 0 7452 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1165
timestamp 1
transform 1 0 108284 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1170
timestamp 1
transform 1 0 108744 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1197
timestamp 1
transform 1 0 111228 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1210
timestamp 1
transform 1 0 112424 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_1219
timestamp 1
transform 1 0 113252 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1232
timestamp 1
transform 1 0 114448 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1250
timestamp 1
transform 1 0 116104 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1258
timestamp 1
transform 1 0 116840 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1268
timestamp 1
transform 1 0 117760 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1275
timestamp 1
transform 1 0 118404 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636968456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636968456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636968456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636968456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636968456
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_65
timestamp 1
transform 1 0 7084 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_1165
timestamp 1
transform 1 0 108284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1173
timestamp 1
transform 1 0 109020 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1177
timestamp 1
transform 1 0 109388 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_1188
timestamp 1
transform 1 0 110400 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1191
timestamp 1
transform 1 0 110676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1195
timestamp 1
transform 1 0 111044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1203
timestamp 1
transform 1 0 111780 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1207
timestamp 1
transform 1 0 112148 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1231
timestamp 1
transform 1 0 114356 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_1247
timestamp 1
transform 1 0 115828 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1256
timestamp 1
transform 1 0 116656 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_8
timestamp 1636968456
transform 1 0 1840 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_20
timestamp 1636968456
transform 1 0 2944 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_32
timestamp 1636968456
transform 1 0 4048 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_44
timestamp 1636968456
transform 1 0 5152 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636968456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_69
timestamp 1
transform 1 0 7452 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_1165
timestamp 1
transform 1 0 108284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1184
timestamp 1
transform 1 0 110032 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1196
timestamp 1
transform 1 0 111136 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1205
timestamp 1
transform 1 0 111964 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1213
timestamp 1
transform 1 0 112700 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1219
timestamp 1
transform 1 0 113252 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1228
timestamp 1
transform 1 0 114080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1236
timestamp 1
transform 1 0 114816 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1245
timestamp 1
transform 1 0 115644 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1275
timestamp 1
transform 1 0 118404 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636968456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636968456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636968456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636968456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1636968456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_65
timestamp 1
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1165
timestamp 1
transform 1 0 108284 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1173
timestamp 1
transform 1 0 109020 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1179
timestamp 1
transform 1 0 109572 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1189
timestamp 1
transform 1 0 110492 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1198
timestamp 1
transform 1 0 111320 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1202
timestamp 1
transform 1 0 111688 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1228
timestamp 1
transform 1 0 114080 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1245
timestamp 1
transform 1 0 115644 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1262
timestamp 1636968456
transform 1 0 117208 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_1274
timestamp 1
transform 1 0 118312 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636968456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636968456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1636968456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1636968456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1636968456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_69
timestamp 1
transform 1 0 7452 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1187
timestamp 1
transform 1 0 110308 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1197
timestamp 1
transform 1 0 111228 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1205
timestamp 1
transform 1 0 111964 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_1215
timestamp 1
transform 1 0 112884 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1260
timestamp 1636968456
transform 1 0 117024 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1272
timestamp 1
transform 1 0 118128 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1275
timestamp 1
transform 1 0 118404 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636968456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636968456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636968456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1636968456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1636968456
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_65
timestamp 1
transform 1 0 7084 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_1165
timestamp 1
transform 1 0 108284 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1173
timestamp 1
transform 1 0 109020 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1179
timestamp 1
transform 1 0 109572 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1184
timestamp 1
transform 1 0 110032 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1191
timestamp 1
transform 1 0 110676 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1201
timestamp 1
transform 1 0 111596 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1215
timestamp 1
transform 1 0 112884 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1242
timestamp 1
transform 1 0 115368 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1256
timestamp 1636968456
transform 1 0 116656 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_1268
timestamp 1
transform 1 0 117760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1276
timestamp 1
transform 1 0 118496 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_8
timestamp 1636968456
transform 1 0 1840 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_20
timestamp 1636968456
transform 1 0 2944 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_32
timestamp 1636968456
transform 1 0 4048 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_44
timestamp 1636968456
transform 1 0 5152 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1636968456
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_69
timestamp 1
transform 1 0 7452 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_1165
timestamp 1
transform 1 0 108284 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1173
timestamp 1
transform 1 0 109020 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1179
timestamp 1
transform 1 0 109572 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_1196
timestamp 1
transform 1 0 111136 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_1204
timestamp 1
transform 1 0 111872 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_1213
timestamp 1
transform 1 0 112700 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1217
timestamp 1
transform 1 0 113068 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_1219
timestamp 1
transform 1 0 113252 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_1229
timestamp 1
transform 1 0 114172 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1234
timestamp 1636968456
transform 1 0 114632 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1246
timestamp 1636968456
transform 1 0 115736 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1258
timestamp 1636968456
transform 1 0 116840 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_1270
timestamp 1
transform 1 0 117944 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_1275
timestamp 1
transform 1 0 118404 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_8
timestamp 1636968456
transform 1 0 1840 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_20
timestamp 1
transform 1 0 2944 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636968456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1636968456
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1636968456
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_65
timestamp 1
transform 1 0 7084 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_66_1165
timestamp 1
transform 1 0 108284 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_1188
timestamp 1
transform 1 0 110400 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_1191
timestamp 1
transform 1 0 110676 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_1199
timestamp 1
transform 1 0 111412 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1207
timestamp 1636968456
transform 1 0 112148 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1219
timestamp 1636968456
transform 1 0 113252 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1231
timestamp 1636968456
transform 1 0 114356 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_1243
timestamp 1
transform 1 0 115460 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1247
timestamp 1636968456
transform 1 0 115828 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1259
timestamp 1636968456
transform 1 0 116932 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_1271
timestamp 1
transform 1 0 118036 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636968456
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636968456
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1636968456
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1636968456
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636968456
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_69
timestamp 1
transform 1 0 7452 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1165
timestamp 1
transform 1 0 108284 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_1173
timestamp 1
transform 1 0 109020 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_67_1189
timestamp 1
transform 1 0 110492 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1197
timestamp 1636968456
transform 1 0 111228 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1209
timestamp 1
transform 1 0 112332 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_1217
timestamp 1
transform 1 0 113068 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1219
timestamp 1636968456
transform 1 0 113252 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1231
timestamp 1636968456
transform 1 0 114356 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1243
timestamp 1636968456
transform 1 0 115460 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1255
timestamp 1636968456
transform 1 0 116564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_1267
timestamp 1
transform 1 0 117668 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_1273
timestamp 1
transform 1 0 118220 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_1275
timestamp 1
transform 1 0 118404 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636968456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636968456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636968456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636968456
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636968456
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_65
timestamp 1
transform 1 0 7084 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_1165
timestamp 1
transform 1 0 108284 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1193
timestamp 1636968456
transform 1 0 110860 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1205
timestamp 1636968456
transform 1 0 111964 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1217
timestamp 1636968456
transform 1 0 113068 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1229
timestamp 1636968456
transform 1 0 114172 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_1241
timestamp 1
transform 1 0 115276 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1245
timestamp 1
transform 1 0 115644 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1247
timestamp 1636968456
transform 1 0 115828 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1259
timestamp 1636968456
transform 1 0 116932 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_1271
timestamp 1
transform 1 0 118036 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636968456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636968456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636968456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636968456
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636968456
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_69
timestamp 1
transform 1 0 7452 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1165
timestamp 1636968456
transform 1 0 108284 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_1187
timestamp 1
transform 1 0 110308 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1198
timestamp 1636968456
transform 1 0 111320 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_1210
timestamp 1
transform 1 0 112424 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1219
timestamp 1636968456
transform 1 0 113252 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1231
timestamp 1636968456
transform 1 0 114356 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1243
timestamp 1636968456
transform 1 0 115460 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1255
timestamp 1636968456
transform 1 0 116564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_1267
timestamp 1
transform 1 0 117668 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_1273
timestamp 1
transform 1 0 118220 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_1275
timestamp 1
transform 1 0 118404 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_8
timestamp 1636968456
transform 1 0 1840 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_20
timestamp 1
transform 1 0 2944 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636968456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636968456
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636968456
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_65
timestamp 1
transform 1 0 7084 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1198
timestamp 1636968456
transform 1 0 111320 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1210
timestamp 1636968456
transform 1 0 112424 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1222
timestamp 1636968456
transform 1 0 113528 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1234
timestamp 1636968456
transform 1 0 114632 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1247
timestamp 1636968456
transform 1 0 115828 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1259
timestamp 1636968456
transform 1 0 116932 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_1271
timestamp 1
transform 1 0 118036 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_8
timestamp 1636968456
transform 1 0 1840 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_20
timestamp 1636968456
transform 1 0 2944 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_32
timestamp 1636968456
transform 1 0 4048 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_44
timestamp 1636968456
transform 1 0 5152 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636968456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_69
timestamp 1
transform 1 0 7452 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1165
timestamp 1636968456
transform 1 0 108284 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_1177
timestamp 1
transform 1 0 109388 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1186
timestamp 1
transform 1 0 110216 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1196
timestamp 1636968456
transform 1 0 111136 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_1208
timestamp 1
transform 1 0 112240 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1216
timestamp 1
transform 1 0 112976 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1219
timestamp 1636968456
transform 1 0 113252 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1231
timestamp 1636968456
transform 1 0 114356 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1243
timestamp 1636968456
transform 1 0 115460 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1255
timestamp 1636968456
transform 1 0 116564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_1267
timestamp 1
transform 1 0 117668 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_1273
timestamp 1
transform 1 0 118220 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1275
timestamp 1
transform 1 0 118404 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636968456
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636968456
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636968456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636968456
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636968456
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_65
timestamp 1
transform 1 0 7084 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_1170
timestamp 1
transform 1 0 108744 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_1185
timestamp 1
transform 1 0 110124 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_1189
timestamp 1
transform 1 0 110492 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1194
timestamp 1636968456
transform 1 0 110952 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1206
timestamp 1636968456
transform 1 0 112056 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1218
timestamp 1636968456
transform 1 0 113160 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1230
timestamp 1636968456
transform 1 0 114264 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_1242
timestamp 1
transform 1 0 115368 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1247
timestamp 1636968456
transform 1 0 115828 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1259
timestamp 1636968456
transform 1 0 116932 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_1271
timestamp 1
transform 1 0 118036 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636968456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636968456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636968456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636968456
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636968456
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_69
timestamp 1
transform 1 0 7452 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_1165
timestamp 1
transform 1 0 108284 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1188
timestamp 1636968456
transform 1 0 110400 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1200
timestamp 1636968456
transform 1 0 111504 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_1212
timestamp 1
transform 1 0 112608 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1219
timestamp 1636968456
transform 1 0 113252 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1231
timestamp 1636968456
transform 1 0 114356 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1243
timestamp 1636968456
transform 1 0 115460 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1255
timestamp 1636968456
transform 1 0 116564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_1267
timestamp 1
transform 1 0 117668 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_1273
timestamp 1
transform 1 0 118220 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_1275
timestamp 1
transform 1 0 118404 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636968456
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636968456
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636968456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636968456
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636968456
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_65
timestamp 1
transform 1 0 7084 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1165
timestamp 1
transform 1 0 108284 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_1171
timestamp 1
transform 1 0 108836 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_1183
timestamp 1
transform 1 0 109940 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1189
timestamp 1
transform 1 0 110492 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1191
timestamp 1636968456
transform 1 0 110676 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1203
timestamp 1636968456
transform 1 0 111780 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1215
timestamp 1636968456
transform 1 0 112884 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1227
timestamp 1636968456
transform 1 0 113988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_1239
timestamp 1
transform 1 0 115092 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1245
timestamp 1
transform 1 0 115644 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1247
timestamp 1636968456
transform 1 0 115828 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1259
timestamp 1636968456
transform 1 0 116932 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_1271
timestamp 1
transform 1 0 118036 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_8
timestamp 1636968456
transform 1 0 1840 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_20
timestamp 1636968456
transform 1 0 2944 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_32
timestamp 1636968456
transform 1 0 4048 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_44
timestamp 1636968456
transform 1 0 5152 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636968456
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_69
timestamp 1
transform 1 0 7452 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_1165
timestamp 1
transform 1 0 108284 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_1173
timestamp 1
transform 1 0 109020 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1189
timestamp 1636968456
transform 1 0 110492 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1201
timestamp 1636968456
transform 1 0 111596 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_1213
timestamp 1
transform 1 0 112700 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_1217
timestamp 1
transform 1 0 113068 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1219
timestamp 1636968456
transform 1 0 113252 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1231
timestamp 1636968456
transform 1 0 114356 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1243
timestamp 1636968456
transform 1 0 115460 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1255
timestamp 1636968456
transform 1 0 116564 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_1267
timestamp 1
transform 1 0 117668 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_1273
timestamp 1
transform 1 0 118220 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_1275
timestamp 1
transform 1 0 118404 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636968456
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636968456
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636968456
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1636968456
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1636968456
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_65
timestamp 1
transform 1 0 7084 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_76_1170
timestamp 1
transform 1 0 108744 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1178
timestamp 1
transform 1 0 109480 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1189
timestamp 1
transform 1 0 110492 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1191
timestamp 1636968456
transform 1 0 110676 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1203
timestamp 1636968456
transform 1 0 111780 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1215
timestamp 1636968456
transform 1 0 112884 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1227
timestamp 1636968456
transform 1 0 113988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1239
timestamp 1
transform 1 0 115092 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1245
timestamp 1
transform 1 0 115644 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1247
timestamp 1636968456
transform 1 0 115828 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1259
timestamp 1636968456
transform 1 0 116932 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1271
timestamp 1
transform 1 0 118036 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_8
timestamp 1636968456
transform 1 0 1840 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_20
timestamp 1636968456
transform 1 0 2944 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_32
timestamp 1636968456
transform 1 0 4048 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_44
timestamp 1636968456
transform 1 0 5152 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1636968456
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_69
timestamp 1
transform 1 0 7452 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1170
timestamp 1636968456
transform 1 0 108744 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1182
timestamp 1636968456
transform 1 0 109848 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1194
timestamp 1636968456
transform 1 0 110952 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1206
timestamp 1636968456
transform 1 0 112056 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1219
timestamp 1636968456
transform 1 0 113252 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1231
timestamp 1636968456
transform 1 0 114356 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1243
timestamp 1636968456
transform 1 0 115460 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1255
timestamp 1636968456
transform 1 0 116564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_1267
timestamp 1
transform 1 0 117668 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_1273
timestamp 1
transform 1 0 118220 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_1275
timestamp 1
transform 1 0 118404 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636968456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636968456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636968456
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1636968456
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1636968456
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_65
timestamp 1
transform 1 0 7084 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1165
timestamp 1636968456
transform 1 0 108284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_1180
timestamp 1
transform 1 0 109664 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_1188
timestamp 1
transform 1 0 110400 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1191
timestamp 1636968456
transform 1 0 110676 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1203
timestamp 1636968456
transform 1 0 111780 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1215
timestamp 1636968456
transform 1 0 112884 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1227
timestamp 1636968456
transform 1 0 113988 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_1239
timestamp 1
transform 1 0 115092 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_1245
timestamp 1
transform 1 0 115644 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1247
timestamp 1636968456
transform 1 0 115828 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1259
timestamp 1636968456
transform 1 0 116932 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_1271
timestamp 1
transform 1 0 118036 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636968456
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636968456
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636968456
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1636968456
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1636968456
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_69
timestamp 1
transform 1 0 7452 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_1167
timestamp 1
transform 1 0 108468 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1193
timestamp 1636968456
transform 1 0 110860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1205
timestamp 1636968456
transform 1 0 111964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_1217
timestamp 1
transform 1 0 113068 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1219
timestamp 1636968456
transform 1 0 113252 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1231
timestamp 1636968456
transform 1 0 114356 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1243
timestamp 1636968456
transform 1 0 115460 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1255
timestamp 1636968456
transform 1 0 116564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_1267
timestamp 1
transform 1 0 117668 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_1273
timestamp 1
transform 1 0 118220 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_1275
timestamp 1
transform 1 0 118404 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636968456
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636968456
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636968456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1636968456
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1636968456
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_65
timestamp 1
transform 1 0 7084 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1168
timestamp 1
transform 1 0 108560 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1189
timestamp 1
transform 1 0 110492 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1191
timestamp 1636968456
transform 1 0 110676 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1203
timestamp 1636968456
transform 1 0 111780 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1215
timestamp 1636968456
transform 1 0 112884 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1227
timestamp 1636968456
transform 1 0 113988 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_1239
timestamp 1
transform 1 0 115092 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1245
timestamp 1
transform 1 0 115644 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1247
timestamp 1636968456
transform 1 0 115828 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1259
timestamp 1636968456
transform 1 0 116932 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_1271
timestamp 1
transform 1 0 118036 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636968456
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636968456
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1636968456
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1636968456
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1636968456
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_69
timestamp 1
transform 1 0 7452 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_1165
timestamp 1
transform 1 0 108284 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_1173
timestamp 1
transform 1 0 109020 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1182
timestamp 1636968456
transform 1 0 109848 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1194
timestamp 1636968456
transform 1 0 110952 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1206
timestamp 1636968456
transform 1 0 112056 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1219
timestamp 1636968456
transform 1 0 113252 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1231
timestamp 1636968456
transform 1 0 114356 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1243
timestamp 1636968456
transform 1 0 115460 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1255
timestamp 1636968456
transform 1 0 116564 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_1267
timestamp 1
transform 1 0 117668 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_1273
timestamp 1
transform 1 0 118220 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_1275
timestamp 1
transform 1 0 118404 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636968456
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636968456
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636968456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1636968456
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1636968456
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_65
timestamp 1
transform 1 0 7084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_82_1165
timestamp 1
transform 1 0 108284 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1189
timestamp 1
transform 1 0 110492 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1193
timestamp 1636968456
transform 1 0 110860 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1205
timestamp 1636968456
transform 1 0 111964 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1217
timestamp 1636968456
transform 1 0 113068 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1229
timestamp 1636968456
transform 1 0 114172 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_1241
timestamp 1
transform 1 0 115276 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1245
timestamp 1
transform 1 0 115644 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1247
timestamp 1636968456
transform 1 0 115828 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1259
timestamp 1636968456
transform 1 0 116932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_1271
timestamp 1
transform 1 0 118036 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636968456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636968456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636968456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1636968456
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1636968456
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_69
timestamp 1
transform 1 0 7452 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1165
timestamp 1636968456
transform 1 0 108284 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1177
timestamp 1636968456
transform 1 0 109388 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1189
timestamp 1636968456
transform 1 0 110492 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1201
timestamp 1636968456
transform 1 0 111596 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_1213
timestamp 1
transform 1 0 112700 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_1217
timestamp 1
transform 1 0 113068 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1219
timestamp 1636968456
transform 1 0 113252 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1231
timestamp 1636968456
transform 1 0 114356 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1243
timestamp 1636968456
transform 1 0 115460 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1255
timestamp 1636968456
transform 1 0 116564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_1267
timestamp 1
transform 1 0 117668 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_1273
timestamp 1
transform 1 0 118220 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_1275
timestamp 1
transform 1 0 118404 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636968456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636968456
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636968456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1636968456
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1636968456
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_65
timestamp 1
transform 1 0 7084 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_84_1165
timestamp 1
transform 1 0 108284 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_84_1188
timestamp 1
transform 1 0 110400 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1191
timestamp 1636968456
transform 1 0 110676 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1203
timestamp 1636968456
transform 1 0 111780 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1215
timestamp 1636968456
transform 1 0 112884 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1227
timestamp 1636968456
transform 1 0 113988 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_1239
timestamp 1
transform 1 0 115092 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_1245
timestamp 1
transform 1 0 115644 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1247
timestamp 1636968456
transform 1 0 115828 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1259
timestamp 1636968456
transform 1 0 116932 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_1271
timestamp 1
transform 1 0 118036 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1636968456
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1636968456
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1636968456
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1636968456
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1636968456
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_69
timestamp 1
transform 1 0 7452 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1165
timestamp 1636968456
transform 1 0 108284 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1177
timestamp 1636968456
transform 1 0 109388 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1189
timestamp 1636968456
transform 1 0 110492 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1201
timestamp 1636968456
transform 1 0 111596 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_1213
timestamp 1
transform 1 0 112700 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_1217
timestamp 1
transform 1 0 113068 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1219
timestamp 1636968456
transform 1 0 113252 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1231
timestamp 1636968456
transform 1 0 114356 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1243
timestamp 1636968456
transform 1 0 115460 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1255
timestamp 1636968456
transform 1 0 116564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_1267
timestamp 1
transform 1 0 117668 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_1273
timestamp 1
transform 1 0 118220 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_1275
timestamp 1
transform 1 0 118404 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636968456
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636968456
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636968456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1636968456
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1636968456
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_65
timestamp 1
transform 1 0 7084 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_86_1170
timestamp 1
transform 1 0 108744 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1178
timestamp 1636968456
transform 1 0 109480 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1191
timestamp 1636968456
transform 1 0 110676 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1203
timestamp 1636968456
transform 1 0 111780 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1215
timestamp 1636968456
transform 1 0 112884 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1227
timestamp 1636968456
transform 1 0 113988 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_1239
timestamp 1
transform 1 0 115092 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_1245
timestamp 1
transform 1 0 115644 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1247
timestamp 1636968456
transform 1 0 115828 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1259
timestamp 1636968456
transform 1 0 116932 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_1271
timestamp 1
transform 1 0 118036 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636968456
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636968456
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1636968456
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1636968456
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1636968456
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_69
timestamp 1
transform 1 0 7452 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1165
timestamp 1636968456
transform 1 0 108284 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1177
timestamp 1636968456
transform 1 0 109388 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1189
timestamp 1636968456
transform 1 0 110492 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1201
timestamp 1636968456
transform 1 0 111596 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_1213
timestamp 1
transform 1 0 112700 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_1217
timestamp 1
transform 1 0 113068 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1219
timestamp 1636968456
transform 1 0 113252 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1231
timestamp 1636968456
transform 1 0 114356 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1243
timestamp 1636968456
transform 1 0 115460 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1255
timestamp 1636968456
transform 1 0 116564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_1267
timestamp 1
transform 1 0 117668 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_1273
timestamp 1
transform 1 0 118220 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_1275
timestamp 1
transform 1 0 118404 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636968456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636968456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636968456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1636968456
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1636968456
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_65
timestamp 1
transform 1 0 7084 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1170
timestamp 1636968456
transform 1 0 108744 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_1182
timestamp 1
transform 1 0 109848 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1191
timestamp 1636968456
transform 1 0 110676 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1203
timestamp 1636968456
transform 1 0 111780 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1215
timestamp 1636968456
transform 1 0 112884 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1227
timestamp 1636968456
transform 1 0 113988 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_1239
timestamp 1
transform 1 0 115092 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_1245
timestamp 1
transform 1 0 115644 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1247
timestamp 1636968456
transform 1 0 115828 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1259
timestamp 1636968456
transform 1 0 116932 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_1271
timestamp 1
transform 1 0 118036 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636968456
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636968456
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1636968456
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1636968456
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1636968456
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_69
timestamp 1
transform 1 0 7452 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1176
timestamp 1636968456
transform 1 0 109296 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1188
timestamp 1636968456
transform 1 0 110400 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1200
timestamp 1636968456
transform 1 0 111504 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_1212
timestamp 1
transform 1 0 112608 0 -1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1219
timestamp 1636968456
transform 1 0 113252 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1231
timestamp 1636968456
transform 1 0 114356 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1243
timestamp 1636968456
transform 1 0 115460 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1255
timestamp 1636968456
transform 1 0 116564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_1267
timestamp 1
transform 1 0 117668 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_1273
timestamp 1
transform 1 0 118220 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_1275
timestamp 1
transform 1 0 118404 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1636968456
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1636968456
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636968456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1636968456
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1636968456
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_65
timestamp 1
transform 1 0 7084 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_1185
timestamp 1
transform 1 0 110124 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_1189
timestamp 1
transform 1 0 110492 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1191
timestamp 1636968456
transform 1 0 110676 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1203
timestamp 1636968456
transform 1 0 111780 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1215
timestamp 1636968456
transform 1 0 112884 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1227
timestamp 1636968456
transform 1 0 113988 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_1239
timestamp 1
transform 1 0 115092 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_1245
timestamp 1
transform 1 0 115644 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1247
timestamp 1636968456
transform 1 0 115828 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1259
timestamp 1636968456
transform 1 0 116932 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_1271
timestamp 1
transform 1 0 118036 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636968456
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636968456
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1636968456
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1636968456
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1636968456
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_69
timestamp 1
transform 1 0 7452 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_91_1167
timestamp 1
transform 1 0 108468 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1181
timestamp 1636968456
transform 1 0 109756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1193
timestamp 1636968456
transform 1 0 110860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1205
timestamp 1636968456
transform 1 0 111964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_1217
timestamp 1
transform 1 0 113068 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1219
timestamp 1636968456
transform 1 0 113252 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1231
timestamp 1636968456
transform 1 0 114356 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1243
timestamp 1636968456
transform 1 0 115460 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1255
timestamp 1636968456
transform 1 0 116564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_1267
timestamp 1
transform 1 0 117668 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_1273
timestamp 1
transform 1 0 118220 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_1275
timestamp 1
transform 1 0 118404 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1636968456
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1636968456
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636968456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1636968456
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1636968456
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_65
timestamp 1
transform 1 0 7084 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1191
timestamp 1636968456
transform 1 0 110676 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1203
timestamp 1636968456
transform 1 0 111780 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1215
timestamp 1636968456
transform 1 0 112884 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1227
timestamp 1636968456
transform 1 0 113988 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_1239
timestamp 1
transform 1 0 115092 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_1245
timestamp 1
transform 1 0 115644 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1247
timestamp 1636968456
transform 1 0 115828 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1259
timestamp 1636968456
transform 1 0 116932 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_1271
timestamp 1
transform 1 0 118036 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636968456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636968456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636968456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1636968456
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1636968456
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_69
timestamp 1
transform 1 0 7452 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1174
timestamp 1636968456
transform 1 0 109112 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1186
timestamp 1636968456
transform 1 0 110216 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1198
timestamp 1636968456
transform 1 0 111320 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_1210
timestamp 1
transform 1 0 112424 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1219
timestamp 1636968456
transform 1 0 113252 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1231
timestamp 1636968456
transform 1 0 114356 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1243
timestamp 1636968456
transform 1 0 115460 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1255
timestamp 1636968456
transform 1 0 116564 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_1267
timestamp 1
transform 1 0 117668 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_1273
timestamp 1
transform 1 0 118220 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_1275
timestamp 1
transform 1 0 118404 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636968456
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636968456
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636968456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1636968456
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1636968456
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_65
timestamp 1
transform 1 0 7084 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_94_1187
timestamp 1
transform 1 0 110308 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1191
timestamp 1636968456
transform 1 0 110676 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1203
timestamp 1636968456
transform 1 0 111780 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1215
timestamp 1636968456
transform 1 0 112884 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1227
timestamp 1636968456
transform 1 0 113988 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_1239
timestamp 1
transform 1 0 115092 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_1245
timestamp 1
transform 1 0 115644 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1247
timestamp 1636968456
transform 1 0 115828 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1259
timestamp 1636968456
transform 1 0 116932 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_1271
timestamp 1
transform 1 0 118036 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1636968456
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1636968456
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1636968456
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1636968456
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1636968456
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_69
timestamp 1
transform 1 0 7452 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1167
timestamp 1636968456
transform 1 0 108468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1179
timestamp 1636968456
transform 1 0 109572 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1191
timestamp 1636968456
transform 1 0 110676 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1203
timestamp 1636968456
transform 1 0 111780 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_1215
timestamp 1
transform 1 0 112884 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1219
timestamp 1636968456
transform 1 0 113252 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1231
timestamp 1636968456
transform 1 0 114356 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1243
timestamp 1636968456
transform 1 0 115460 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1255
timestamp 1636968456
transform 1 0 116564 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_1267
timestamp 1
transform 1 0 117668 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_1273
timestamp 1
transform 1 0 118220 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_1275
timestamp 1
transform 1 0 118404 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636968456
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636968456
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636968456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1636968456
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1636968456
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_65
timestamp 1
transform 1 0 7084 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1170
timestamp 1636968456
transform 1 0 108744 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_1182
timestamp 1
transform 1 0 109848 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1191
timestamp 1636968456
transform 1 0 110676 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1203
timestamp 1636968456
transform 1 0 111780 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1215
timestamp 1636968456
transform 1 0 112884 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1227
timestamp 1636968456
transform 1 0 113988 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_1239
timestamp 1
transform 1 0 115092 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_1245
timestamp 1
transform 1 0 115644 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1247
timestamp 1636968456
transform 1 0 115828 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1259
timestamp 1636968456
transform 1 0 116932 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_1271
timestamp 1
transform 1 0 118036 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636968456
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636968456
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1636968456
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1636968456
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1636968456
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_69
timestamp 1
transform 1 0 7452 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1165
timestamp 1636968456
transform 1 0 108284 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1177
timestamp 1636968456
transform 1 0 109388 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1189
timestamp 1636968456
transform 1 0 110492 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1201
timestamp 1636968456
transform 1 0 111596 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_1213
timestamp 1
transform 1 0 112700 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_1217
timestamp 1
transform 1 0 113068 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1219
timestamp 1636968456
transform 1 0 113252 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1231
timestamp 1636968456
transform 1 0 114356 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1243
timestamp 1636968456
transform 1 0 115460 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1255
timestamp 1636968456
transform 1 0 116564 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_1267
timestamp 1
transform 1 0 117668 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_1273
timestamp 1
transform 1 0 118220 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_1275
timestamp 1
transform 1 0 118404 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636968456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636968456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636968456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1636968456
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1636968456
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_65
timestamp 1
transform 1 0 7084 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1165
timestamp 1636968456
transform 1 0 108284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1177
timestamp 1636968456
transform 1 0 109388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_1189
timestamp 1
transform 1 0 110492 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1191
timestamp 1636968456
transform 1 0 110676 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1203
timestamp 1636968456
transform 1 0 111780 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1215
timestamp 1636968456
transform 1 0 112884 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1227
timestamp 1636968456
transform 1 0 113988 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_1239
timestamp 1
transform 1 0 115092 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_1245
timestamp 1
transform 1 0 115644 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1247
timestamp 1636968456
transform 1 0 115828 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1259
timestamp 1636968456
transform 1 0 116932 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_1271
timestamp 1
transform 1 0 118036 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636968456
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636968456
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1636968456
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1636968456
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1636968456
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_69
timestamp 1
transform 1 0 7452 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1165
timestamp 1636968456
transform 1 0 108284 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1177
timestamp 1636968456
transform 1 0 109388 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1189
timestamp 1636968456
transform 1 0 110492 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1201
timestamp 1636968456
transform 1 0 111596 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_1213
timestamp 1
transform 1 0 112700 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_1217
timestamp 1
transform 1 0 113068 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1219
timestamp 1636968456
transform 1 0 113252 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1231
timestamp 1636968456
transform 1 0 114356 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1243
timestamp 1636968456
transform 1 0 115460 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1255
timestamp 1636968456
transform 1 0 116564 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_1267
timestamp 1
transform 1 0 117668 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_1273
timestamp 1
transform 1 0 118220 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_1275
timestamp 1
transform 1 0 118404 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1636968456
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1636968456
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1636968456
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1636968456
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1636968456
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_65
timestamp 1
transform 1 0 7084 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1165
timestamp 1636968456
transform 1 0 108284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1177
timestamp 1636968456
transform 1 0 109388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_1189
timestamp 1
transform 1 0 110492 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1191
timestamp 1636968456
transform 1 0 110676 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1203
timestamp 1636968456
transform 1 0 111780 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1215
timestamp 1636968456
transform 1 0 112884 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1227
timestamp 1636968456
transform 1 0 113988 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_1239
timestamp 1
transform 1 0 115092 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_1245
timestamp 1
transform 1 0 115644 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1247
timestamp 1636968456
transform 1 0 115828 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1259
timestamp 1636968456
transform 1 0 116932 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_1271
timestamp 1
transform 1 0 118036 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636968456
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636968456
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_27
timestamp 1636968456
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1636968456
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1636968456
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_69
timestamp 1
transform 1 0 7452 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1165
timestamp 1636968456
transform 1 0 108284 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1177
timestamp 1636968456
transform 1 0 109388 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1189
timestamp 1636968456
transform 1 0 110492 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1201
timestamp 1636968456
transform 1 0 111596 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_1213
timestamp 1
transform 1 0 112700 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_1217
timestamp 1
transform 1 0 113068 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1219
timestamp 1636968456
transform 1 0 113252 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1231
timestamp 1636968456
transform 1 0 114356 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1243
timestamp 1636968456
transform 1 0 115460 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1255
timestamp 1636968456
transform 1 0 116564 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_1267
timestamp 1
transform 1 0 117668 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_1273
timestamp 1
transform 1 0 118220 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_1275
timestamp 1
transform 1 0 118404 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1636968456
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1636968456
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1636968456
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1636968456
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1636968456
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_65
timestamp 1
transform 1 0 7084 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_102_1185
timestamp 1
transform 1 0 110124 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_1189
timestamp 1
transform 1 0 110492 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1191
timestamp 1636968456
transform 1 0 110676 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1203
timestamp 1636968456
transform 1 0 111780 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1215
timestamp 1636968456
transform 1 0 112884 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1227
timestamp 1636968456
transform 1 0 113988 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_1239
timestamp 1
transform 1 0 115092 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_1245
timestamp 1
transform 1 0 115644 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1247
timestamp 1636968456
transform 1 0 115828 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1259
timestamp 1636968456
transform 1 0 116932 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_1271
timestamp 1
transform 1 0 118036 0 1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636968456
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636968456
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1636968456
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_39
timestamp 1636968456
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1636968456
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_69
timestamp 1
transform 1 0 7452 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1165
timestamp 1636968456
transform 1 0 108284 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1177
timestamp 1636968456
transform 1 0 109388 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1189
timestamp 1636968456
transform 1 0 110492 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1201
timestamp 1636968456
transform 1 0 111596 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_1213
timestamp 1
transform 1 0 112700 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_1217
timestamp 1
transform 1 0 113068 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1219
timestamp 1636968456
transform 1 0 113252 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1231
timestamp 1636968456
transform 1 0 114356 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1243
timestamp 1636968456
transform 1 0 115460 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1255
timestamp 1636968456
transform 1 0 116564 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_1267
timestamp 1
transform 1 0 117668 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_1273
timestamp 1
transform 1 0 118220 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_1275
timestamp 1
transform 1 0 118404 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1636968456
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1636968456
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1636968456
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1636968456
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1636968456
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_65
timestamp 1
transform 1 0 7084 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1165
timestamp 1636968456
transform 1 0 108284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1177
timestamp 1636968456
transform 1 0 109388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_1189
timestamp 1
transform 1 0 110492 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1191
timestamp 1636968456
transform 1 0 110676 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1203
timestamp 1636968456
transform 1 0 111780 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1215
timestamp 1636968456
transform 1 0 112884 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1227
timestamp 1636968456
transform 1 0 113988 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_1239
timestamp 1
transform 1 0 115092 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_1245
timestamp 1
transform 1 0 115644 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1247
timestamp 1636968456
transform 1 0 115828 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1259
timestamp 1636968456
transform 1 0 116932 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_1271
timestamp 1
transform 1 0 118036 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_105_3
timestamp 1636968456
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_15
timestamp 1636968456
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_27
timestamp 1636968456
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_39
timestamp 1636968456
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1636968456
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_69
timestamp 1
transform 1 0 7452 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1165
timestamp 1636968456
transform 1 0 108284 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1177
timestamp 1636968456
transform 1 0 109388 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1189
timestamp 1636968456
transform 1 0 110492 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1201
timestamp 1636968456
transform 1 0 111596 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_1213
timestamp 1
transform 1 0 112700 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_1217
timestamp 1
transform 1 0 113068 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1219
timestamp 1636968456
transform 1 0 113252 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1231
timestamp 1636968456
transform 1 0 114356 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1243
timestamp 1636968456
transform 1 0 115460 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1255
timestamp 1636968456
transform 1 0 116564 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_1267
timestamp 1
transform 1 0 117668 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_1273
timestamp 1
transform 1 0 118220 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_1275
timestamp 1
transform 1 0 118404 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636968456
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636968456
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636968456
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1636968456
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1636968456
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_65
timestamp 1
transform 1 0 7084 0 1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1165
timestamp 1636968456
transform 1 0 108284 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1177
timestamp 1636968456
transform 1 0 109388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_1189
timestamp 1
transform 1 0 110492 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1191
timestamp 1636968456
transform 1 0 110676 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1203
timestamp 1636968456
transform 1 0 111780 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1215
timestamp 1636968456
transform 1 0 112884 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1227
timestamp 1636968456
transform 1 0 113988 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_1239
timestamp 1
transform 1 0 115092 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_1245
timestamp 1
transform 1 0 115644 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1247
timestamp 1636968456
transform 1 0 115828 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1259
timestamp 1636968456
transform 1 0 116932 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_1271
timestamp 1
transform 1 0 118036 0 1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636968456
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636968456
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1636968456
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_39
timestamp 1636968456
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1636968456
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_69
timestamp 1
transform 1 0 7452 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1165
timestamp 1636968456
transform 1 0 108284 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1177
timestamp 1636968456
transform 1 0 109388 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1189
timestamp 1636968456
transform 1 0 110492 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1201
timestamp 1636968456
transform 1 0 111596 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_1213
timestamp 1
transform 1 0 112700 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_1217
timestamp 1
transform 1 0 113068 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1219
timestamp 1636968456
transform 1 0 113252 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1231
timestamp 1636968456
transform 1 0 114356 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1243
timestamp 1636968456
transform 1 0 115460 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1255
timestamp 1636968456
transform 1 0 116564 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_1267
timestamp 1
transform 1 0 117668 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_1273
timestamp 1
transform 1 0 118220 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_107_1275
timestamp 1
transform 1 0 118404 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636968456
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636968456
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636968456
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1636968456
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1636968456
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_65
timestamp 1
transform 1 0 7084 0 1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1165
timestamp 1636968456
transform 1 0 108284 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1177
timestamp 1636968456
transform 1 0 109388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_1189
timestamp 1
transform 1 0 110492 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1191
timestamp 1636968456
transform 1 0 110676 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1203
timestamp 1636968456
transform 1 0 111780 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1215
timestamp 1636968456
transform 1 0 112884 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1227
timestamp 1636968456
transform 1 0 113988 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_1239
timestamp 1
transform 1 0 115092 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_1245
timestamp 1
transform 1 0 115644 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1247
timestamp 1636968456
transform 1 0 115828 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1259
timestamp 1636968456
transform 1 0 116932 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_1271
timestamp 1
transform 1 0 118036 0 1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1636968456
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1636968456
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_27
timestamp 1636968456
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_39
timestamp 1636968456
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1636968456
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_69
timestamp 1
transform 1 0 7452 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1165
timestamp 1636968456
transform 1 0 108284 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1177
timestamp 1636968456
transform 1 0 109388 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1189
timestamp 1636968456
transform 1 0 110492 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1201
timestamp 1636968456
transform 1 0 111596 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_1213
timestamp 1
transform 1 0 112700 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_1217
timestamp 1
transform 1 0 113068 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1219
timestamp 1636968456
transform 1 0 113252 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1231
timestamp 1636968456
transform 1 0 114356 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1243
timestamp 1636968456
transform 1 0 115460 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1255
timestamp 1636968456
transform 1 0 116564 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_1267
timestamp 1
transform 1 0 117668 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_1273
timestamp 1
transform 1 0 118220 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_109_1275
timestamp 1
transform 1 0 118404 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_110_3
timestamp 1636968456
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_15
timestamp 1636968456
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636968456
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1636968456
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1636968456
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_65
timestamp 1
transform 1 0 7084 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1165
timestamp 1636968456
transform 1 0 108284 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1177
timestamp 1636968456
transform 1 0 109388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_1189
timestamp 1
transform 1 0 110492 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1191
timestamp 1636968456
transform 1 0 110676 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1203
timestamp 1636968456
transform 1 0 111780 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1215
timestamp 1636968456
transform 1 0 112884 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1227
timestamp 1636968456
transform 1 0 113988 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_1239
timestamp 1
transform 1 0 115092 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_1245
timestamp 1
transform 1 0 115644 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1247
timestamp 1636968456
transform 1 0 115828 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1259
timestamp 1636968456
transform 1 0 116932 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_1271
timestamp 1
transform 1 0 118036 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636968456
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636968456
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1636968456
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_39
timestamp 1636968456
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1636968456
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_69
timestamp 1
transform 1 0 7452 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1165
timestamp 1636968456
transform 1 0 108284 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1177
timestamp 1636968456
transform 1 0 109388 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1189
timestamp 1636968456
transform 1 0 110492 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1201
timestamp 1636968456
transform 1 0 111596 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_1213
timestamp 1
transform 1 0 112700 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_1217
timestamp 1
transform 1 0 113068 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1219
timestamp 1636968456
transform 1 0 113252 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1231
timestamp 1636968456
transform 1 0 114356 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1243
timestamp 1636968456
transform 1 0 115460 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1255
timestamp 1636968456
transform 1 0 116564 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_1267
timestamp 1
transform 1 0 117668 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_1273
timestamp 1
transform 1 0 118220 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_111_1275
timestamp 1
transform 1 0 118404 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1636968456
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1636968456
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636968456
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1636968456
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1636968456
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_65
timestamp 1
transform 1 0 7084 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1165
timestamp 1636968456
transform 1 0 108284 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1177
timestamp 1636968456
transform 1 0 109388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_1189
timestamp 1
transform 1 0 110492 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1191
timestamp 1636968456
transform 1 0 110676 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1203
timestamp 1636968456
transform 1 0 111780 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1215
timestamp 1636968456
transform 1 0 112884 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1227
timestamp 1636968456
transform 1 0 113988 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_1239
timestamp 1
transform 1 0 115092 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_1245
timestamp 1
transform 1 0 115644 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1247
timestamp 1636968456
transform 1 0 115828 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1259
timestamp 1636968456
transform 1 0 116932 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_1271
timestamp 1
transform 1 0 118036 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636968456
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636968456
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636968456
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1636968456
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1636968456
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_69
timestamp 1
transform 1 0 7452 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1165
timestamp 1636968456
transform 1 0 108284 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1177
timestamp 1636968456
transform 1 0 109388 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1189
timestamp 1636968456
transform 1 0 110492 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1201
timestamp 1636968456
transform 1 0 111596 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_1213
timestamp 1
transform 1 0 112700 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_1217
timestamp 1
transform 1 0 113068 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1219
timestamp 1636968456
transform 1 0 113252 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1231
timestamp 1636968456
transform 1 0 114356 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1243
timestamp 1636968456
transform 1 0 115460 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1255
timestamp 1636968456
transform 1 0 116564 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_1267
timestamp 1
transform 1 0 117668 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_1273
timestamp 1
transform 1 0 118220 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_113_1275
timestamp 1
transform 1 0 118404 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636968456
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636968456
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636968456
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1636968456
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1636968456
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_65
timestamp 1
transform 1 0 7084 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1165
timestamp 1636968456
transform 1 0 108284 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1177
timestamp 1636968456
transform 1 0 109388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_1189
timestamp 1
transform 1 0 110492 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1191
timestamp 1636968456
transform 1 0 110676 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1203
timestamp 1636968456
transform 1 0 111780 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1215
timestamp 1636968456
transform 1 0 112884 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1227
timestamp 1636968456
transform 1 0 113988 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_1239
timestamp 1
transform 1 0 115092 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_1245
timestamp 1
transform 1 0 115644 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1247
timestamp 1636968456
transform 1 0 115828 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1259
timestamp 1636968456
transform 1 0 116932 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_1271
timestamp 1
transform 1 0 118036 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_115_3
timestamp 1636968456
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_15
timestamp 1636968456
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_27
timestamp 1636968456
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_39
timestamp 1636968456
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1636968456
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_115_69
timestamp 1
transform 1 0 7452 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1165
timestamp 1636968456
transform 1 0 108284 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1177
timestamp 1636968456
transform 1 0 109388 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1189
timestamp 1636968456
transform 1 0 110492 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1201
timestamp 1636968456
transform 1 0 111596 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_1213
timestamp 1
transform 1 0 112700 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_1217
timestamp 1
transform 1 0 113068 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1219
timestamp 1636968456
transform 1 0 113252 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1231
timestamp 1636968456
transform 1 0 114356 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1243
timestamp 1636968456
transform 1 0 115460 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1255
timestamp 1636968456
transform 1 0 116564 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_1267
timestamp 1
transform 1 0 117668 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_1273
timestamp 1
transform 1 0 118220 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_115_1275
timestamp 1
transform 1 0 118404 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636968456
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636968456
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636968456
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1636968456
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_53
timestamp 1636968456
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_65
timestamp 1
transform 1 0 7084 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1165
timestamp 1636968456
transform 1 0 108284 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1177
timestamp 1636968456
transform 1 0 109388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_1189
timestamp 1
transform 1 0 110492 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1191
timestamp 1636968456
transform 1 0 110676 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1203
timestamp 1636968456
transform 1 0 111780 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1215
timestamp 1636968456
transform 1 0 112884 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1227
timestamp 1636968456
transform 1 0 113988 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_1239
timestamp 1
transform 1 0 115092 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_1245
timestamp 1
transform 1 0 115644 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1247
timestamp 1636968456
transform 1 0 115828 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1259
timestamp 1636968456
transform 1 0 116932 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_1271
timestamp 1
transform 1 0 118036 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636968456
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636968456
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_27
timestamp 1636968456
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_39
timestamp 1636968456
transform 1 0 4692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_51
timestamp 1
transform 1 0 5796 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1636968456
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_69
timestamp 1
transform 1 0 7452 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1165
timestamp 1636968456
transform 1 0 108284 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1177
timestamp 1636968456
transform 1 0 109388 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1189
timestamp 1636968456
transform 1 0 110492 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1201
timestamp 1636968456
transform 1 0 111596 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_1213
timestamp 1
transform 1 0 112700 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1217
timestamp 1
transform 1 0 113068 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1219
timestamp 1636968456
transform 1 0 113252 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1231
timestamp 1636968456
transform 1 0 114356 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1243
timestamp 1636968456
transform 1 0 115460 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1255
timestamp 1636968456
transform 1 0 116564 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_1267
timestamp 1
transform 1 0 117668 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1273
timestamp 1
transform 1 0 118220 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_117_1275
timestamp 1
transform 1 0 118404 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636968456
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636968456
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636968456
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1636968456
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1636968456
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_65
timestamp 1
transform 1 0 7084 0 1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1165
timestamp 1636968456
transform 1 0 108284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1177
timestamp 1636968456
transform 1 0 109388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1189
timestamp 1
transform 1 0 110492 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1191
timestamp 1636968456
transform 1 0 110676 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1203
timestamp 1636968456
transform 1 0 111780 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1215
timestamp 1636968456
transform 1 0 112884 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1227
timestamp 1636968456
transform 1 0 113988 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1239
timestamp 1
transform 1 0 115092 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1245
timestamp 1
transform 1 0 115644 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1247
timestamp 1636968456
transform 1 0 115828 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1259
timestamp 1636968456
transform 1 0 116932 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1271
timestamp 1
transform 1 0 118036 0 1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636968456
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636968456
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1636968456
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_39
timestamp 1636968456
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1636968456
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_69
timestamp 1
transform 1 0 7452 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1186
timestamp 1636968456
transform 1 0 110216 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1198
timestamp 1636968456
transform 1 0 111320 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_1210
timestamp 1
transform 1 0 112424 0 -1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1219
timestamp 1636968456
transform 1 0 113252 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1231
timestamp 1636968456
transform 1 0 114356 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1243
timestamp 1636968456
transform 1 0 115460 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1255
timestamp 1636968456
transform 1 0 116564 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1267
timestamp 1
transform 1 0 117668 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1273
timestamp 1
transform 1 0 118220 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_119_1275
timestamp 1
transform 1 0 118404 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1636968456
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1636968456
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636968456
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1636968456
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1636968456
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_65
timestamp 1
transform 1 0 7084 0 1 67456
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1165
timestamp 1636968456
transform 1 0 108284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1177
timestamp 1636968456
transform 1 0 109388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1189
timestamp 1
transform 1 0 110492 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1191
timestamp 1636968456
transform 1 0 110676 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1203
timestamp 1636968456
transform 1 0 111780 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1215
timestamp 1636968456
transform 1 0 112884 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1227
timestamp 1636968456
transform 1 0 113988 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1239
timestamp 1
transform 1 0 115092 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1245
timestamp 1
transform 1 0 115644 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1247
timestamp 1636968456
transform 1 0 115828 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1259
timestamp 1636968456
transform 1 0 116932 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1271
timestamp 1
transform 1 0 118036 0 1 67456
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636968456
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636968456
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1636968456
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_39
timestamp 1636968456
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1636968456
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_69
timestamp 1
transform 1 0 7452 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1165
timestamp 1636968456
transform 1 0 108284 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1177
timestamp 1636968456
transform 1 0 109388 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1189
timestamp 1636968456
transform 1 0 110492 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1201
timestamp 1636968456
transform 1 0 111596 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_1213
timestamp 1
transform 1 0 112700 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1217
timestamp 1
transform 1 0 113068 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1219
timestamp 1636968456
transform 1 0 113252 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1231
timestamp 1636968456
transform 1 0 114356 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1243
timestamp 1636968456
transform 1 0 115460 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1255
timestamp 1636968456
transform 1 0 116564 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1267
timestamp 1
transform 1 0 117668 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1273
timestamp 1
transform 1 0 118220 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_121_1275
timestamp 1
transform 1 0 118404 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1636968456
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1636968456
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636968456
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1636968456
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1636968456
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_65
timestamp 1
transform 1 0 7084 0 1 68544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1165
timestamp 1636968456
transform 1 0 108284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1177
timestamp 1636968456
transform 1 0 109388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1189
timestamp 1
transform 1 0 110492 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1191
timestamp 1636968456
transform 1 0 110676 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1203
timestamp 1636968456
transform 1 0 111780 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1215
timestamp 1636968456
transform 1 0 112884 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1227
timestamp 1636968456
transform 1 0 113988 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1239
timestamp 1
transform 1 0 115092 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1245
timestamp 1
transform 1 0 115644 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1247
timestamp 1636968456
transform 1 0 115828 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1259
timestamp 1636968456
transform 1 0 116932 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1271
timestamp 1
transform 1 0 118036 0 1 68544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636968456
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636968456
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636968456
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_39
timestamp 1636968456
transform 1 0 4692 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1
transform 1 0 5796 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1636968456
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_69
timestamp 1
transform 1 0 7452 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1165
timestamp 1636968456
transform 1 0 108284 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1177
timestamp 1636968456
transform 1 0 109388 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1189
timestamp 1636968456
transform 1 0 110492 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1201
timestamp 1636968456
transform 1 0 111596 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_1213
timestamp 1
transform 1 0 112700 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1217
timestamp 1
transform 1 0 113068 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1219
timestamp 1636968456
transform 1 0 113252 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1231
timestamp 1636968456
transform 1 0 114356 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1243
timestamp 1636968456
transform 1 0 115460 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1255
timestamp 1636968456
transform 1 0 116564 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1267
timestamp 1
transform 1 0 117668 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1273
timestamp 1
transform 1 0 118220 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_123_1275
timestamp 1
transform 1 0 118404 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636968456
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636968456
transform 1 0 2484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 1
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1636968456
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_41
timestamp 1636968456
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_53
timestamp 1636968456
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_65
timestamp 1
transform 1 0 7084 0 1 69632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1165
timestamp 1636968456
transform 1 0 108284 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1177
timestamp 1636968456
transform 1 0 109388 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1189
timestamp 1
transform 1 0 110492 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1191
timestamp 1636968456
transform 1 0 110676 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1203
timestamp 1636968456
transform 1 0 111780 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1215
timestamp 1636968456
transform 1 0 112884 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1227
timestamp 1636968456
transform 1 0 113988 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1239
timestamp 1
transform 1 0 115092 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1245
timestamp 1
transform 1 0 115644 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1247
timestamp 1636968456
transform 1 0 115828 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1259
timestamp 1636968456
transform 1 0 116932 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1271
timestamp 1
transform 1 0 118036 0 1 69632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_125_3
timestamp 1636968456
transform 1 0 1380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_15
timestamp 1636968456
transform 1 0 2484 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_27
timestamp 1636968456
transform 1 0 3588 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_39
timestamp 1636968456
transform 1 0 4692 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1
transform 1 0 5796 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1636968456
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_125_69
timestamp 1
transform 1 0 7452 0 -1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1165
timestamp 1636968456
transform 1 0 108284 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1177
timestamp 1636968456
transform 1 0 109388 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1189
timestamp 1636968456
transform 1 0 110492 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1201
timestamp 1636968456
transform 1 0 111596 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_1213
timestamp 1
transform 1 0 112700 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1217
timestamp 1
transform 1 0 113068 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1219
timestamp 1636968456
transform 1 0 113252 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1231
timestamp 1636968456
transform 1 0 114356 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1243
timestamp 1636968456
transform 1 0 115460 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1255
timestamp 1636968456
transform 1 0 116564 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1267
timestamp 1
transform 1 0 117668 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1273
timestamp 1
transform 1 0 118220 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_125_1275
timestamp 1
transform 1 0 118404 0 -1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636968456
transform 1 0 1380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636968456
transform 1 0 2484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 1
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636968456
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1636968456
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_53
timestamp 1636968456
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_65
timestamp 1
transform 1 0 7084 0 1 70720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1165
timestamp 1636968456
transform 1 0 108284 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1177
timestamp 1636968456
transform 1 0 109388 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1189
timestamp 1
transform 1 0 110492 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1191
timestamp 1636968456
transform 1 0 110676 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1203
timestamp 1636968456
transform 1 0 111780 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1215
timestamp 1636968456
transform 1 0 112884 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1227
timestamp 1636968456
transform 1 0 113988 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1239
timestamp 1
transform 1 0 115092 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1245
timestamp 1
transform 1 0 115644 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1247
timestamp 1636968456
transform 1 0 115828 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1259
timestamp 1636968456
transform 1 0 116932 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1271
timestamp 1
transform 1 0 118036 0 1 70720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1636968456
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1636968456
transform 1 0 2484 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_27
timestamp 1636968456
transform 1 0 3588 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_39
timestamp 1636968456
transform 1 0 4692 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_51
timestamp 1
transform 1 0 5796 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1636968456
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_69
timestamp 1
transform 1 0 7452 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1165
timestamp 1636968456
transform 1 0 108284 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1177
timestamp 1636968456
transform 1 0 109388 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1189
timestamp 1636968456
transform 1 0 110492 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1201
timestamp 1636968456
transform 1 0 111596 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_1213
timestamp 1
transform 1 0 112700 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1217
timestamp 1
transform 1 0 113068 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1219
timestamp 1636968456
transform 1 0 113252 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1231
timestamp 1636968456
transform 1 0 114356 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1243
timestamp 1636968456
transform 1 0 115460 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1255
timestamp 1636968456
transform 1 0 116564 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_1267
timestamp 1
transform 1 0 117668 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1273
timestamp 1
transform 1 0 118220 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_127_1275
timestamp 1
transform 1 0 118404 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636968456
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636968456
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1636968456
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_41
timestamp 1636968456
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_53
timestamp 1636968456
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_65
timestamp 1
transform 1 0 7084 0 1 71808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1165
timestamp 1636968456
transform 1 0 108284 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1177
timestamp 1636968456
transform 1 0 109388 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1189
timestamp 1
transform 1 0 110492 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1191
timestamp 1636968456
transform 1 0 110676 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1203
timestamp 1636968456
transform 1 0 111780 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1215
timestamp 1636968456
transform 1 0 112884 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1227
timestamp 1636968456
transform 1 0 113988 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_1239
timestamp 1
transform 1 0 115092 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1245
timestamp 1
transform 1 0 115644 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1247
timestamp 1636968456
transform 1 0 115828 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1259
timestamp 1636968456
transform 1 0 116932 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_1271
timestamp 1
transform 1 0 118036 0 1 71808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_129_3
timestamp 1636968456
transform 1 0 1380 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_15
timestamp 1636968456
transform 1 0 2484 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_27
timestamp 1636968456
transform 1 0 3588 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_39
timestamp 1636968456
transform 1 0 4692 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_51
timestamp 1
transform 1 0 5796 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_57
timestamp 1636968456
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_69
timestamp 1
transform 1 0 7452 0 -1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1165
timestamp 1636968456
transform 1 0 108284 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1177
timestamp 1636968456
transform 1 0 109388 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1189
timestamp 1636968456
transform 1 0 110492 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1201
timestamp 1636968456
transform 1 0 111596 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_1213
timestamp 1
transform 1 0 112700 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1217
timestamp 1
transform 1 0 113068 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1219
timestamp 1636968456
transform 1 0 113252 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1231
timestamp 1636968456
transform 1 0 114356 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1243
timestamp 1636968456
transform 1 0 115460 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1255
timestamp 1636968456
transform 1 0 116564 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_1267
timestamp 1
transform 1 0 117668 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1273
timestamp 1
transform 1 0 118220 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_129_1275
timestamp 1
transform 1 0 118404 0 -1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_130_3
timestamp 1636968456
transform 1 0 1380 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_15
timestamp 1636968456
transform 1 0 2484 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1636968456
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_41
timestamp 1636968456
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_53
timestamp 1636968456
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_65
timestamp 1
transform 1 0 7084 0 1 72896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1165
timestamp 1636968456
transform 1 0 108284 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1177
timestamp 1636968456
transform 1 0 109388 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1189
timestamp 1
transform 1 0 110492 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1191
timestamp 1636968456
transform 1 0 110676 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1203
timestamp 1636968456
transform 1 0 111780 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1215
timestamp 1636968456
transform 1 0 112884 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1227
timestamp 1636968456
transform 1 0 113988 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_1239
timestamp 1
transform 1 0 115092 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1245
timestamp 1
transform 1 0 115644 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1247
timestamp 1636968456
transform 1 0 115828 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1259
timestamp 1636968456
transform 1 0 116932 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_1271
timestamp 1
transform 1 0 118036 0 1 72896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_131_3
timestamp 1636968456
transform 1 0 1380 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_15
timestamp 1636968456
transform 1 0 2484 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_27
timestamp 1636968456
transform 1 0 3588 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_39
timestamp 1636968456
transform 1 0 4692 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_51
timestamp 1
transform 1 0 5796 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_57
timestamp 1636968456
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_69
timestamp 1
transform 1 0 7452 0 -1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1165
timestamp 1636968456
transform 1 0 108284 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1177
timestamp 1636968456
transform 1 0 109388 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1189
timestamp 1636968456
transform 1 0 110492 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1201
timestamp 1636968456
transform 1 0 111596 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_1213
timestamp 1
transform 1 0 112700 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1217
timestamp 1
transform 1 0 113068 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1219
timestamp 1636968456
transform 1 0 113252 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1231
timestamp 1636968456
transform 1 0 114356 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1243
timestamp 1636968456
transform 1 0 115460 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1255
timestamp 1636968456
transform 1 0 116564 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1267
timestamp 1
transform 1 0 117668 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1273
timestamp 1
transform 1 0 118220 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_131_1275
timestamp 1
transform 1 0 118404 0 -1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_132_3
timestamp 1636968456
transform 1 0 1380 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_15
timestamp 1636968456
transform 1 0 2484 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1636968456
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_41
timestamp 1636968456
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_53
timestamp 1636968456
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_65
timestamp 1
transform 1 0 7084 0 1 73984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1165
timestamp 1636968456
transform 1 0 108284 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1177
timestamp 1636968456
transform 1 0 109388 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1189
timestamp 1
transform 1 0 110492 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1191
timestamp 1636968456
transform 1 0 110676 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1203
timestamp 1636968456
transform 1 0 111780 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1215
timestamp 1636968456
transform 1 0 112884 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1227
timestamp 1636968456
transform 1 0 113988 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_1239
timestamp 1
transform 1 0 115092 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1245
timestamp 1
transform 1 0 115644 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1247
timestamp 1636968456
transform 1 0 115828 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1259
timestamp 1636968456
transform 1 0 116932 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_1271
timestamp 1
transform 1 0 118036 0 1 73984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636968456
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636968456
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1636968456
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_39
timestamp 1636968456
transform 1 0 4692 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_51
timestamp 1
transform 1 0 5796 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_55
timestamp 1
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_57
timestamp 1636968456
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_69
timestamp 1
transform 1 0 7452 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1165
timestamp 1636968456
transform 1 0 108284 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1177
timestamp 1636968456
transform 1 0 109388 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1189
timestamp 1636968456
transform 1 0 110492 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1201
timestamp 1636968456
transform 1 0 111596 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_1213
timestamp 1
transform 1 0 112700 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1217
timestamp 1
transform 1 0 113068 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1219
timestamp 1636968456
transform 1 0 113252 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1231
timestamp 1636968456
transform 1 0 114356 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1243
timestamp 1636968456
transform 1 0 115460 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1255
timestamp 1636968456
transform 1 0 116564 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_1267
timestamp 1
transform 1 0 117668 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1273
timestamp 1
transform 1 0 118220 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_133_1275
timestamp 1
transform 1 0 118404 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_134_3
timestamp 1636968456
transform 1 0 1380 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_15
timestamp 1636968456
transform 1 0 2484 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1636968456
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_41
timestamp 1636968456
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_53
timestamp 1636968456
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_65
timestamp 1
transform 1 0 7084 0 1 75072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1165
timestamp 1636968456
transform 1 0 108284 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1177
timestamp 1636968456
transform 1 0 109388 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1189
timestamp 1
transform 1 0 110492 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1191
timestamp 1636968456
transform 1 0 110676 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1203
timestamp 1636968456
transform 1 0 111780 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1215
timestamp 1636968456
transform 1 0 112884 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1227
timestamp 1636968456
transform 1 0 113988 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_1239
timestamp 1
transform 1 0 115092 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1245
timestamp 1
transform 1 0 115644 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1247
timestamp 1636968456
transform 1 0 115828 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1259
timestamp 1636968456
transform 1 0 116932 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_1271
timestamp 1
transform 1 0 118036 0 1 75072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_135_3
timestamp 1636968456
transform 1 0 1380 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_15
timestamp 1636968456
transform 1 0 2484 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_27
timestamp 1636968456
transform 1 0 3588 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_39
timestamp 1636968456
transform 1 0 4692 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_51
timestamp 1
transform 1 0 5796 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_55
timestamp 1
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_57
timestamp 1636968456
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_135_69
timestamp 1
transform 1 0 7452 0 -1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1165
timestamp 1636968456
transform 1 0 108284 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1177
timestamp 1636968456
transform 1 0 109388 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1189
timestamp 1636968456
transform 1 0 110492 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1201
timestamp 1636968456
transform 1 0 111596 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_1213
timestamp 1
transform 1 0 112700 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1217
timestamp 1
transform 1 0 113068 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1219
timestamp 1636968456
transform 1 0 113252 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1231
timestamp 1636968456
transform 1 0 114356 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1243
timestamp 1636968456
transform 1 0 115460 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1255
timestamp 1636968456
transform 1 0 116564 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1267
timestamp 1
transform 1 0 117668 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1273
timestamp 1
transform 1 0 118220 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_135_1275
timestamp 1
transform 1 0 118404 0 -1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1636968456
transform 1 0 1380 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1636968456
transform 1 0 2484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1636968456
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_41
timestamp 1636968456
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_53
timestamp 1636968456
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_65
timestamp 1
transform 1 0 7084 0 1 76160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1165
timestamp 1636968456
transform 1 0 108284 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1177
timestamp 1636968456
transform 1 0 109388 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1189
timestamp 1
transform 1 0 110492 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1191
timestamp 1636968456
transform 1 0 110676 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1203
timestamp 1636968456
transform 1 0 111780 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1215
timestamp 1636968456
transform 1 0 112884 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1227
timestamp 1636968456
transform 1 0 113988 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_1239
timestamp 1
transform 1 0 115092 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1245
timestamp 1
transform 1 0 115644 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1247
timestamp 1636968456
transform 1 0 115828 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1259
timestamp 1636968456
transform 1 0 116932 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_1271
timestamp 1
transform 1 0 118036 0 1 76160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_137_3
timestamp 1636968456
transform 1 0 1380 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_15
timestamp 1636968456
transform 1 0 2484 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_27
timestamp 1636968456
transform 1 0 3588 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_39
timestamp 1636968456
transform 1 0 4692 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_57
timestamp 1636968456
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_137_69
timestamp 1
transform 1 0 7452 0 -1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1165
timestamp 1636968456
transform 1 0 108284 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1177
timestamp 1636968456
transform 1 0 109388 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1189
timestamp 1636968456
transform 1 0 110492 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1201
timestamp 1636968456
transform 1 0 111596 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_1213
timestamp 1
transform 1 0 112700 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1217
timestamp 1
transform 1 0 113068 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1219
timestamp 1636968456
transform 1 0 113252 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1231
timestamp 1636968456
transform 1 0 114356 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1243
timestamp 1636968456
transform 1 0 115460 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1255
timestamp 1636968456
transform 1 0 116564 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_1267
timestamp 1
transform 1 0 117668 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1273
timestamp 1
transform 1 0 118220 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_137_1275
timestamp 1
transform 1 0 118404 0 -1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636968456
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636968456
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1636968456
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_41
timestamp 1636968456
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_53
timestamp 1636968456
transform 1 0 5980 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_65
timestamp 1
transform 1 0 7084 0 1 77248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1165
timestamp 1636968456
transform 1 0 108284 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1177
timestamp 1636968456
transform 1 0 109388 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1189
timestamp 1
transform 1 0 110492 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1191
timestamp 1636968456
transform 1 0 110676 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1203
timestamp 1636968456
transform 1 0 111780 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1215
timestamp 1636968456
transform 1 0 112884 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1227
timestamp 1636968456
transform 1 0 113988 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_1239
timestamp 1
transform 1 0 115092 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1245
timestamp 1
transform 1 0 115644 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1247
timestamp 1636968456
transform 1 0 115828 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1259
timestamp 1636968456
transform 1 0 116932 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_1271
timestamp 1
transform 1 0 118036 0 1 77248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_139_3
timestamp 1636968456
transform 1 0 1380 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_15
timestamp 1636968456
transform 1 0 2484 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_27
timestamp 1636968456
transform 1 0 3588 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_39
timestamp 1636968456
transform 1 0 4692 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_139_51
timestamp 1
transform 1 0 5796 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_139_55
timestamp 1
transform 1 0 6164 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_57
timestamp 1636968456
transform 1 0 6348 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_139_69
timestamp 1
transform 1 0 7452 0 -1 78336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1165
timestamp 1636968456
transform 1 0 108284 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1177
timestamp 1636968456
transform 1 0 109388 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1189
timestamp 1636968456
transform 1 0 110492 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1201
timestamp 1636968456
transform 1 0 111596 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_139_1213
timestamp 1
transform 1 0 112700 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_139_1217
timestamp 1
transform 1 0 113068 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1219
timestamp 1636968456
transform 1 0 113252 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1231
timestamp 1636968456
transform 1 0 114356 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1243
timestamp 1636968456
transform 1 0 115460 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1255
timestamp 1636968456
transform 1 0 116564 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_1267
timestamp 1
transform 1 0 117668 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_1273
timestamp 1
transform 1 0 118220 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_139_1275
timestamp 1
transform 1 0 118404 0 -1 78336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_140_3
timestamp 1636968456
transform 1 0 1380 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_15
timestamp 1636968456
transform 1 0 2484 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 1
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_29
timestamp 1636968456
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_41
timestamp 1636968456
transform 1 0 4876 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_53
timestamp 1636968456
transform 1 0 5980 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_65
timestamp 1
transform 1 0 7084 0 1 78336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1165
timestamp 1636968456
transform 1 0 108284 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1177
timestamp 1636968456
transform 1 0 109388 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_1189
timestamp 1
transform 1 0 110492 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1191
timestamp 1636968456
transform 1 0 110676 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1203
timestamp 1636968456
transform 1 0 111780 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1215
timestamp 1636968456
transform 1 0 112884 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1227
timestamp 1636968456
transform 1 0 113988 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_1239
timestamp 1
transform 1 0 115092 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_1245
timestamp 1
transform 1 0 115644 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1247
timestamp 1636968456
transform 1 0 115828 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1259
timestamp 1636968456
transform 1 0 116932 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_1271
timestamp 1
transform 1 0 118036 0 1 78336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_141_3
timestamp 1636968456
transform 1 0 1380 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_15
timestamp 1636968456
transform 1 0 2484 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_27
timestamp 1636968456
transform 1 0 3588 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_39
timestamp 1636968456
transform 1 0 4692 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_141_51
timestamp 1
transform 1 0 5796 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_141_55
timestamp 1
transform 1 0 6164 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_57
timestamp 1636968456
transform 1 0 6348 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_141_69
timestamp 1
transform 1 0 7452 0 -1 79424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1165
timestamp 1636968456
transform 1 0 108284 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1177
timestamp 1636968456
transform 1 0 109388 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1189
timestamp 1636968456
transform 1 0 110492 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1201
timestamp 1636968456
transform 1 0 111596 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_141_1213
timestamp 1
transform 1 0 112700 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_141_1217
timestamp 1
transform 1 0 113068 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1219
timestamp 1636968456
transform 1 0 113252 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1231
timestamp 1636968456
transform 1 0 114356 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1243
timestamp 1636968456
transform 1 0 115460 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1255
timestamp 1636968456
transform 1 0 116564 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_1267
timestamp 1
transform 1 0 117668 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_1273
timestamp 1
transform 1 0 118220 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_141_1275
timestamp 1
transform 1 0 118404 0 -1 79424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_142_3
timestamp 1636968456
transform 1 0 1380 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_15
timestamp 1636968456
transform 1 0 2484 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 1
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_29
timestamp 1636968456
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_41
timestamp 1636968456
transform 1 0 4876 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_53
timestamp 1636968456
transform 1 0 5980 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_65
timestamp 1
transform 1 0 7084 0 1 79424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1165
timestamp 1636968456
transform 1 0 108284 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1177
timestamp 1636968456
transform 1 0 109388 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_1189
timestamp 1
transform 1 0 110492 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1191
timestamp 1636968456
transform 1 0 110676 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1203
timestamp 1636968456
transform 1 0 111780 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1215
timestamp 1636968456
transform 1 0 112884 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1227
timestamp 1636968456
transform 1 0 113988 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_1239
timestamp 1
transform 1 0 115092 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_1245
timestamp 1
transform 1 0 115644 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1247
timestamp 1636968456
transform 1 0 115828 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1259
timestamp 1636968456
transform 1 0 116932 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_1271
timestamp 1
transform 1 0 118036 0 1 79424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_143_3
timestamp 1636968456
transform 1 0 1380 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_15
timestamp 1636968456
transform 1 0 2484 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_27
timestamp 1636968456
transform 1 0 3588 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_39
timestamp 1636968456
transform 1 0 4692 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_143_51
timestamp 1
transform 1 0 5796 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_143_55
timestamp 1
transform 1 0 6164 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_57
timestamp 1636968456
transform 1 0 6348 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_143_69
timestamp 1
transform 1 0 7452 0 -1 80512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1165
timestamp 1636968456
transform 1 0 108284 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1177
timestamp 1636968456
transform 1 0 109388 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1189
timestamp 1636968456
transform 1 0 110492 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1201
timestamp 1636968456
transform 1 0 111596 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_143_1213
timestamp 1
transform 1 0 112700 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_143_1217
timestamp 1
transform 1 0 113068 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1219
timestamp 1636968456
transform 1 0 113252 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1231
timestamp 1636968456
transform 1 0 114356 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1243
timestamp 1636968456
transform 1 0 115460 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1255
timestamp 1636968456
transform 1 0 116564 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_1267
timestamp 1
transform 1 0 117668 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_1273
timestamp 1
transform 1 0 118220 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_143_1275
timestamp 1
transform 1 0 118404 0 -1 80512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_144_3
timestamp 1636968456
transform 1 0 1380 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636968456
transform 1 0 2484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 1
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_29
timestamp 1636968456
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_41
timestamp 1636968456
transform 1 0 4876 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_53
timestamp 1636968456
transform 1 0 5980 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_65
timestamp 1
transform 1 0 7084 0 1 80512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1165
timestamp 1636968456
transform 1 0 108284 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1177
timestamp 1636968456
transform 1 0 109388 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_1189
timestamp 1
transform 1 0 110492 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1191
timestamp 1636968456
transform 1 0 110676 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1203
timestamp 1636968456
transform 1 0 111780 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1215
timestamp 1636968456
transform 1 0 112884 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1227
timestamp 1636968456
transform 1 0 113988 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_1239
timestamp 1
transform 1 0 115092 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_1245
timestamp 1
transform 1 0 115644 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1247
timestamp 1636968456
transform 1 0 115828 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1259
timestamp 1636968456
transform 1 0 116932 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_1271
timestamp 1
transform 1 0 118036 0 1 80512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_145_3
timestamp 1636968456
transform 1 0 1380 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_15
timestamp 1636968456
transform 1 0 2484 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_27
timestamp 1636968456
transform 1 0 3588 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_39
timestamp 1636968456
transform 1 0 4692 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_145_51
timestamp 1
transform 1 0 5796 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_145_55
timestamp 1
transform 1 0 6164 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_57
timestamp 1636968456
transform 1 0 6348 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_145_69
timestamp 1
transform 1 0 7452 0 -1 81600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1165
timestamp 1636968456
transform 1 0 108284 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1177
timestamp 1636968456
transform 1 0 109388 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1189
timestamp 1636968456
transform 1 0 110492 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1201
timestamp 1636968456
transform 1 0 111596 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_145_1213
timestamp 1
transform 1 0 112700 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_145_1217
timestamp 1
transform 1 0 113068 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1219
timestamp 1636968456
transform 1 0 113252 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1231
timestamp 1636968456
transform 1 0 114356 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1243
timestamp 1636968456
transform 1 0 115460 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1255
timestamp 1636968456
transform 1 0 116564 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_1267
timestamp 1
transform 1 0 117668 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_1273
timestamp 1
transform 1 0 118220 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_145_1275
timestamp 1
transform 1 0 118404 0 -1 81600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_3
timestamp 1636968456
transform 1 0 1380 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_15
timestamp 1636968456
transform 1 0 2484 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 1
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636968456
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_41
timestamp 1636968456
transform 1 0 4876 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_53
timestamp 1636968456
transform 1 0 5980 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_65
timestamp 1
transform 1 0 7084 0 1 81600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1165
timestamp 1636968456
transform 1 0 108284 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1177
timestamp 1636968456
transform 1 0 109388 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_1189
timestamp 1
transform 1 0 110492 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1191
timestamp 1636968456
transform 1 0 110676 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1203
timestamp 1636968456
transform 1 0 111780 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1215
timestamp 1636968456
transform 1 0 112884 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1227
timestamp 1636968456
transform 1 0 113988 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_1239
timestamp 1
transform 1 0 115092 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_1245
timestamp 1
transform 1 0 115644 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1247
timestamp 1636968456
transform 1 0 115828 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1259
timestamp 1636968456
transform 1 0 116932 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_1271
timestamp 1
transform 1 0 118036 0 1 81600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_147_3
timestamp 1636968456
transform 1 0 1380 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_15
timestamp 1636968456
transform 1 0 2484 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_27
timestamp 1636968456
transform 1 0 3588 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_39
timestamp 1636968456
transform 1 0 4692 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_147_51
timestamp 1
transform 1 0 5796 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_147_55
timestamp 1
transform 1 0 6164 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_57
timestamp 1636968456
transform 1 0 6348 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_147_69
timestamp 1
transform 1 0 7452 0 -1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1165
timestamp 1636968456
transform 1 0 108284 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1177
timestamp 1636968456
transform 1 0 109388 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1189
timestamp 1636968456
transform 1 0 110492 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1201
timestamp 1636968456
transform 1 0 111596 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_147_1213
timestamp 1
transform 1 0 112700 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_147_1217
timestamp 1
transform 1 0 113068 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1219
timestamp 1636968456
transform 1 0 113252 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1231
timestamp 1636968456
transform 1 0 114356 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1243
timestamp 1636968456
transform 1 0 115460 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1255
timestamp 1636968456
transform 1 0 116564 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_1267
timestamp 1
transform 1 0 117668 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_1273
timestamp 1
transform 1 0 118220 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_147_1275
timestamp 1
transform 1 0 118404 0 -1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636968456
transform 1 0 1380 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636968456
transform 1 0 2484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 1
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636968456
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_41
timestamp 1636968456
transform 1 0 4876 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_53
timestamp 1636968456
transform 1 0 5980 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_65
timestamp 1
transform 1 0 7084 0 1 82688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1165
timestamp 1636968456
transform 1 0 108284 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1177
timestamp 1636968456
transform 1 0 109388 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_1189
timestamp 1
transform 1 0 110492 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1191
timestamp 1636968456
transform 1 0 110676 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1203
timestamp 1636968456
transform 1 0 111780 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1215
timestamp 1636968456
transform 1 0 112884 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1227
timestamp 1636968456
transform 1 0 113988 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_1239
timestamp 1
transform 1 0 115092 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_1245
timestamp 1
transform 1 0 115644 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1247
timestamp 1636968456
transform 1 0 115828 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1259
timestamp 1636968456
transform 1 0 116932 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_1271
timestamp 1
transform 1 0 118036 0 1 82688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_149_3
timestamp 1636968456
transform 1 0 1380 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_15
timestamp 1636968456
transform 1 0 2484 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_27
timestamp 1636968456
transform 1 0 3588 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_39
timestamp 1636968456
transform 1 0 4692 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_149_51
timestamp 1
transform 1 0 5796 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_55
timestamp 1
transform 1 0 6164 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_57
timestamp 1636968456
transform 1 0 6348 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_149_69
timestamp 1
transform 1 0 7452 0 -1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1165
timestamp 1636968456
transform 1 0 108284 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1177
timestamp 1636968456
transform 1 0 109388 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1189
timestamp 1636968456
transform 1 0 110492 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1201
timestamp 1636968456
transform 1 0 111596 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_149_1213
timestamp 1
transform 1 0 112700 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_1217
timestamp 1
transform 1 0 113068 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1219
timestamp 1636968456
transform 1 0 113252 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1231
timestamp 1636968456
transform 1 0 114356 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1243
timestamp 1636968456
transform 1 0 115460 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1255
timestamp 1636968456
transform 1 0 116564 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_1267
timestamp 1
transform 1 0 117668 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_1273
timestamp 1
transform 1 0 118220 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_149_1275
timestamp 1
transform 1 0 118404 0 -1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_150_3
timestamp 1636968456
transform 1 0 1380 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_15
timestamp 1636968456
transform 1 0 2484 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 1
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636968456
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_41
timestamp 1636968456
transform 1 0 4876 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_53
timestamp 1636968456
transform 1 0 5980 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_65
timestamp 1
transform 1 0 7084 0 1 83776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1165
timestamp 1636968456
transform 1 0 108284 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1177
timestamp 1636968456
transform 1 0 109388 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_1189
timestamp 1
transform 1 0 110492 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1191
timestamp 1636968456
transform 1 0 110676 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1203
timestamp 1636968456
transform 1 0 111780 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1215
timestamp 1636968456
transform 1 0 112884 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1227
timestamp 1636968456
transform 1 0 113988 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_1239
timestamp 1
transform 1 0 115092 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_1245
timestamp 1
transform 1 0 115644 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1247
timestamp 1636968456
transform 1 0 115828 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1259
timestamp 1636968456
transform 1 0 116932 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_1271
timestamp 1
transform 1 0 118036 0 1 83776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_151_3
timestamp 1636968456
transform 1 0 1380 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_15
timestamp 1636968456
transform 1 0 2484 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_27
timestamp 1636968456
transform 1 0 3588 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_39
timestamp 1636968456
transform 1 0 4692 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_51
timestamp 1
transform 1 0 5796 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_55
timestamp 1
transform 1 0 6164 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_57
timestamp 1636968456
transform 1 0 6348 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_151_69
timestamp 1
transform 1 0 7452 0 -1 84864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1165
timestamp 1636968456
transform 1 0 108284 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1177
timestamp 1636968456
transform 1 0 109388 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1189
timestamp 1636968456
transform 1 0 110492 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1201
timestamp 1636968456
transform 1 0 111596 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_1213
timestamp 1
transform 1 0 112700 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_1217
timestamp 1
transform 1 0 113068 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1219
timestamp 1636968456
transform 1 0 113252 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1231
timestamp 1636968456
transform 1 0 114356 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1243
timestamp 1636968456
transform 1 0 115460 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1255
timestamp 1636968456
transform 1 0 116564 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_1267
timestamp 1
transform 1 0 117668 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_1273
timestamp 1
transform 1 0 118220 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_151_1275
timestamp 1
transform 1 0 118404 0 -1 84864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_152_3
timestamp 1636968456
transform 1 0 1380 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_15
timestamp 1636968456
transform 1 0 2484 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 1
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_29
timestamp 1636968456
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_41
timestamp 1636968456
transform 1 0 4876 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_53
timestamp 1636968456
transform 1 0 5980 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_65
timestamp 1
transform 1 0 7084 0 1 84864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1165
timestamp 1636968456
transform 1 0 108284 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1177
timestamp 1636968456
transform 1 0 109388 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_1189
timestamp 1
transform 1 0 110492 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1191
timestamp 1636968456
transform 1 0 110676 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1203
timestamp 1636968456
transform 1 0 111780 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1215
timestamp 1636968456
transform 1 0 112884 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1227
timestamp 1636968456
transform 1 0 113988 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_1239
timestamp 1
transform 1 0 115092 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_1245
timestamp 1
transform 1 0 115644 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1247
timestamp 1636968456
transform 1 0 115828 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1259
timestamp 1636968456
transform 1 0 116932 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_1271
timestamp 1
transform 1 0 118036 0 1 84864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_153_3
timestamp 1636968456
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_15
timestamp 1636968456
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_27
timestamp 1636968456
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_39
timestamp 1636968456
transform 1 0 4692 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_51
timestamp 1
transform 1 0 5796 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_55
timestamp 1
transform 1 0 6164 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_57
timestamp 1636968456
transform 1 0 6348 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_153_69
timestamp 1
transform 1 0 7452 0 -1 85952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1165
timestamp 1636968456
transform 1 0 108284 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1177
timestamp 1636968456
transform 1 0 109388 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1189
timestamp 1636968456
transform 1 0 110492 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1201
timestamp 1636968456
transform 1 0 111596 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_1213
timestamp 1
transform 1 0 112700 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_1217
timestamp 1
transform 1 0 113068 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1219
timestamp 1636968456
transform 1 0 113252 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1231
timestamp 1636968456
transform 1 0 114356 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1243
timestamp 1636968456
transform 1 0 115460 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1255
timestamp 1636968456
transform 1 0 116564 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_1267
timestamp 1
transform 1 0 117668 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_1273
timestamp 1
transform 1 0 118220 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_153_1275
timestamp 1
transform 1 0 118404 0 -1 85952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_154_3
timestamp 1636968456
transform 1 0 1380 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_15
timestamp 1636968456
transform 1 0 2484 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_27
timestamp 1
transform 1 0 3588 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_29
timestamp 1636968456
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_41
timestamp 1636968456
transform 1 0 4876 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_53
timestamp 1636968456
transform 1 0 5980 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_65
timestamp 1
transform 1 0 7084 0 1 85952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1165
timestamp 1636968456
transform 1 0 108284 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1177
timestamp 1636968456
transform 1 0 109388 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_1189
timestamp 1
transform 1 0 110492 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1191
timestamp 1636968456
transform 1 0 110676 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1203
timestamp 1636968456
transform 1 0 111780 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1215
timestamp 1636968456
transform 1 0 112884 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1227
timestamp 1636968456
transform 1 0 113988 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_1239
timestamp 1
transform 1 0 115092 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_1245
timestamp 1
transform 1 0 115644 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1247
timestamp 1636968456
transform 1 0 115828 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1259
timestamp 1636968456
transform 1 0 116932 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_1271
timestamp 1
transform 1 0 118036 0 1 85952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_155_3
timestamp 1636968456
transform 1 0 1380 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_15
timestamp 1636968456
transform 1 0 2484 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_27
timestamp 1636968456
transform 1 0 3588 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_39
timestamp 1636968456
transform 1 0 4692 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_155_51
timestamp 1
transform 1 0 5796 0 -1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_155_55
timestamp 1
transform 1 0 6164 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_57
timestamp 1636968456
transform 1 0 6348 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_155_69
timestamp 1
transform 1 0 7452 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1168
timestamp 1636968456
transform 1 0 108560 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1180
timestamp 1636968456
transform 1 0 109664 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1192
timestamp 1636968456
transform 1 0 110768 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1204
timestamp 1636968456
transform 1 0 111872 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_155_1216
timestamp 1
transform 1 0 112976 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1219
timestamp 1636968456
transform 1 0 113252 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1231
timestamp 1636968456
transform 1 0 114356 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1243
timestamp 1636968456
transform 1 0 115460 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1255
timestamp 1636968456
transform 1 0 116564 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_1267
timestamp 1
transform 1 0 117668 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_1273
timestamp 1
transform 1 0 118220 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_155_1275
timestamp 1
transform 1 0 118404 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_156_3
timestamp 1636968456
transform 1 0 1380 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_15
timestamp 1636968456
transform 1 0 2484 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_27
timestamp 1
transform 1 0 3588 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_29
timestamp 1636968456
transform 1 0 3772 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_41
timestamp 1636968456
transform 1 0 4876 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_53
timestamp 1636968456
transform 1 0 5980 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_65
timestamp 1
transform 1 0 7084 0 1 87040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1165
timestamp 1636968456
transform 1 0 108284 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1177
timestamp 1636968456
transform 1 0 109388 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_1189
timestamp 1
transform 1 0 110492 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1191
timestamp 1636968456
transform 1 0 110676 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1203
timestamp 1636968456
transform 1 0 111780 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1215
timestamp 1636968456
transform 1 0 112884 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1227
timestamp 1636968456
transform 1 0 113988 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_1239
timestamp 1
transform 1 0 115092 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_1245
timestamp 1
transform 1 0 115644 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1247
timestamp 1636968456
transform 1 0 115828 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1259
timestamp 1636968456
transform 1 0 116932 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_1271
timestamp 1
transform 1 0 118036 0 1 87040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_157_3
timestamp 1636968456
transform 1 0 1380 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_15
timestamp 1636968456
transform 1 0 2484 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_27
timestamp 1636968456
transform 1 0 3588 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_39
timestamp 1636968456
transform 1 0 4692 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_157_51
timestamp 1
transform 1 0 5796 0 -1 88128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_157_55
timestamp 1
transform 1 0 6164 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_57
timestamp 1636968456
transform 1 0 6348 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_157_69
timestamp 1
transform 1 0 7452 0 -1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1165
timestamp 1636968456
transform 1 0 108284 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1177
timestamp 1636968456
transform 1 0 109388 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1189
timestamp 1636968456
transform 1 0 110492 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1201
timestamp 1636968456
transform 1 0 111596 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_157_1213
timestamp 1
transform 1 0 112700 0 -1 88128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_157_1217
timestamp 1
transform 1 0 113068 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1219
timestamp 1636968456
transform 1 0 113252 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1231
timestamp 1636968456
transform 1 0 114356 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1243
timestamp 1636968456
transform 1 0 115460 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1255
timestamp 1636968456
transform 1 0 116564 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_1267
timestamp 1
transform 1 0 117668 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_1273
timestamp 1
transform 1 0 118220 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_157_1275
timestamp 1
transform 1 0 118404 0 -1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_158_3
timestamp 1636968456
transform 1 0 1380 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_15
timestamp 1636968456
transform 1 0 2484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_27
timestamp 1
transform 1 0 3588 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_29
timestamp 1636968456
transform 1 0 3772 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_41
timestamp 1636968456
transform 1 0 4876 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_53
timestamp 1636968456
transform 1 0 5980 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_65
timestamp 1
transform 1 0 7084 0 1 88128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1165
timestamp 1636968456
transform 1 0 108284 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1177
timestamp 1636968456
transform 1 0 109388 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_1189
timestamp 1
transform 1 0 110492 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1191
timestamp 1636968456
transform 1 0 110676 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1203
timestamp 1636968456
transform 1 0 111780 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1215
timestamp 1636968456
transform 1 0 112884 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1227
timestamp 1636968456
transform 1 0 113988 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_1239
timestamp 1
transform 1 0 115092 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_1245
timestamp 1
transform 1 0 115644 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1247
timestamp 1636968456
transform 1 0 115828 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1259
timestamp 1636968456
transform 1 0 116932 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_1271
timestamp 1
transform 1 0 118036 0 1 88128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_159_3
timestamp 1636968456
transform 1 0 1380 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_15
timestamp 1636968456
transform 1 0 2484 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_27
timestamp 1636968456
transform 1 0 3588 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_39
timestamp 1636968456
transform 1 0 4692 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_159_51
timestamp 1
transform 1 0 5796 0 -1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_159_55
timestamp 1
transform 1 0 6164 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_57
timestamp 1636968456
transform 1 0 6348 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_159_69
timestamp 1
transform 1 0 7452 0 -1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1165
timestamp 1636968456
transform 1 0 108284 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1177
timestamp 1636968456
transform 1 0 109388 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1189
timestamp 1636968456
transform 1 0 110492 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1201
timestamp 1636968456
transform 1 0 111596 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_159_1213
timestamp 1
transform 1 0 112700 0 -1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_159_1217
timestamp 1
transform 1 0 113068 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1219
timestamp 1636968456
transform 1 0 113252 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1231
timestamp 1636968456
transform 1 0 114356 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1243
timestamp 1636968456
transform 1 0 115460 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1255
timestamp 1636968456
transform 1 0 116564 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_1267
timestamp 1
transform 1 0 117668 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_1273
timestamp 1
transform 1 0 118220 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_159_1275
timestamp 1
transform 1 0 118404 0 -1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_160_3
timestamp 1636968456
transform 1 0 1380 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_15
timestamp 1636968456
transform 1 0 2484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_27
timestamp 1
transform 1 0 3588 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_29
timestamp 1636968456
transform 1 0 3772 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_41
timestamp 1636968456
transform 1 0 4876 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_53
timestamp 1636968456
transform 1 0 5980 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_65
timestamp 1
transform 1 0 7084 0 1 89216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1165
timestamp 1636968456
transform 1 0 108284 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1177
timestamp 1636968456
transform 1 0 109388 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_1189
timestamp 1
transform 1 0 110492 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1191
timestamp 1636968456
transform 1 0 110676 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1203
timestamp 1636968456
transform 1 0 111780 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1215
timestamp 1636968456
transform 1 0 112884 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1227
timestamp 1636968456
transform 1 0 113988 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_1239
timestamp 1
transform 1 0 115092 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_1245
timestamp 1
transform 1 0 115644 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1247
timestamp 1636968456
transform 1 0 115828 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1259
timestamp 1636968456
transform 1 0 116932 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_1271
timestamp 1
transform 1 0 118036 0 1 89216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_161_3
timestamp 1636968456
transform 1 0 1380 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_15
timestamp 1636968456
transform 1 0 2484 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_27
timestamp 1636968456
transform 1 0 3588 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_39
timestamp 1636968456
transform 1 0 4692 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_161_51
timestamp 1
transform 1 0 5796 0 -1 90304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_161_55
timestamp 1
transform 1 0 6164 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_57
timestamp 1636968456
transform 1 0 6348 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_161_69
timestamp 1
transform 1 0 7452 0 -1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1165
timestamp 1636968456
transform 1 0 108284 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1177
timestamp 1636968456
transform 1 0 109388 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1189
timestamp 1636968456
transform 1 0 110492 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1201
timestamp 1636968456
transform 1 0 111596 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_161_1213
timestamp 1
transform 1 0 112700 0 -1 90304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_161_1217
timestamp 1
transform 1 0 113068 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1219
timestamp 1636968456
transform 1 0 113252 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1231
timestamp 1636968456
transform 1 0 114356 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1243
timestamp 1636968456
transform 1 0 115460 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1255
timestamp 1636968456
transform 1 0 116564 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_1267
timestamp 1
transform 1 0 117668 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_1273
timestamp 1
transform 1 0 118220 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_161_1275
timestamp 1
transform 1 0 118404 0 -1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_162_3
timestamp 1636968456
transform 1 0 1380 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_15
timestamp 1636968456
transform 1 0 2484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_27
timestamp 1
transform 1 0 3588 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_29
timestamp 1636968456
transform 1 0 3772 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_41
timestamp 1636968456
transform 1 0 4876 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_53
timestamp 1636968456
transform 1 0 5980 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_65
timestamp 1
transform 1 0 7084 0 1 90304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1165
timestamp 1636968456
transform 1 0 108284 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1177
timestamp 1636968456
transform 1 0 109388 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_1189
timestamp 1
transform 1 0 110492 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1191
timestamp 1636968456
transform 1 0 110676 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1203
timestamp 1636968456
transform 1 0 111780 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1215
timestamp 1636968456
transform 1 0 112884 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1227
timestamp 1636968456
transform 1 0 113988 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_1239
timestamp 1
transform 1 0 115092 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_1245
timestamp 1
transform 1 0 115644 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1247
timestamp 1636968456
transform 1 0 115828 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1259
timestamp 1636968456
transform 1 0 116932 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_1271
timestamp 1
transform 1 0 118036 0 1 90304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_163_3
timestamp 1636968456
transform 1 0 1380 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_15
timestamp 1636968456
transform 1 0 2484 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_27
timestamp 1636968456
transform 1 0 3588 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_39
timestamp 1636968456
transform 1 0 4692 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_163_51
timestamp 1
transform 1 0 5796 0 -1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_163_55
timestamp 1
transform 1 0 6164 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_57
timestamp 1636968456
transform 1 0 6348 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_163_69
timestamp 1
transform 1 0 7452 0 -1 91392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1165
timestamp 1636968456
transform 1 0 108284 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1177
timestamp 1636968456
transform 1 0 109388 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1189
timestamp 1636968456
transform 1 0 110492 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1201
timestamp 1636968456
transform 1 0 111596 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_163_1213
timestamp 1
transform 1 0 112700 0 -1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_163_1217
timestamp 1
transform 1 0 113068 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1219
timestamp 1636968456
transform 1 0 113252 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1231
timestamp 1636968456
transform 1 0 114356 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1243
timestamp 1636968456
transform 1 0 115460 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1255
timestamp 1636968456
transform 1 0 116564 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_1267
timestamp 1
transform 1 0 117668 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_1273
timestamp 1
transform 1 0 118220 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_163_1275
timestamp 1
transform 1 0 118404 0 -1 91392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_164_3
timestamp 1636968456
transform 1 0 1380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_15
timestamp 1636968456
transform 1 0 2484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_27
timestamp 1
transform 1 0 3588 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_29
timestamp 1636968456
transform 1 0 3772 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_41
timestamp 1636968456
transform 1 0 4876 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_53
timestamp 1636968456
transform 1 0 5980 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_65
timestamp 1
transform 1 0 7084 0 1 91392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1165
timestamp 1636968456
transform 1 0 108284 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1177
timestamp 1636968456
transform 1 0 109388 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_1189
timestamp 1
transform 1 0 110492 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1191
timestamp 1636968456
transform 1 0 110676 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1203
timestamp 1636968456
transform 1 0 111780 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1215
timestamp 1636968456
transform 1 0 112884 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1227
timestamp 1636968456
transform 1 0 113988 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_1239
timestamp 1
transform 1 0 115092 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_1245
timestamp 1
transform 1 0 115644 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1247
timestamp 1636968456
transform 1 0 115828 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1259
timestamp 1636968456
transform 1 0 116932 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_1271
timestamp 1
transform 1 0 118036 0 1 91392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_165_3
timestamp 1636968456
transform 1 0 1380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_15
timestamp 1636968456
transform 1 0 2484 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_165_27
timestamp 1
transform 1 0 3588 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_29
timestamp 1636968456
transform 1 0 3772 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_41
timestamp 1636968456
transform 1 0 4876 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_53
timestamp 1
transform 1 0 5980 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_57
timestamp 1636968456
transform 1 0 6348 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_69
timestamp 1636968456
transform 1 0 7452 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_81
timestamp 1
transform 1 0 8556 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_85
timestamp 1636968456
transform 1 0 8924 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_97
timestamp 1636968456
transform 1 0 10028 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_109
timestamp 1
transform 1 0 11132 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_113
timestamp 1636968456
transform 1 0 11500 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_125
timestamp 1636968456
transform 1 0 12604 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_137
timestamp 1
transform 1 0 13708 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_141
timestamp 1636968456
transform 1 0 14076 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_153
timestamp 1636968456
transform 1 0 15180 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_165
timestamp 1
transform 1 0 16284 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_169
timestamp 1636968456
transform 1 0 16652 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_181
timestamp 1636968456
transform 1 0 17756 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_193
timestamp 1
transform 1 0 18860 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_197
timestamp 1636968456
transform 1 0 19228 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_209
timestamp 1636968456
transform 1 0 20332 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_221
timestamp 1
transform 1 0 21436 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_225
timestamp 1636968456
transform 1 0 21804 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_237
timestamp 1636968456
transform 1 0 22908 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_249
timestamp 1
transform 1 0 24012 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_253
timestamp 1636968456
transform 1 0 24380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_265
timestamp 1636968456
transform 1 0 25484 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_277
timestamp 1
transform 1 0 26588 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_281
timestamp 1636968456
transform 1 0 26956 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_293
timestamp 1636968456
transform 1 0 28060 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_305
timestamp 1
transform 1 0 29164 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_309
timestamp 1636968456
transform 1 0 29532 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_321
timestamp 1636968456
transform 1 0 30636 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_333
timestamp 1
transform 1 0 31740 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_337
timestamp 1636968456
transform 1 0 32108 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_349
timestamp 1636968456
transform 1 0 33212 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_361
timestamp 1
transform 1 0 34316 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_365
timestamp 1636968456
transform 1 0 34684 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_377
timestamp 1636968456
transform 1 0 35788 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_389
timestamp 1
transform 1 0 36892 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_393
timestamp 1636968456
transform 1 0 37260 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_405
timestamp 1636968456
transform 1 0 38364 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_417
timestamp 1
transform 1 0 39468 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_421
timestamp 1636968456
transform 1 0 39836 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_433
timestamp 1636968456
transform 1 0 40940 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_445
timestamp 1
transform 1 0 42044 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_449
timestamp 1636968456
transform 1 0 42412 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_461
timestamp 1636968456
transform 1 0 43516 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_473
timestamp 1
transform 1 0 44620 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_165_477
timestamp 1
transform 1 0 44988 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_165_503
timestamp 1
transform 1 0 47380 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_165_505
timestamp 1
transform 1 0 47564 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_165_528
timestamp 1
transform 1 0 49680 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_165_533
timestamp 1
transform 1 0 50140 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_552
timestamp 1
transform 1 0 51888 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_165_561
timestamp 1
transform 1 0 52716 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_165_565
timestamp 1
transform 1 0 53084 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_165_584
timestamp 1
transform 1 0 54832 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_165_589
timestamp 1
transform 1 0 55292 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_165_597
timestamp 1
transform 1 0 56028 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_617
timestamp 1
transform 1 0 57868 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_165_625
timestamp 1
transform 1 0 58604 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_165_645
timestamp 1
transform 1 0 60444 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_664
timestamp 1
transform 1 0 62192 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_165_673
timestamp 1
transform 1 0 63020 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_165_699
timestamp 1
transform 1 0 65412 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_701
timestamp 1636968456
transform 1 0 65596 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_713
timestamp 1636968456
transform 1 0 66700 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_725
timestamp 1
transform 1 0 67804 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_165_729
timestamp 1
transform 1 0 68172 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_165_746
timestamp 1
transform 1 0 69736 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_757
timestamp 1
transform 1 0 70748 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_165_782
timestamp 1
transform 1 0 73048 0 -1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_165_803
timestamp 1
transform 1 0 74980 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_165_811
timestamp 1
transform 1 0 75716 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_813
timestamp 1636968456
transform 1 0 75900 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_825
timestamp 1
transform 1 0 77004 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_165_829
timestamp 1
transform 1 0 77372 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_165_836
timestamp 1
transform 1 0 78016 0 -1 92480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_165_841
timestamp 1636968456
transform 1 0 78476 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_853
timestamp 1636968456
transform 1 0 79580 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_865
timestamp 1
transform 1 0 80684 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_869
timestamp 1636968456
transform 1 0 81052 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_881
timestamp 1636968456
transform 1 0 82156 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_893
timestamp 1
transform 1 0 83260 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_897
timestamp 1636968456
transform 1 0 83628 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_909
timestamp 1636968456
transform 1 0 84732 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_921
timestamp 1
transform 1 0 85836 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_925
timestamp 1636968456
transform 1 0 86204 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_937
timestamp 1636968456
transform 1 0 87308 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_949
timestamp 1
transform 1 0 88412 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_165_953
timestamp 1
transform 1 0 88780 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_959
timestamp 1
transform 1 0 89332 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_962
timestamp 1636968456
transform 1 0 89608 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_974
timestamp 1
transform 1 0 90712 0 -1 92480
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_165_981
timestamp 1636968456
transform 1 0 91356 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_993
timestamp 1636968456
transform 1 0 92460 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1005
timestamp 1
transform 1 0 93564 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1009
timestamp 1636968456
transform 1 0 93932 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1021
timestamp 1636968456
transform 1 0 95036 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1033
timestamp 1
transform 1 0 96140 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1037
timestamp 1636968456
transform 1 0 96508 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1049
timestamp 1636968456
transform 1 0 97612 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1061
timestamp 1
transform 1 0 98716 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_165_1065
timestamp 1
transform 1 0 99084 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1073
timestamp 1
transform 1 0 99820 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1078
timestamp 1636968456
transform 1 0 100280 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_165_1090
timestamp 1
transform 1 0 101384 0 -1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1093
timestamp 1636968456
transform 1 0 101660 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1105
timestamp 1636968456
transform 1 0 102764 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1117
timestamp 1
transform 1 0 103868 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1121
timestamp 1636968456
transform 1 0 104236 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1133
timestamp 1636968456
transform 1 0 105340 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1145
timestamp 1
transform 1 0 106444 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1149
timestamp 1636968456
transform 1 0 106812 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1161
timestamp 1636968456
transform 1 0 107916 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1173
timestamp 1
transform 1 0 109020 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1177
timestamp 1636968456
transform 1 0 109388 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1189
timestamp 1636968456
transform 1 0 110492 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1201
timestamp 1
transform 1 0 111596 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1205
timestamp 1636968456
transform 1 0 111964 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1217
timestamp 1636968456
transform 1 0 113068 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1229
timestamp 1
transform 1 0 114172 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1233
timestamp 1636968456
transform 1 0 114540 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1245
timestamp 1636968456
transform 1 0 115644 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_165_1257
timestamp 1
transform 1 0 116748 0 -1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1261
timestamp 1636968456
transform 1 0 117116 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_1273
timestamp 1
transform 1 0 118220 0 -1 92480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_166_3
timestamp 1636968456
transform 1 0 1380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_15
timestamp 1636968456
transform 1 0 2484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_27
timestamp 1
transform 1 0 3588 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_29
timestamp 1636968456
transform 1 0 3772 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_41
timestamp 1636968456
transform 1 0 4876 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_53
timestamp 1636968456
transform 1 0 5980 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_65
timestamp 1636968456
transform 1 0 7084 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_77
timestamp 1
transform 1 0 8188 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_83
timestamp 1
transform 1 0 8740 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_85
timestamp 1636968456
transform 1 0 8924 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_97
timestamp 1636968456
transform 1 0 10028 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_109
timestamp 1636968456
transform 1 0 11132 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_121
timestamp 1636968456
transform 1 0 12236 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_133
timestamp 1
transform 1 0 13340 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_139
timestamp 1
transform 1 0 13892 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_141
timestamp 1636968456
transform 1 0 14076 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_153
timestamp 1636968456
transform 1 0 15180 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_165
timestamp 1636968456
transform 1 0 16284 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_177
timestamp 1636968456
transform 1 0 17388 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_189
timestamp 1
transform 1 0 18492 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_195
timestamp 1
transform 1 0 19044 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_197
timestamp 1636968456
transform 1 0 19228 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_209
timestamp 1636968456
transform 1 0 20332 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_221
timestamp 1636968456
transform 1 0 21436 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_233
timestamp 1636968456
transform 1 0 22540 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_245
timestamp 1
transform 1 0 23644 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_251
timestamp 1
transform 1 0 24196 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_253
timestamp 1636968456
transform 1 0 24380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_265
timestamp 1636968456
transform 1 0 25484 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_277
timestamp 1636968456
transform 1 0 26588 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_289
timestamp 1636968456
transform 1 0 27692 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_301
timestamp 1
transform 1 0 28796 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_307
timestamp 1
transform 1 0 29348 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_309
timestamp 1636968456
transform 1 0 29532 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_321
timestamp 1636968456
transform 1 0 30636 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_333
timestamp 1636968456
transform 1 0 31740 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_345
timestamp 1636968456
transform 1 0 32844 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_357
timestamp 1
transform 1 0 33948 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_363
timestamp 1
transform 1 0 34500 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_365
timestamp 1636968456
transform 1 0 34684 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_377
timestamp 1636968456
transform 1 0 35788 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_389
timestamp 1636968456
transform 1 0 36892 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_401
timestamp 1636968456
transform 1 0 37996 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_413
timestamp 1
transform 1 0 39100 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_419
timestamp 1
transform 1 0 39652 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_421
timestamp 1636968456
transform 1 0 39836 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_433
timestamp 1636968456
transform 1 0 40940 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_445
timestamp 1636968456
transform 1 0 42044 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_457
timestamp 1636968456
transform 1 0 43148 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_469
timestamp 1
transform 1 0 44252 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_475
timestamp 1
transform 1 0 44804 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_166_477
timestamp 1
transform 1 0 44988 0 1 92480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_166_517
timestamp 1636968456
transform 1 0 48668 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_166_529
timestamp 1
transform 1 0 49772 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_166_533
timestamp 1
transform 1 0 50140 0 1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_166_537
timestamp 1
transform 1 0 50508 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_166_593
timestamp 1
transform 1 0 55660 0 1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_166_601
timestamp 1
transform 1 0 56396 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_166_636
timestamp 1
transform 1 0 59616 0 1 92480
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_166_645
timestamp 1636968456
transform 1 0 60444 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_166_657
timestamp 1
transform 1 0 61548 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_166_695
timestamp 1
transform 1 0 65044 0 1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_166_699
timestamp 1
transform 1 0 65412 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_166_749
timestamp 1
transform 1 0 70012 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_755
timestamp 1
transform 1 0 70564 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_791
timestamp 1636968456
transform 1 0 73876 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_803
timestamp 1
transform 1 0 74980 0 1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_166_811
timestamp 1
transform 1 0 75716 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_813
timestamp 1636968456
transform 1 0 75900 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_166_825
timestamp 1
transform 1 0 77004 0 1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_166_852
timestamp 1636968456
transform 1 0 79488 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_166_864
timestamp 1
transform 1 0 80592 0 1 92480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_166_869
timestamp 1636968456
transform 1 0 81052 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_881
timestamp 1636968456
transform 1 0 82156 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_893
timestamp 1636968456
transform 1 0 83260 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_905
timestamp 1636968456
transform 1 0 84364 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_917
timestamp 1
transform 1 0 85468 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_923
timestamp 1
transform 1 0 86020 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_925
timestamp 1636968456
transform 1 0 86204 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_937
timestamp 1636968456
transform 1 0 87308 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_949
timestamp 1636968456
transform 1 0 88412 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_961
timestamp 1636968456
transform 1 0 89516 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_973
timestamp 1
transform 1 0 90620 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_979
timestamp 1
transform 1 0 91172 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_981
timestamp 1636968456
transform 1 0 91356 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_993
timestamp 1636968456
transform 1 0 92460 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1005
timestamp 1636968456
transform 1 0 93564 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1017
timestamp 1636968456
transform 1 0 94668 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_1029
timestamp 1
transform 1 0 95772 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_1035
timestamp 1
transform 1 0 96324 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1037
timestamp 1636968456
transform 1 0 96508 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1049
timestamp 1636968456
transform 1 0 97612 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1061
timestamp 1636968456
transform 1 0 98716 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1073
timestamp 1636968456
transform 1 0 99820 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_1085
timestamp 1
transform 1 0 100924 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_1091
timestamp 1
transform 1 0 101476 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1093
timestamp 1636968456
transform 1 0 101660 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1105
timestamp 1636968456
transform 1 0 102764 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1117
timestamp 1636968456
transform 1 0 103868 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1129
timestamp 1636968456
transform 1 0 104972 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_1141
timestamp 1
transform 1 0 106076 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_1147
timestamp 1
transform 1 0 106628 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1149
timestamp 1636968456
transform 1 0 106812 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1161
timestamp 1636968456
transform 1 0 107916 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1173
timestamp 1636968456
transform 1 0 109020 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1185
timestamp 1636968456
transform 1 0 110124 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_1197
timestamp 1
transform 1 0 111228 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_1203
timestamp 1
transform 1 0 111780 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1205
timestamp 1636968456
transform 1 0 111964 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1217
timestamp 1636968456
transform 1 0 113068 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1229
timestamp 1636968456
transform 1 0 114172 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1241
timestamp 1636968456
transform 1 0 115276 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_1253
timestamp 1
transform 1 0 116380 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_1259
timestamp 1
transform 1 0 116932 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1261
timestamp 1636968456
transform 1 0 117116 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_166_1273
timestamp 1
transform 1 0 118220 0 1 92480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_167_3
timestamp 1636968456
transform 1 0 1380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_15
timestamp 1636968456
transform 1 0 2484 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_27
timestamp 1636968456
transform 1 0 3588 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_39
timestamp 1636968456
transform 1 0 4692 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_51
timestamp 1
transform 1 0 5796 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_55
timestamp 1
transform 1 0 6164 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_57
timestamp 1636968456
transform 1 0 6348 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_69
timestamp 1636968456
transform 1 0 7452 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_81
timestamp 1636968456
transform 1 0 8556 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_93
timestamp 1636968456
transform 1 0 9660 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_105
timestamp 1
transform 1 0 10764 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_111
timestamp 1
transform 1 0 11316 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_113
timestamp 1636968456
transform 1 0 11500 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_125
timestamp 1636968456
transform 1 0 12604 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_137
timestamp 1636968456
transform 1 0 13708 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_149
timestamp 1636968456
transform 1 0 14812 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_161
timestamp 1
transform 1 0 15916 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_167
timestamp 1
transform 1 0 16468 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_169
timestamp 1636968456
transform 1 0 16652 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_181
timestamp 1636968456
transform 1 0 17756 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_193
timestamp 1636968456
transform 1 0 18860 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_205
timestamp 1636968456
transform 1 0 19964 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_217
timestamp 1
transform 1 0 21068 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_223
timestamp 1
transform 1 0 21620 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_225
timestamp 1636968456
transform 1 0 21804 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_237
timestamp 1636968456
transform 1 0 22908 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_249
timestamp 1636968456
transform 1 0 24012 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_261
timestamp 1636968456
transform 1 0 25116 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_273
timestamp 1
transform 1 0 26220 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_279
timestamp 1
transform 1 0 26772 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_281
timestamp 1636968456
transform 1 0 26956 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_293
timestamp 1636968456
transform 1 0 28060 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_305
timestamp 1636968456
transform 1 0 29164 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_317
timestamp 1636968456
transform 1 0 30268 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_329
timestamp 1
transform 1 0 31372 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_335
timestamp 1
transform 1 0 31924 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_337
timestamp 1636968456
transform 1 0 32108 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_349
timestamp 1636968456
transform 1 0 33212 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_361
timestamp 1636968456
transform 1 0 34316 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_373
timestamp 1636968456
transform 1 0 35420 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_385
timestamp 1
transform 1 0 36524 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_391
timestamp 1
transform 1 0 37076 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_393
timestamp 1636968456
transform 1 0 37260 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_405
timestamp 1636968456
transform 1 0 38364 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_417
timestamp 1636968456
transform 1 0 39468 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_429
timestamp 1636968456
transform 1 0 40572 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_441
timestamp 1
transform 1 0 41676 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_447
timestamp 1
transform 1 0 42228 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_449
timestamp 1636968456
transform 1 0 42412 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_461
timestamp 1636968456
transform 1 0 43516 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_473
timestamp 1
transform 1 0 44620 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_167_492
timestamp 1
transform 1 0 46368 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_496
timestamp 1
transform 1 0 46736 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_167_501
timestamp 1
transform 1 0 47196 0 -1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_167_505
timestamp 1636968456
transform 1 0 47564 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_517
timestamp 1
transform 1 0 48668 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_521
timestamp 1
transform 1 0 49036 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_542
timestamp 1636968456
transform 1 0 50968 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_554
timestamp 1
transform 1 0 52072 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_167_561
timestamp 1
transform 1 0 52716 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_167_569
timestamp 1
transform 1 0 53452 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_167_581
timestamp 1
transform 1 0 54556 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_167_604
timestamp 1
transform 1 0 56672 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_167_617
timestamp 1
transform 1 0 57868 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_623
timestamp 1
transform 1 0 58420 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_167_673
timestamp 1
transform 1 0 63020 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_718
timestamp 1
transform 1 0 67160 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_167_726
timestamp 1
transform 1 0 67896 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_167_747
timestamp 1
transform 1 0 69828 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_167_783
timestamp 1
transform 1 0 73140 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_167_789
timestamp 1
transform 1 0 73692 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_808
timestamp 1636968456
transform 1 0 75440 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_820
timestamp 1636968456
transform 1 0 76544 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_832
timestamp 1
transform 1 0 77648 0 -1 93568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_167_841
timestamp 1636968456
transform 1 0 78476 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_853
timestamp 1636968456
transform 1 0 79580 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_865
timestamp 1636968456
transform 1 0 80684 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_877
timestamp 1636968456
transform 1 0 81788 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_889
timestamp 1
transform 1 0 82892 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_895
timestamp 1
transform 1 0 83444 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_897
timestamp 1636968456
transform 1 0 83628 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_909
timestamp 1636968456
transform 1 0 84732 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_921
timestamp 1636968456
transform 1 0 85836 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_933
timestamp 1636968456
transform 1 0 86940 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_945
timestamp 1
transform 1 0 88044 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_951
timestamp 1
transform 1 0 88596 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_953
timestamp 1636968456
transform 1 0 88780 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_965
timestamp 1636968456
transform 1 0 89884 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_977
timestamp 1636968456
transform 1 0 90988 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_989
timestamp 1636968456
transform 1 0 92092 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_1001
timestamp 1
transform 1 0 93196 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_1007
timestamp 1
transform 1 0 93748 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1009
timestamp 1636968456
transform 1 0 93932 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1021
timestamp 1636968456
transform 1 0 95036 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1033
timestamp 1636968456
transform 1 0 96140 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1045
timestamp 1636968456
transform 1 0 97244 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_1057
timestamp 1
transform 1 0 98348 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_1063
timestamp 1
transform 1 0 98900 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1065
timestamp 1636968456
transform 1 0 99084 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1077
timestamp 1636968456
transform 1 0 100188 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1089
timestamp 1636968456
transform 1 0 101292 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1101
timestamp 1636968456
transform 1 0 102396 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_1113
timestamp 1
transform 1 0 103500 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_1119
timestamp 1
transform 1 0 104052 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1121
timestamp 1636968456
transform 1 0 104236 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1133
timestamp 1636968456
transform 1 0 105340 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1145
timestamp 1636968456
transform 1 0 106444 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1157
timestamp 1636968456
transform 1 0 107548 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_1169
timestamp 1
transform 1 0 108652 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_1175
timestamp 1
transform 1 0 109204 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1177
timestamp 1636968456
transform 1 0 109388 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1189
timestamp 1636968456
transform 1 0 110492 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1201
timestamp 1636968456
transform 1 0 111596 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1213
timestamp 1636968456
transform 1 0 112700 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_1225
timestamp 1
transform 1 0 113804 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_1231
timestamp 1
transform 1 0 114356 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1233
timestamp 1636968456
transform 1 0 114540 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1245
timestamp 1636968456
transform 1 0 115644 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1257
timestamp 1636968456
transform 1 0 116748 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_1269
timestamp 1
transform 1 0 117852 0 -1 93568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_168_3
timestamp 1636968456
transform 1 0 1380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_15
timestamp 1636968456
transform 1 0 2484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_27
timestamp 1
transform 1 0 3588 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_29
timestamp 1636968456
transform 1 0 3772 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_41
timestamp 1636968456
transform 1 0 4876 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_53
timestamp 1636968456
transform 1 0 5980 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_65
timestamp 1636968456
transform 1 0 7084 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_77
timestamp 1
transform 1 0 8188 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_83
timestamp 1
transform 1 0 8740 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_85
timestamp 1636968456
transform 1 0 8924 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_97
timestamp 1636968456
transform 1 0 10028 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_109
timestamp 1636968456
transform 1 0 11132 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_121
timestamp 1636968456
transform 1 0 12236 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_133
timestamp 1
transform 1 0 13340 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_139
timestamp 1
transform 1 0 13892 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_141
timestamp 1636968456
transform 1 0 14076 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_153
timestamp 1636968456
transform 1 0 15180 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_165
timestamp 1636968456
transform 1 0 16284 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_177
timestamp 1636968456
transform 1 0 17388 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_189
timestamp 1
transform 1 0 18492 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_195
timestamp 1
transform 1 0 19044 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_197
timestamp 1636968456
transform 1 0 19228 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_209
timestamp 1636968456
transform 1 0 20332 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_221
timestamp 1636968456
transform 1 0 21436 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_233
timestamp 1636968456
transform 1 0 22540 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_245
timestamp 1
transform 1 0 23644 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_251
timestamp 1
transform 1 0 24196 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_253
timestamp 1636968456
transform 1 0 24380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_265
timestamp 1636968456
transform 1 0 25484 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_277
timestamp 1636968456
transform 1 0 26588 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_289
timestamp 1636968456
transform 1 0 27692 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_301
timestamp 1
transform 1 0 28796 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_307
timestamp 1
transform 1 0 29348 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_309
timestamp 1636968456
transform 1 0 29532 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_321
timestamp 1636968456
transform 1 0 30636 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_333
timestamp 1636968456
transform 1 0 31740 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_345
timestamp 1636968456
transform 1 0 32844 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_357
timestamp 1
transform 1 0 33948 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_363
timestamp 1
transform 1 0 34500 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_365
timestamp 1636968456
transform 1 0 34684 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_377
timestamp 1636968456
transform 1 0 35788 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_389
timestamp 1636968456
transform 1 0 36892 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_401
timestamp 1636968456
transform 1 0 37996 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_413
timestamp 1
transform 1 0 39100 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_419
timestamp 1
transform 1 0 39652 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_421
timestamp 1636968456
transform 1 0 39836 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_433
timestamp 1636968456
transform 1 0 40940 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_445
timestamp 1636968456
transform 1 0 42044 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_457
timestamp 1636968456
transform 1 0 43148 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_469
timestamp 1
transform 1 0 44252 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_475
timestamp 1
transform 1 0 44804 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_477
timestamp 1636968456
transform 1 0 44988 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_489
timestamp 1636968456
transform 1 0 46092 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_501
timestamp 1636968456
transform 1 0 47196 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_513
timestamp 1636968456
transform 1 0 48300 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_525
timestamp 1
transform 1 0 49404 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_531
timestamp 1
transform 1 0 49956 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_533
timestamp 1636968456
transform 1 0 50140 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_545
timestamp 1636968456
transform 1 0 51244 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_557
timestamp 1636968456
transform 1 0 52348 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_569
timestamp 1636968456
transform 1 0 53452 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_581
timestamp 1
transform 1 0 54556 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_168_585
timestamp 1
transform 1 0 54924 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_168_589
timestamp 1
transform 1 0 55292 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_168_610
timestamp 1
transform 1 0 57224 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_654
timestamp 1
transform 1 0 61272 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_168_676
timestamp 1
transform 1 0 63296 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_168_686
timestamp 1
transform 1 0 64216 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_168_699
timestamp 1
transform 1 0 65412 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_168_713
timestamp 1
transform 1 0 66700 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_168_719
timestamp 1
transform 1 0 67252 0 1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_168_727
timestamp 1
transform 1 0 67988 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_168_741
timestamp 1
transform 1 0 69276 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_168_750
timestamp 1
transform 1 0 70104 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_168_762
timestamp 1
transform 1 0 71208 0 1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_168_770
timestamp 1
transform 1 0 71944 0 1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_168_775
timestamp 1636968456
transform 1 0 72404 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_787
timestamp 1636968456
transform 1 0 73508 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_799
timestamp 1636968456
transform 1 0 74612 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_811
timestamp 1
transform 1 0 75716 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_813
timestamp 1636968456
transform 1 0 75900 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_825
timestamp 1636968456
transform 1 0 77004 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_837
timestamp 1636968456
transform 1 0 78108 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_849
timestamp 1636968456
transform 1 0 79212 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_861
timestamp 1
transform 1 0 80316 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_867
timestamp 1
transform 1 0 80868 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_869
timestamp 1636968456
transform 1 0 81052 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_881
timestamp 1636968456
transform 1 0 82156 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_893
timestamp 1636968456
transform 1 0 83260 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_905
timestamp 1636968456
transform 1 0 84364 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_917
timestamp 1
transform 1 0 85468 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_923
timestamp 1
transform 1 0 86020 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_925
timestamp 1636968456
transform 1 0 86204 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_937
timestamp 1636968456
transform 1 0 87308 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_949
timestamp 1636968456
transform 1 0 88412 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_961
timestamp 1636968456
transform 1 0 89516 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_973
timestamp 1
transform 1 0 90620 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_979
timestamp 1
transform 1 0 91172 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_981
timestamp 1636968456
transform 1 0 91356 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_993
timestamp 1636968456
transform 1 0 92460 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1005
timestamp 1636968456
transform 1 0 93564 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1017
timestamp 1636968456
transform 1 0 94668 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_1029
timestamp 1
transform 1 0 95772 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_1035
timestamp 1
transform 1 0 96324 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1037
timestamp 1636968456
transform 1 0 96508 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1049
timestamp 1636968456
transform 1 0 97612 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1061
timestamp 1636968456
transform 1 0 98716 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1073
timestamp 1636968456
transform 1 0 99820 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_1085
timestamp 1
transform 1 0 100924 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_1091
timestamp 1
transform 1 0 101476 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1093
timestamp 1636968456
transform 1 0 101660 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1105
timestamp 1636968456
transform 1 0 102764 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1117
timestamp 1636968456
transform 1 0 103868 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1129
timestamp 1636968456
transform 1 0 104972 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_1141
timestamp 1
transform 1 0 106076 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_1147
timestamp 1
transform 1 0 106628 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1149
timestamp 1636968456
transform 1 0 106812 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1161
timestamp 1636968456
transform 1 0 107916 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1173
timestamp 1636968456
transform 1 0 109020 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1185
timestamp 1636968456
transform 1 0 110124 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_1197
timestamp 1
transform 1 0 111228 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_1203
timestamp 1
transform 1 0 111780 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1205
timestamp 1636968456
transform 1 0 111964 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1217
timestamp 1636968456
transform 1 0 113068 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1229
timestamp 1636968456
transform 1 0 114172 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1241
timestamp 1636968456
transform 1 0 115276 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_1253
timestamp 1
transform 1 0 116380 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_1259
timestamp 1
transform 1 0 116932 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1261
timestamp 1636968456
transform 1 0 117116 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_168_1273
timestamp 1
transform 1 0 118220 0 1 93568
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_169_3
timestamp 1636968456
transform 1 0 1380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_15
timestamp 1636968456
transform 1 0 2484 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_27
timestamp 1636968456
transform 1 0 3588 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_39
timestamp 1636968456
transform 1 0 4692 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_51
timestamp 1
transform 1 0 5796 0 -1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_169_55
timestamp 1
transform 1 0 6164 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_57
timestamp 1636968456
transform 1 0 6348 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_69
timestamp 1636968456
transform 1 0 7452 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_81
timestamp 1636968456
transform 1 0 8556 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_93
timestamp 1636968456
transform 1 0 9660 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_105
timestamp 1
transform 1 0 10764 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_111
timestamp 1
transform 1 0 11316 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_113
timestamp 1636968456
transform 1 0 11500 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_125
timestamp 1636968456
transform 1 0 12604 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_137
timestamp 1636968456
transform 1 0 13708 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_149
timestamp 1636968456
transform 1 0 14812 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_161
timestamp 1
transform 1 0 15916 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_167
timestamp 1
transform 1 0 16468 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_169
timestamp 1636968456
transform 1 0 16652 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_181
timestamp 1636968456
transform 1 0 17756 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_193
timestamp 1636968456
transform 1 0 18860 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_205
timestamp 1636968456
transform 1 0 19964 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_217
timestamp 1
transform 1 0 21068 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_223
timestamp 1
transform 1 0 21620 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_225
timestamp 1636968456
transform 1 0 21804 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_237
timestamp 1636968456
transform 1 0 22908 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_249
timestamp 1636968456
transform 1 0 24012 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_261
timestamp 1636968456
transform 1 0 25116 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_273
timestamp 1
transform 1 0 26220 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_279
timestamp 1
transform 1 0 26772 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_281
timestamp 1636968456
transform 1 0 26956 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_293
timestamp 1636968456
transform 1 0 28060 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_305
timestamp 1636968456
transform 1 0 29164 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_317
timestamp 1636968456
transform 1 0 30268 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_329
timestamp 1
transform 1 0 31372 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_335
timestamp 1
transform 1 0 31924 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_337
timestamp 1636968456
transform 1 0 32108 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_349
timestamp 1636968456
transform 1 0 33212 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_361
timestamp 1636968456
transform 1 0 34316 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_373
timestamp 1636968456
transform 1 0 35420 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_385
timestamp 1
transform 1 0 36524 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_391
timestamp 1
transform 1 0 37076 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_393
timestamp 1636968456
transform 1 0 37260 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_405
timestamp 1636968456
transform 1 0 38364 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_417
timestamp 1636968456
transform 1 0 39468 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_429
timestamp 1636968456
transform 1 0 40572 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_441
timestamp 1
transform 1 0 41676 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_447
timestamp 1
transform 1 0 42228 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_449
timestamp 1636968456
transform 1 0 42412 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_461
timestamp 1636968456
transform 1 0 43516 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_473
timestamp 1636968456
transform 1 0 44620 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_485
timestamp 1636968456
transform 1 0 45724 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_497
timestamp 1
transform 1 0 46828 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_503
timestamp 1
transform 1 0 47380 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_505
timestamp 1636968456
transform 1 0 47564 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_517
timestamp 1636968456
transform 1 0 48668 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_529
timestamp 1636968456
transform 1 0 49772 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_541
timestamp 1636968456
transform 1 0 50876 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_553
timestamp 1
transform 1 0 51980 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_559
timestamp 1
transform 1 0 52532 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_561
timestamp 1636968456
transform 1 0 52716 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_573
timestamp 1
transform 1 0 53820 0 -1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_169_608
timestamp 1
transform 1 0 57040 0 -1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_169_617
timestamp 1
transform 1 0 57868 0 -1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_169_628
timestamp 1
transform 1 0 58880 0 -1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_169_655
timestamp 1
transform 1 0 61364 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_169_661
timestamp 1
transform 1 0 61916 0 -1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_169_669
timestamp 1
transform 1 0 62652 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_169_673
timestamp 1
transform 1 0 63020 0 -1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_169_689
timestamp 1
transform 1 0 64492 0 -1 94656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_169_700
timestamp 1636968456
transform 1 0 65504 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_712
timestamp 1636968456
transform 1 0 66608 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_724
timestamp 1
transform 1 0 67712 0 -1 94656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_169_729
timestamp 1636968456
transform 1 0 68172 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_741
timestamp 1636968456
transform 1 0 69276 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_753
timestamp 1636968456
transform 1 0 70380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_765
timestamp 1636968456
transform 1 0 71484 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_777
timestamp 1
transform 1 0 72588 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_783
timestamp 1
transform 1 0 73140 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_785
timestamp 1636968456
transform 1 0 73324 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_797
timestamp 1636968456
transform 1 0 74428 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_809
timestamp 1636968456
transform 1 0 75532 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_821
timestamp 1636968456
transform 1 0 76636 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_833
timestamp 1
transform 1 0 77740 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_839
timestamp 1
transform 1 0 78292 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_841
timestamp 1636968456
transform 1 0 78476 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_853
timestamp 1636968456
transform 1 0 79580 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_865
timestamp 1636968456
transform 1 0 80684 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_877
timestamp 1636968456
transform 1 0 81788 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_889
timestamp 1
transform 1 0 82892 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_895
timestamp 1
transform 1 0 83444 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_897
timestamp 1636968456
transform 1 0 83628 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_909
timestamp 1636968456
transform 1 0 84732 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_921
timestamp 1636968456
transform 1 0 85836 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_933
timestamp 1636968456
transform 1 0 86940 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_945
timestamp 1
transform 1 0 88044 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_951
timestamp 1
transform 1 0 88596 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_953
timestamp 1636968456
transform 1 0 88780 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_965
timestamp 1636968456
transform 1 0 89884 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_977
timestamp 1636968456
transform 1 0 90988 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_989
timestamp 1636968456
transform 1 0 92092 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_1001
timestamp 1
transform 1 0 93196 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_1007
timestamp 1
transform 1 0 93748 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1009
timestamp 1636968456
transform 1 0 93932 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1021
timestamp 1636968456
transform 1 0 95036 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1033
timestamp 1636968456
transform 1 0 96140 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1045
timestamp 1636968456
transform 1 0 97244 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_1057
timestamp 1
transform 1 0 98348 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_1063
timestamp 1
transform 1 0 98900 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1065
timestamp 1636968456
transform 1 0 99084 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1077
timestamp 1636968456
transform 1 0 100188 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1089
timestamp 1636968456
transform 1 0 101292 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1101
timestamp 1636968456
transform 1 0 102396 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_1113
timestamp 1
transform 1 0 103500 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_1119
timestamp 1
transform 1 0 104052 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1121
timestamp 1636968456
transform 1 0 104236 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1133
timestamp 1636968456
transform 1 0 105340 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1145
timestamp 1636968456
transform 1 0 106444 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1157
timestamp 1636968456
transform 1 0 107548 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_1169
timestamp 1
transform 1 0 108652 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_1175
timestamp 1
transform 1 0 109204 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1177
timestamp 1636968456
transform 1 0 109388 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1189
timestamp 1636968456
transform 1 0 110492 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1201
timestamp 1636968456
transform 1 0 111596 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1213
timestamp 1636968456
transform 1 0 112700 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_1225
timestamp 1
transform 1 0 113804 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_1231
timestamp 1
transform 1 0 114356 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1233
timestamp 1636968456
transform 1 0 114540 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1245
timestamp 1636968456
transform 1 0 115644 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1257
timestamp 1636968456
transform 1 0 116748 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_1269
timestamp 1
transform 1 0 117852 0 -1 94656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_170_3
timestamp 1636968456
transform 1 0 1380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_15
timestamp 1636968456
transform 1 0 2484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_27
timestamp 1
transform 1 0 3588 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_29
timestamp 1636968456
transform 1 0 3772 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_41
timestamp 1636968456
transform 1 0 4876 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_53
timestamp 1636968456
transform 1 0 5980 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_65
timestamp 1636968456
transform 1 0 7084 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_77
timestamp 1
transform 1 0 8188 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_83
timestamp 1
transform 1 0 8740 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_85
timestamp 1636968456
transform 1 0 8924 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_97
timestamp 1636968456
transform 1 0 10028 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_109
timestamp 1636968456
transform 1 0 11132 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_121
timestamp 1636968456
transform 1 0 12236 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_133
timestamp 1
transform 1 0 13340 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_139
timestamp 1
transform 1 0 13892 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_141
timestamp 1636968456
transform 1 0 14076 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_153
timestamp 1636968456
transform 1 0 15180 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_165
timestamp 1636968456
transform 1 0 16284 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_177
timestamp 1636968456
transform 1 0 17388 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_189
timestamp 1
transform 1 0 18492 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_195
timestamp 1
transform 1 0 19044 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_197
timestamp 1636968456
transform 1 0 19228 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_209
timestamp 1636968456
transform 1 0 20332 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_221
timestamp 1636968456
transform 1 0 21436 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_233
timestamp 1636968456
transform 1 0 22540 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_245
timestamp 1
transform 1 0 23644 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_251
timestamp 1
transform 1 0 24196 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_253
timestamp 1636968456
transform 1 0 24380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_265
timestamp 1636968456
transform 1 0 25484 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_277
timestamp 1636968456
transform 1 0 26588 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_289
timestamp 1636968456
transform 1 0 27692 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_301
timestamp 1
transform 1 0 28796 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_307
timestamp 1
transform 1 0 29348 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_309
timestamp 1636968456
transform 1 0 29532 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_321
timestamp 1636968456
transform 1 0 30636 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_333
timestamp 1636968456
transform 1 0 31740 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_345
timestamp 1636968456
transform 1 0 32844 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_357
timestamp 1
transform 1 0 33948 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_363
timestamp 1
transform 1 0 34500 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_365
timestamp 1636968456
transform 1 0 34684 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_377
timestamp 1636968456
transform 1 0 35788 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_389
timestamp 1636968456
transform 1 0 36892 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_401
timestamp 1636968456
transform 1 0 37996 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_413
timestamp 1
transform 1 0 39100 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_419
timestamp 1
transform 1 0 39652 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_421
timestamp 1636968456
transform 1 0 39836 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_433
timestamp 1636968456
transform 1 0 40940 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_445
timestamp 1636968456
transform 1 0 42044 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_457
timestamp 1636968456
transform 1 0 43148 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_469
timestamp 1
transform 1 0 44252 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_475
timestamp 1
transform 1 0 44804 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_477
timestamp 1636968456
transform 1 0 44988 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_489
timestamp 1636968456
transform 1 0 46092 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_501
timestamp 1636968456
transform 1 0 47196 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_513
timestamp 1636968456
transform 1 0 48300 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_525
timestamp 1
transform 1 0 49404 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_531
timestamp 1
transform 1 0 49956 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_533
timestamp 1636968456
transform 1 0 50140 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_545
timestamp 1636968456
transform 1 0 51244 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_557
timestamp 1636968456
transform 1 0 52348 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_569
timestamp 1636968456
transform 1 0 53452 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_581
timestamp 1
transform 1 0 54556 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_587
timestamp 1
transform 1 0 55108 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_170_589
timestamp 1
transform 1 0 55292 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_595
timestamp 1
transform 1 0 55844 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_605
timestamp 1636968456
transform 1 0 56764 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_637
timestamp 1
transform 1 0 59708 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_643
timestamp 1
transform 1 0 60260 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_645
timestamp 1636968456
transform 1 0 60444 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_170_657
timestamp 1
transform 1 0 61548 0 1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_170_661
timestamp 1
transform 1 0 61916 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_682
timestamp 1636968456
transform 1 0 63848 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_694
timestamp 1
transform 1 0 64952 0 1 94656
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_170_741
timestamp 1636968456
transform 1 0 69276 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_170_753
timestamp 1
transform 1 0 70380 0 1 94656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_170_777
timestamp 1636968456
transform 1 0 72588 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_789
timestamp 1636968456
transform 1 0 73692 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_801
timestamp 1
transform 1 0 74796 0 1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_170_809
timestamp 1
transform 1 0 75532 0 1 94656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_170_813
timestamp 1636968456
transform 1 0 75900 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_825
timestamp 1636968456
transform 1 0 77004 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_837
timestamp 1636968456
transform 1 0 78108 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_849
timestamp 1636968456
transform 1 0 79212 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_861
timestamp 1
transform 1 0 80316 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_867
timestamp 1
transform 1 0 80868 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_869
timestamp 1636968456
transform 1 0 81052 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_881
timestamp 1636968456
transform 1 0 82156 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_893
timestamp 1636968456
transform 1 0 83260 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_905
timestamp 1636968456
transform 1 0 84364 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_917
timestamp 1
transform 1 0 85468 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_923
timestamp 1
transform 1 0 86020 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_925
timestamp 1636968456
transform 1 0 86204 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_937
timestamp 1636968456
transform 1 0 87308 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_949
timestamp 1636968456
transform 1 0 88412 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_961
timestamp 1636968456
transform 1 0 89516 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_973
timestamp 1
transform 1 0 90620 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_979
timestamp 1
transform 1 0 91172 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_981
timestamp 1636968456
transform 1 0 91356 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_993
timestamp 1636968456
transform 1 0 92460 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1005
timestamp 1636968456
transform 1 0 93564 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1017
timestamp 1636968456
transform 1 0 94668 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_1029
timestamp 1
transform 1 0 95772 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1035
timestamp 1
transform 1 0 96324 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1037
timestamp 1636968456
transform 1 0 96508 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1049
timestamp 1636968456
transform 1 0 97612 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1061
timestamp 1636968456
transform 1 0 98716 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1073
timestamp 1636968456
transform 1 0 99820 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_1085
timestamp 1
transform 1 0 100924 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1091
timestamp 1
transform 1 0 101476 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1093
timestamp 1636968456
transform 1 0 101660 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1105
timestamp 1636968456
transform 1 0 102764 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1117
timestamp 1636968456
transform 1 0 103868 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1129
timestamp 1636968456
transform 1 0 104972 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_1141
timestamp 1
transform 1 0 106076 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1147
timestamp 1
transform 1 0 106628 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1149
timestamp 1636968456
transform 1 0 106812 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1161
timestamp 1636968456
transform 1 0 107916 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1173
timestamp 1636968456
transform 1 0 109020 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1185
timestamp 1636968456
transform 1 0 110124 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_1197
timestamp 1
transform 1 0 111228 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1203
timestamp 1
transform 1 0 111780 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1205
timestamp 1636968456
transform 1 0 111964 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1217
timestamp 1636968456
transform 1 0 113068 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1229
timestamp 1636968456
transform 1 0 114172 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1241
timestamp 1636968456
transform 1 0 115276 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_1253
timestamp 1
transform 1 0 116380 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1259
timestamp 1
transform 1 0 116932 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1261
timestamp 1636968456
transform 1 0 117116 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_170_1273
timestamp 1
transform 1 0 118220 0 1 94656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_171_3
timestamp 1636968456
transform 1 0 1380 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_15
timestamp 1636968456
transform 1 0 2484 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_27
timestamp 1636968456
transform 1 0 3588 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_39
timestamp 1636968456
transform 1 0 4692 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_171_51
timestamp 1
transform 1 0 5796 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_55
timestamp 1
transform 1 0 6164 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_57
timestamp 1636968456
transform 1 0 6348 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_69
timestamp 1636968456
transform 1 0 7452 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_81
timestamp 1636968456
transform 1 0 8556 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_93
timestamp 1636968456
transform 1 0 9660 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_105
timestamp 1
transform 1 0 10764 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_111
timestamp 1
transform 1 0 11316 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_113
timestamp 1636968456
transform 1 0 11500 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_125
timestamp 1636968456
transform 1 0 12604 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_137
timestamp 1636968456
transform 1 0 13708 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_149
timestamp 1636968456
transform 1 0 14812 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_161
timestamp 1
transform 1 0 15916 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_167
timestamp 1
transform 1 0 16468 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_169
timestamp 1636968456
transform 1 0 16652 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_181
timestamp 1636968456
transform 1 0 17756 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_193
timestamp 1636968456
transform 1 0 18860 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_205
timestamp 1636968456
transform 1 0 19964 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_217
timestamp 1
transform 1 0 21068 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_223
timestamp 1
transform 1 0 21620 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_225
timestamp 1636968456
transform 1 0 21804 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_237
timestamp 1636968456
transform 1 0 22908 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_249
timestamp 1636968456
transform 1 0 24012 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_261
timestamp 1636968456
transform 1 0 25116 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_273
timestamp 1
transform 1 0 26220 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_279
timestamp 1
transform 1 0 26772 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_281
timestamp 1636968456
transform 1 0 26956 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_293
timestamp 1636968456
transform 1 0 28060 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_305
timestamp 1636968456
transform 1 0 29164 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_317
timestamp 1636968456
transform 1 0 30268 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_329
timestamp 1
transform 1 0 31372 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_335
timestamp 1
transform 1 0 31924 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_337
timestamp 1636968456
transform 1 0 32108 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_349
timestamp 1636968456
transform 1 0 33212 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_361
timestamp 1636968456
transform 1 0 34316 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_373
timestamp 1636968456
transform 1 0 35420 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_385
timestamp 1
transform 1 0 36524 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_391
timestamp 1
transform 1 0 37076 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_393
timestamp 1636968456
transform 1 0 37260 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_405
timestamp 1636968456
transform 1 0 38364 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_417
timestamp 1636968456
transform 1 0 39468 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_429
timestamp 1636968456
transform 1 0 40572 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_441
timestamp 1
transform 1 0 41676 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_447
timestamp 1
transform 1 0 42228 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_449
timestamp 1636968456
transform 1 0 42412 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_461
timestamp 1636968456
transform 1 0 43516 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_473
timestamp 1636968456
transform 1 0 44620 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_485
timestamp 1636968456
transform 1 0 45724 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_497
timestamp 1
transform 1 0 46828 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_503
timestamp 1
transform 1 0 47380 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_505
timestamp 1636968456
transform 1 0 47564 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_517
timestamp 1636968456
transform 1 0 48668 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_529
timestamp 1636968456
transform 1 0 49772 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_541
timestamp 1636968456
transform 1 0 50876 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_553
timestamp 1
transform 1 0 51980 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_559
timestamp 1
transform 1 0 52532 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_561
timestamp 1636968456
transform 1 0 52716 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_573
timestamp 1636968456
transform 1 0 53820 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_585
timestamp 1
transform 1 0 54924 0 -1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_171_613
timestamp 1
transform 1 0 57500 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_617
timestamp 1636968456
transform 1 0 57868 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_629
timestamp 1
transform 1 0 58972 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_171_673
timestamp 1
transform 1 0 63020 0 -1 95744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_171_715
timestamp 1636968456
transform 1 0 66884 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_171_727
timestamp 1
transform 1 0 67988 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_769
timestamp 1636968456
transform 1 0 71852 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_171_781
timestamp 1
transform 1 0 72956 0 -1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_171_785
timestamp 1636968456
transform 1 0 73324 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_797
timestamp 1636968456
transform 1 0 74428 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_809
timestamp 1636968456
transform 1 0 75532 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_821
timestamp 1636968456
transform 1 0 76636 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_833
timestamp 1
transform 1 0 77740 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_839
timestamp 1
transform 1 0 78292 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_841
timestamp 1636968456
transform 1 0 78476 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_853
timestamp 1636968456
transform 1 0 79580 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_865
timestamp 1636968456
transform 1 0 80684 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_877
timestamp 1636968456
transform 1 0 81788 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_889
timestamp 1
transform 1 0 82892 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_895
timestamp 1
transform 1 0 83444 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_897
timestamp 1636968456
transform 1 0 83628 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_909
timestamp 1636968456
transform 1 0 84732 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_921
timestamp 1636968456
transform 1 0 85836 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_933
timestamp 1636968456
transform 1 0 86940 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_945
timestamp 1
transform 1 0 88044 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_951
timestamp 1
transform 1 0 88596 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_953
timestamp 1636968456
transform 1 0 88780 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_965
timestamp 1636968456
transform 1 0 89884 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_977
timestamp 1636968456
transform 1 0 90988 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_989
timestamp 1636968456
transform 1 0 92092 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_1001
timestamp 1
transform 1 0 93196 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_1007
timestamp 1
transform 1 0 93748 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1009
timestamp 1636968456
transform 1 0 93932 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1021
timestamp 1636968456
transform 1 0 95036 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1033
timestamp 1636968456
transform 1 0 96140 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1045
timestamp 1636968456
transform 1 0 97244 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_1057
timestamp 1
transform 1 0 98348 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_1063
timestamp 1
transform 1 0 98900 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1065
timestamp 1636968456
transform 1 0 99084 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1077
timestamp 1636968456
transform 1 0 100188 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1089
timestamp 1636968456
transform 1 0 101292 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1101
timestamp 1636968456
transform 1 0 102396 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_1113
timestamp 1
transform 1 0 103500 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_1119
timestamp 1
transform 1 0 104052 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1121
timestamp 1636968456
transform 1 0 104236 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1133
timestamp 1636968456
transform 1 0 105340 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1145
timestamp 1636968456
transform 1 0 106444 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1157
timestamp 1636968456
transform 1 0 107548 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_1169
timestamp 1
transform 1 0 108652 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_1175
timestamp 1
transform 1 0 109204 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1177
timestamp 1636968456
transform 1 0 109388 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1189
timestamp 1636968456
transform 1 0 110492 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1201
timestamp 1636968456
transform 1 0 111596 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1213
timestamp 1636968456
transform 1 0 112700 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_1225
timestamp 1
transform 1 0 113804 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_1231
timestamp 1
transform 1 0 114356 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1233
timestamp 1636968456
transform 1 0 114540 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1245
timestamp 1636968456
transform 1 0 115644 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1257
timestamp 1636968456
transform 1 0 116748 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_1269
timestamp 1
transform 1 0 117852 0 -1 95744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_172_3
timestamp 1636968456
transform 1 0 1380 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_15
timestamp 1636968456
transform 1 0 2484 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_27
timestamp 1
transform 1 0 3588 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_29
timestamp 1636968456
transform 1 0 3772 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_41
timestamp 1636968456
transform 1 0 4876 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_53
timestamp 1636968456
transform 1 0 5980 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_65
timestamp 1636968456
transform 1 0 7084 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_77
timestamp 1
transform 1 0 8188 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_83
timestamp 1
transform 1 0 8740 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_85
timestamp 1636968456
transform 1 0 8924 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_97
timestamp 1636968456
transform 1 0 10028 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_109
timestamp 1636968456
transform 1 0 11132 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_121
timestamp 1636968456
transform 1 0 12236 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_133
timestamp 1
transform 1 0 13340 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_139
timestamp 1
transform 1 0 13892 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_141
timestamp 1636968456
transform 1 0 14076 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_153
timestamp 1636968456
transform 1 0 15180 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_165
timestamp 1636968456
transform 1 0 16284 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_177
timestamp 1636968456
transform 1 0 17388 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_189
timestamp 1
transform 1 0 18492 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_195
timestamp 1
transform 1 0 19044 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_197
timestamp 1636968456
transform 1 0 19228 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_209
timestamp 1636968456
transform 1 0 20332 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_221
timestamp 1636968456
transform 1 0 21436 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_233
timestamp 1636968456
transform 1 0 22540 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_245
timestamp 1
transform 1 0 23644 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_251
timestamp 1
transform 1 0 24196 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_253
timestamp 1636968456
transform 1 0 24380 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_265
timestamp 1636968456
transform 1 0 25484 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_277
timestamp 1636968456
transform 1 0 26588 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_289
timestamp 1636968456
transform 1 0 27692 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_301
timestamp 1
transform 1 0 28796 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_307
timestamp 1
transform 1 0 29348 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_309
timestamp 1636968456
transform 1 0 29532 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_321
timestamp 1636968456
transform 1 0 30636 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_333
timestamp 1636968456
transform 1 0 31740 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_345
timestamp 1636968456
transform 1 0 32844 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_357
timestamp 1
transform 1 0 33948 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_363
timestamp 1
transform 1 0 34500 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_365
timestamp 1636968456
transform 1 0 34684 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_377
timestamp 1636968456
transform 1 0 35788 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_389
timestamp 1636968456
transform 1 0 36892 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_401
timestamp 1636968456
transform 1 0 37996 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_413
timestamp 1
transform 1 0 39100 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_419
timestamp 1
transform 1 0 39652 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_421
timestamp 1636968456
transform 1 0 39836 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_433
timestamp 1636968456
transform 1 0 40940 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_445
timestamp 1636968456
transform 1 0 42044 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_457
timestamp 1636968456
transform 1 0 43148 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_469
timestamp 1
transform 1 0 44252 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_475
timestamp 1
transform 1 0 44804 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_477
timestamp 1636968456
transform 1 0 44988 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_489
timestamp 1636968456
transform 1 0 46092 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_501
timestamp 1636968456
transform 1 0 47196 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_513
timestamp 1636968456
transform 1 0 48300 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_525
timestamp 1
transform 1 0 49404 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_531
timestamp 1
transform 1 0 49956 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_533
timestamp 1636968456
transform 1 0 50140 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_545
timestamp 1636968456
transform 1 0 51244 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_557
timestamp 1636968456
transform 1 0 52348 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_569
timestamp 1636968456
transform 1 0 53452 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_581
timestamp 1
transform 1 0 54556 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_587
timestamp 1
transform 1 0 55108 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_589
timestamp 1636968456
transform 1 0 55292 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_172_601
timestamp 1
transform 1 0 56396 0 1 95744
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_172_625
timestamp 1636968456
transform 1 0 58604 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_637
timestamp 1
transform 1 0 59708 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_643
timestamp 1
transform 1 0 60260 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_645
timestamp 1636968456
transform 1 0 60444 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_657
timestamp 1636968456
transform 1 0 61548 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_669
timestamp 1636968456
transform 1 0 62652 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_681
timestamp 1636968456
transform 1 0 63756 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_693
timestamp 1
transform 1 0 64860 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_699
timestamp 1
transform 1 0 65412 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_172_701
timestamp 1
transform 1 0 65596 0 1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_172_705
timestamp 1
transform 1 0 65964 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_726
timestamp 1636968456
transform 1 0 67896 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_738
timestamp 1636968456
transform 1 0 69000 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_750
timestamp 1
transform 1 0 70104 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_172_757
timestamp 1
transform 1 0 70748 0 1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_172_765
timestamp 1
transform 1 0 71484 0 1 95744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_172_787
timestamp 1636968456
transform 1 0 73508 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_799
timestamp 1636968456
transform 1 0 74612 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_811
timestamp 1
transform 1 0 75716 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_813
timestamp 1636968456
transform 1 0 75900 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_825
timestamp 1636968456
transform 1 0 77004 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_837
timestamp 1636968456
transform 1 0 78108 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_849
timestamp 1636968456
transform 1 0 79212 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_861
timestamp 1
transform 1 0 80316 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_867
timestamp 1
transform 1 0 80868 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_869
timestamp 1636968456
transform 1 0 81052 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_881
timestamp 1636968456
transform 1 0 82156 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_893
timestamp 1636968456
transform 1 0 83260 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_905
timestamp 1636968456
transform 1 0 84364 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_917
timestamp 1
transform 1 0 85468 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_923
timestamp 1
transform 1 0 86020 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_925
timestamp 1636968456
transform 1 0 86204 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_937
timestamp 1636968456
transform 1 0 87308 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_949
timestamp 1636968456
transform 1 0 88412 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_961
timestamp 1636968456
transform 1 0 89516 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_973
timestamp 1
transform 1 0 90620 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_979
timestamp 1
transform 1 0 91172 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_981
timestamp 1636968456
transform 1 0 91356 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_993
timestamp 1636968456
transform 1 0 92460 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1005
timestamp 1636968456
transform 1 0 93564 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1017
timestamp 1636968456
transform 1 0 94668 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_1029
timestamp 1
transform 1 0 95772 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_1035
timestamp 1
transform 1 0 96324 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1037
timestamp 1636968456
transform 1 0 96508 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1049
timestamp 1636968456
transform 1 0 97612 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1061
timestamp 1636968456
transform 1 0 98716 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1073
timestamp 1636968456
transform 1 0 99820 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_1085
timestamp 1
transform 1 0 100924 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_1091
timestamp 1
transform 1 0 101476 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1093
timestamp 1636968456
transform 1 0 101660 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1105
timestamp 1636968456
transform 1 0 102764 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1117
timestamp 1636968456
transform 1 0 103868 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1129
timestamp 1636968456
transform 1 0 104972 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_1141
timestamp 1
transform 1 0 106076 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_1147
timestamp 1
transform 1 0 106628 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1149
timestamp 1636968456
transform 1 0 106812 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1161
timestamp 1636968456
transform 1 0 107916 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1173
timestamp 1636968456
transform 1 0 109020 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1185
timestamp 1636968456
transform 1 0 110124 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_1197
timestamp 1
transform 1 0 111228 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_1203
timestamp 1
transform 1 0 111780 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1205
timestamp 1636968456
transform 1 0 111964 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1217
timestamp 1636968456
transform 1 0 113068 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1229
timestamp 1636968456
transform 1 0 114172 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1241
timestamp 1636968456
transform 1 0 115276 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_1253
timestamp 1
transform 1 0 116380 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_1259
timestamp 1
transform 1 0 116932 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1261
timestamp 1636968456
transform 1 0 117116 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_172_1273
timestamp 1
transform 1 0 118220 0 1 95744
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_173_3
timestamp 1636968456
transform 1 0 1380 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_15
timestamp 1636968456
transform 1 0 2484 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_27
timestamp 1636968456
transform 1 0 3588 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_39
timestamp 1636968456
transform 1 0 4692 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_173_51
timestamp 1
transform 1 0 5796 0 -1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_173_55
timestamp 1
transform 1 0 6164 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_57
timestamp 1636968456
transform 1 0 6348 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_69
timestamp 1636968456
transform 1 0 7452 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_81
timestamp 1636968456
transform 1 0 8556 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_93
timestamp 1636968456
transform 1 0 9660 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_105
timestamp 1
transform 1 0 10764 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_111
timestamp 1
transform 1 0 11316 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_113
timestamp 1636968456
transform 1 0 11500 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_125
timestamp 1636968456
transform 1 0 12604 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_137
timestamp 1636968456
transform 1 0 13708 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_149
timestamp 1636968456
transform 1 0 14812 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_161
timestamp 1
transform 1 0 15916 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_167
timestamp 1
transform 1 0 16468 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_169
timestamp 1636968456
transform 1 0 16652 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_181
timestamp 1636968456
transform 1 0 17756 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_193
timestamp 1636968456
transform 1 0 18860 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_205
timestamp 1636968456
transform 1 0 19964 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_217
timestamp 1
transform 1 0 21068 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_223
timestamp 1
transform 1 0 21620 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_225
timestamp 1636968456
transform 1 0 21804 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_237
timestamp 1636968456
transform 1 0 22908 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_249
timestamp 1636968456
transform 1 0 24012 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_261
timestamp 1636968456
transform 1 0 25116 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_273
timestamp 1
transform 1 0 26220 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_279
timestamp 1
transform 1 0 26772 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_281
timestamp 1636968456
transform 1 0 26956 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_293
timestamp 1636968456
transform 1 0 28060 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_305
timestamp 1636968456
transform 1 0 29164 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_317
timestamp 1636968456
transform 1 0 30268 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_329
timestamp 1
transform 1 0 31372 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_335
timestamp 1
transform 1 0 31924 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_337
timestamp 1636968456
transform 1 0 32108 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_349
timestamp 1636968456
transform 1 0 33212 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_361
timestamp 1636968456
transform 1 0 34316 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_373
timestamp 1636968456
transform 1 0 35420 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_385
timestamp 1
transform 1 0 36524 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_391
timestamp 1
transform 1 0 37076 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_393
timestamp 1636968456
transform 1 0 37260 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_405
timestamp 1636968456
transform 1 0 38364 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_417
timestamp 1636968456
transform 1 0 39468 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_429
timestamp 1636968456
transform 1 0 40572 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_441
timestamp 1
transform 1 0 41676 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_447
timestamp 1
transform 1 0 42228 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_449
timestamp 1636968456
transform 1 0 42412 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_461
timestamp 1636968456
transform 1 0 43516 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_473
timestamp 1636968456
transform 1 0 44620 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_485
timestamp 1636968456
transform 1 0 45724 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_497
timestamp 1
transform 1 0 46828 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_503
timestamp 1
transform 1 0 47380 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_505
timestamp 1636968456
transform 1 0 47564 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_517
timestamp 1636968456
transform 1 0 48668 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_529
timestamp 1636968456
transform 1 0 49772 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_541
timestamp 1636968456
transform 1 0 50876 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_553
timestamp 1
transform 1 0 51980 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_559
timestamp 1
transform 1 0 52532 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_561
timestamp 1636968456
transform 1 0 52716 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_573
timestamp 1636968456
transform 1 0 53820 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_585
timestamp 1
transform 1 0 54924 0 -1 96832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_173_593
timestamp 1
transform 1 0 55660 0 -1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_173_601
timestamp 1636968456
transform 1 0 56396 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_173_613
timestamp 1
transform 1 0 57500 0 -1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_173_617
timestamp 1636968456
transform 1 0 57868 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_629
timestamp 1636968456
transform 1 0 58972 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_641
timestamp 1636968456
transform 1 0 60076 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_653
timestamp 1636968456
transform 1 0 61180 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_665
timestamp 1
transform 1 0 62284 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_671
timestamp 1
transform 1 0 62836 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_673
timestamp 1636968456
transform 1 0 63020 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_685
timestamp 1636968456
transform 1 0 64124 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_697
timestamp 1636968456
transform 1 0 65228 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_709
timestamp 1636968456
transform 1 0 66332 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_721
timestamp 1
transform 1 0 67436 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_727
timestamp 1
transform 1 0 67988 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_173_729
timestamp 1
transform 1 0 68172 0 -1 96832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_173_737
timestamp 1
transform 1 0 68908 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_742
timestamp 1636968456
transform 1 0 69368 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_754
timestamp 1636968456
transform 1 0 70472 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_766
timestamp 1636968456
transform 1 0 71576 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_778
timestamp 1
transform 1 0 72680 0 -1 96832
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_173_785
timestamp 1636968456
transform 1 0 73324 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_797
timestamp 1636968456
transform 1 0 74428 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_809
timestamp 1636968456
transform 1 0 75532 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_821
timestamp 1636968456
transform 1 0 76636 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_833
timestamp 1
transform 1 0 77740 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_839
timestamp 1
transform 1 0 78292 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_841
timestamp 1636968456
transform 1 0 78476 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_853
timestamp 1636968456
transform 1 0 79580 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_865
timestamp 1636968456
transform 1 0 80684 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_877
timestamp 1636968456
transform 1 0 81788 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_889
timestamp 1
transform 1 0 82892 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_895
timestamp 1
transform 1 0 83444 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_897
timestamp 1636968456
transform 1 0 83628 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_909
timestamp 1636968456
transform 1 0 84732 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_921
timestamp 1636968456
transform 1 0 85836 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_933
timestamp 1636968456
transform 1 0 86940 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_945
timestamp 1
transform 1 0 88044 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_951
timestamp 1
transform 1 0 88596 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_953
timestamp 1636968456
transform 1 0 88780 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_965
timestamp 1636968456
transform 1 0 89884 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_977
timestamp 1636968456
transform 1 0 90988 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_989
timestamp 1636968456
transform 1 0 92092 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_1001
timestamp 1
transform 1 0 93196 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_1007
timestamp 1
transform 1 0 93748 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1009
timestamp 1636968456
transform 1 0 93932 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1021
timestamp 1636968456
transform 1 0 95036 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1033
timestamp 1636968456
transform 1 0 96140 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1045
timestamp 1636968456
transform 1 0 97244 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_1057
timestamp 1
transform 1 0 98348 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_1063
timestamp 1
transform 1 0 98900 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1065
timestamp 1636968456
transform 1 0 99084 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1077
timestamp 1636968456
transform 1 0 100188 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1089
timestamp 1636968456
transform 1 0 101292 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1101
timestamp 1636968456
transform 1 0 102396 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_1113
timestamp 1
transform 1 0 103500 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_1119
timestamp 1
transform 1 0 104052 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1121
timestamp 1636968456
transform 1 0 104236 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1133
timestamp 1636968456
transform 1 0 105340 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1145
timestamp 1636968456
transform 1 0 106444 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1157
timestamp 1636968456
transform 1 0 107548 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_1169
timestamp 1
transform 1 0 108652 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_1175
timestamp 1
transform 1 0 109204 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1177
timestamp 1636968456
transform 1 0 109388 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1189
timestamp 1636968456
transform 1 0 110492 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1201
timestamp 1636968456
transform 1 0 111596 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1213
timestamp 1636968456
transform 1 0 112700 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_1225
timestamp 1
transform 1 0 113804 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_1231
timestamp 1
transform 1 0 114356 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1233
timestamp 1636968456
transform 1 0 114540 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1245
timestamp 1636968456
transform 1 0 115644 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1257
timestamp 1636968456
transform 1 0 116748 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_1269
timestamp 1
transform 1 0 117852 0 -1 96832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_174_3
timestamp 1636968456
transform 1 0 1380 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_15
timestamp 1636968456
transform 1 0 2484 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_174_27
timestamp 1
transform 1 0 3588 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_29
timestamp 1636968456
transform 1 0 3772 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_41
timestamp 1636968456
transform 1 0 4876 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_53
timestamp 1
transform 1 0 5980 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_57
timestamp 1636968456
transform 1 0 6348 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_69
timestamp 1636968456
transform 1 0 7452 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_81
timestamp 1
transform 1 0 8556 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_85
timestamp 1636968456
transform 1 0 8924 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_97
timestamp 1636968456
transform 1 0 10028 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_109
timestamp 1
transform 1 0 11132 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_113
timestamp 1636968456
transform 1 0 11500 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_125
timestamp 1636968456
transform 1 0 12604 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_137
timestamp 1
transform 1 0 13708 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_141
timestamp 1636968456
transform 1 0 14076 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_153
timestamp 1636968456
transform 1 0 15180 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_165
timestamp 1
transform 1 0 16284 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_169
timestamp 1636968456
transform 1 0 16652 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_181
timestamp 1636968456
transform 1 0 17756 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_193
timestamp 1
transform 1 0 18860 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_197
timestamp 1636968456
transform 1 0 19228 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_209
timestamp 1636968456
transform 1 0 20332 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_221
timestamp 1
transform 1 0 21436 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_225
timestamp 1636968456
transform 1 0 21804 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_237
timestamp 1636968456
transform 1 0 22908 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_249
timestamp 1
transform 1 0 24012 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_253
timestamp 1636968456
transform 1 0 24380 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_265
timestamp 1636968456
transform 1 0 25484 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_277
timestamp 1
transform 1 0 26588 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_281
timestamp 1636968456
transform 1 0 26956 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_293
timestamp 1636968456
transform 1 0 28060 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_305
timestamp 1
transform 1 0 29164 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_309
timestamp 1636968456
transform 1 0 29532 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_321
timestamp 1636968456
transform 1 0 30636 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_333
timestamp 1
transform 1 0 31740 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_337
timestamp 1636968456
transform 1 0 32108 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_349
timestamp 1636968456
transform 1 0 33212 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_361
timestamp 1
transform 1 0 34316 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_365
timestamp 1636968456
transform 1 0 34684 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_377
timestamp 1636968456
transform 1 0 35788 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_389
timestamp 1
transform 1 0 36892 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_393
timestamp 1636968456
transform 1 0 37260 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_405
timestamp 1636968456
transform 1 0 38364 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_417
timestamp 1
transform 1 0 39468 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_421
timestamp 1636968456
transform 1 0 39836 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_433
timestamp 1636968456
transform 1 0 40940 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_445
timestamp 1
transform 1 0 42044 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_449
timestamp 1636968456
transform 1 0 42412 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_461
timestamp 1636968456
transform 1 0 43516 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_473
timestamp 1
transform 1 0 44620 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_477
timestamp 1636968456
transform 1 0 44988 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_489
timestamp 1636968456
transform 1 0 46092 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_501
timestamp 1
transform 1 0 47196 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_505
timestamp 1636968456
transform 1 0 47564 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_517
timestamp 1636968456
transform 1 0 48668 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_529
timestamp 1
transform 1 0 49772 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_533
timestamp 1636968456
transform 1 0 50140 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_545
timestamp 1636968456
transform 1 0 51244 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_557
timestamp 1
transform 1 0 52348 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_561
timestamp 1636968456
transform 1 0 52716 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_573
timestamp 1636968456
transform 1 0 53820 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_585
timestamp 1
transform 1 0 54924 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_174_589
timestamp 1
transform 1 0 55292 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_174_615
timestamp 1
transform 1 0 57684 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_174_623
timestamp 1
transform 1 0 58420 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_174_630
timestamp 1
transform 1 0 59064 0 1 96832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_174_638
timestamp 1
transform 1 0 59800 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_174_645
timestamp 1
transform 1 0 60444 0 1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_174_651
timestamp 1636968456
transform 1 0 60996 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_174_663
timestamp 1
transform 1 0 62100 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_174_667
timestamp 1
transform 1 0 62468 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_174_673
timestamp 1
transform 1 0 63020 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_174_679
timestamp 1
transform 1 0 63572 0 1 96832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_174_687
timestamp 1
transform 1 0 64308 0 1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_174_693
timestamp 1
transform 1 0 64860 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_701
timestamp 1636968456
transform 1 0 65596 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_174_713
timestamp 1
transform 1 0 66700 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_174_721
timestamp 1
transform 1 0 67436 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_174_749
timestamp 1
transform 1 0 70012 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_174_757
timestamp 1
transform 1 0 70748 0 1 96832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_174_765
timestamp 1
transform 1 0 71484 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_174_770
timestamp 1
transform 1 0 71944 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_174_777
timestamp 1
transform 1 0 72588 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_783
timestamp 1
transform 1 0 73140 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_785
timestamp 1
transform 1 0 73324 0 1 96832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_174_793
timestamp 1
transform 1 0 74060 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_798
timestamp 1636968456
transform 1 0 74520 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_174_810
timestamp 1
transform 1 0 75624 0 1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_174_813
timestamp 1636968456
transform 1 0 75900 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_825
timestamp 1636968456
transform 1 0 77004 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_837
timestamp 1
transform 1 0 78108 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_841
timestamp 1636968456
transform 1 0 78476 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_853
timestamp 1636968456
transform 1 0 79580 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_865
timestamp 1
transform 1 0 80684 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_869
timestamp 1636968456
transform 1 0 81052 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_881
timestamp 1636968456
transform 1 0 82156 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_893
timestamp 1
transform 1 0 83260 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_897
timestamp 1636968456
transform 1 0 83628 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_909
timestamp 1636968456
transform 1 0 84732 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_921
timestamp 1
transform 1 0 85836 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_925
timestamp 1636968456
transform 1 0 86204 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_937
timestamp 1636968456
transform 1 0 87308 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_949
timestamp 1
transform 1 0 88412 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_953
timestamp 1636968456
transform 1 0 88780 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_965
timestamp 1636968456
transform 1 0 89884 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_977
timestamp 1
transform 1 0 90988 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_981
timestamp 1636968456
transform 1 0 91356 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_993
timestamp 1636968456
transform 1 0 92460 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1005
timestamp 1
transform 1 0 93564 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1009
timestamp 1636968456
transform 1 0 93932 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1021
timestamp 1636968456
transform 1 0 95036 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1033
timestamp 1
transform 1 0 96140 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1037
timestamp 1636968456
transform 1 0 96508 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1049
timestamp 1636968456
transform 1 0 97612 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1061
timestamp 1
transform 1 0 98716 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1065
timestamp 1636968456
transform 1 0 99084 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1077
timestamp 1636968456
transform 1 0 100188 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1089
timestamp 1
transform 1 0 101292 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1093
timestamp 1636968456
transform 1 0 101660 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1105
timestamp 1636968456
transform 1 0 102764 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1117
timestamp 1
transform 1 0 103868 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1121
timestamp 1636968456
transform 1 0 104236 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1133
timestamp 1636968456
transform 1 0 105340 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1145
timestamp 1
transform 1 0 106444 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_174_1149
timestamp 1
transform 1 0 106812 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_1155
timestamp 1
transform 1 0 107364 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1164
timestamp 1636968456
transform 1 0 108192 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1177
timestamp 1636968456
transform 1 0 109388 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1189
timestamp 1636968456
transform 1 0 110492 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1201
timestamp 1
transform 1 0 111596 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1205
timestamp 1636968456
transform 1 0 111964 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1217
timestamp 1636968456
transform 1 0 113068 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1229
timestamp 1
transform 1 0 114172 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1233
timestamp 1636968456
transform 1 0 114540 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1245
timestamp 1636968456
transform 1 0 115644 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_174_1257
timestamp 1
transform 1 0 116748 0 1 96832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1261
timestamp 1636968456
transform 1 0 117116 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_174_1273
timestamp 1
transform 1 0 118220 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 1656 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1656 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 1656 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 1656 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform -1 0 1656 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 1656 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1
transform -1 0 117208 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1
transform 1 0 118036 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1
transform 1 0 118312 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1
transform 1 0 118036 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1
transform 1 0 31648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1
transform 1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1
transform 1 0 44528 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1
transform 1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1
transform -1 0 46736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1
transform 1 0 47748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1
transform 1 0 49036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1
transform -1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1
transform -1 0 35144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1
transform 1 0 37444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1
transform -1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1
transform 1 0 40020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1
transform 1 0 41952 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1
transform 1 0 50324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1
transform 1 0 61916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1
transform 1 0 63204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1
transform -1 0 64124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1
transform -1 0 65412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1
transform -1 0 66700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1
transform 1 0 67712 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1
transform 1 0 51612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1
transform -1 0 52532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1
transform 1 0 53544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1
transform -1 0 55108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1
transform 1 0 56120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1
transform 1 0 57408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1
transform -1 0 58328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1
transform -1 0 59616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1
transform -1 0 60904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1
transform 1 0 118312 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1
transform 1 0 118312 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1
transform 1 0 118312 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1
transform 1 0 118036 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input50
timestamp 1
transform 1 0 107640 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  load_slew78
timestamp 1
transform -1 0 109020 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew79
timestamp 1
transform 1 0 109296 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew80
timestamp 1
transform 1 0 109020 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew81
timestamp 1
transform 1 0 109020 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew82
timestamp 1
transform -1 0 109296 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew83
timestamp 1
transform -1 0 108652 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew84
timestamp 1
transform 1 0 109756 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew85
timestamp 1
transform -1 0 108560 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew86
timestamp 1
transform -1 0 109756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew87
timestamp 1
transform 1 0 109756 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew88
timestamp 1
transform 1 0 110860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew89
timestamp 1
transform -1 0 110492 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew90
timestamp 1
transform -1 0 110308 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  load_slew91
timestamp 1
transform -1 0 110032 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  load_slew92
timestamp 1
transform -1 0 110216 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew93
timestamp 1
transform 1 0 110216 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew94
timestamp 1
transform -1 0 110216 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  load_slew95
timestamp 1
transform -1 0 110584 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew96
timestamp 1
transform -1 0 110216 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew99
timestamp 1
transform -1 0 109940 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  load_slew100
timestamp 1
transform -1 0 109020 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  load_slew101
timestamp 1
transform 1 0 109020 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  max_cap67
timestamp 1
transform -1 0 115644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap68
timestamp 1
transform -1 0 114448 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap70
timestamp 1
transform 1 0 117852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap71
timestamp 1
transform -1 0 115552 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap72
timestamp 1
transform -1 0 112148 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap75
timestamp 1
transform -1 0 115736 0 1 27200
box -38 -48 314 592
use sky130_sram_1kbyte_1rw1r_32x256_8  mem_i .volare/volare/sky130/versions/0fe599b2afb6708d281543108caf8310912f54af/sky130A/libs.ref/sky130_sram_macros/mag
timestamp 1723858470
transform 1 0 10000 0 1 10000
box 0 0 95956 79500
use sky130_fd_sc_hd__conb_1  mem_i_113
timestamp 1
transform -1 0 108560 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i_114
timestamp 1
transform 1 0 7360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i_115
timestamp 1
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i_116
timestamp 1
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i_117
timestamp 1
transform 1 0 29532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i_118
timestamp 1
transform 1 0 30176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1
transform -1 0 55844 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1
transform -1 0 68080 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1
transform -1 0 69368 0 -1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1
transform 1 0 70288 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1
transform -1 0 71944 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1
transform -1 0 72588 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1
transform 1 0 74152 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1
transform -1 0 58236 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1
transform -1 0 59064 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1
transform -1 0 60996 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1
transform -1 0 60352 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1
transform -1 0 62928 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1
transform -1 0 63572 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1
transform -1 0 64860 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1
transform -1 0 65504 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1
transform -1 0 67436 0 1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_175
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 118864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_176
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 118864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_177
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 118864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_178
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 118864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_179
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 118864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_180
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 118864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_181
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 118864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_182
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 118864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_183
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 118864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_184
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 118864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_349
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_659
timestamp 1
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_350
timestamp 1
transform 1 0 108008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_20
timestamp 1
transform -1 0 118864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_185
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_505
timestamp 1
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_351
timestamp 1
transform 1 0 108008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_21
timestamp 1
transform -1 0 118864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_186
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_506
timestamp 1
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_352
timestamp 1
transform 1 0 108008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_22
timestamp 1
transform -1 0 118864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_187
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_507
timestamp 1
transform -1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_353
timestamp 1
transform 1 0 108008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_23
timestamp 1
transform -1 0 118864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_188
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_508
timestamp 1
transform -1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_354
timestamp 1
transform 1 0 108008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_24
timestamp 1
transform -1 0 118864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_189
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_509
timestamp 1
transform -1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_355
timestamp 1
transform 1 0 108008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_25
timestamp 1
transform -1 0 118864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_190
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_510
timestamp 1
transform -1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_356
timestamp 1
transform 1 0 108008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_26
timestamp 1
transform -1 0 118864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_191
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_511
timestamp 1
transform -1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_357
timestamp 1
transform 1 0 108008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_27
timestamp 1
transform -1 0 118864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_192
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_512
timestamp 1
transform -1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_358
timestamp 1
transform 1 0 108008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_28
timestamp 1
transform -1 0 118864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_193
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_513
timestamp 1
transform -1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_359
timestamp 1
transform 1 0 108008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_29
timestamp 1
transform -1 0 118864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_194
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_514
timestamp 1
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_360
timestamp 1
transform 1 0 108008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_30
timestamp 1
transform -1 0 118864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_195
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_515
timestamp 1
transform -1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_361
timestamp 1
transform 1 0 108008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_31
timestamp 1
transform -1 0 118864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_196
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_516
timestamp 1
transform -1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_362
timestamp 1
transform 1 0 108008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_32
timestamp 1
transform -1 0 118864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_197
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_517
timestamp 1
transform -1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_363
timestamp 1
transform 1 0 108008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_33
timestamp 1
transform -1 0 118864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_198
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_518
timestamp 1
transform -1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_364
timestamp 1
transform 1 0 108008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_34
timestamp 1
transform -1 0 118864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_199
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_519
timestamp 1
transform -1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_365
timestamp 1
transform 1 0 108008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_35
timestamp 1
transform -1 0 118864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_200
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_520
timestamp 1
transform -1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_366
timestamp 1
transform 1 0 108008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_36
timestamp 1
transform -1 0 118864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_201
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_521
timestamp 1
transform -1 0 7912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_367
timestamp 1
transform 1 0 108008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_37
timestamp 1
transform -1 0 118864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_202
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_522
timestamp 1
transform -1 0 7912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_368
timestamp 1
transform 1 0 108008 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_38
timestamp 1
transform -1 0 118864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_203
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_523
timestamp 1
transform -1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_369
timestamp 1
transform 1 0 108008 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_39
timestamp 1
transform -1 0 118864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_204
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_524
timestamp 1
transform -1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_370
timestamp 1
transform 1 0 108008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_40
timestamp 1
transform -1 0 118864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_205
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_525
timestamp 1
transform -1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_371
timestamp 1
transform 1 0 108008 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_41
timestamp 1
transform -1 0 118864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_206
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_526
timestamp 1
transform -1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_372
timestamp 1
transform 1 0 108008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_42
timestamp 1
transform -1 0 118864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_207
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_527
timestamp 1
transform -1 0 7912 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_373
timestamp 1
transform 1 0 108008 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_43
timestamp 1
transform -1 0 118864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_208
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_528
timestamp 1
transform -1 0 7912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_374
timestamp 1
transform 1 0 108008 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_44
timestamp 1
transform -1 0 118864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_209
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_529
timestamp 1
transform -1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_375
timestamp 1
transform 1 0 108008 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_45
timestamp 1
transform -1 0 118864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_210
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_530
timestamp 1
transform -1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_376
timestamp 1
transform 1 0 108008 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_46
timestamp 1
transform -1 0 118864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_211
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_531
timestamp 1
transform -1 0 7912 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_377
timestamp 1
transform 1 0 108008 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_47
timestamp 1
transform -1 0 118864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_212
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_532
timestamp 1
transform -1 0 7912 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_378
timestamp 1
transform 1 0 108008 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_48
timestamp 1
transform -1 0 118864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_213
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_533
timestamp 1
transform -1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_379
timestamp 1
transform 1 0 108008 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_49
timestamp 1
transform -1 0 118864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_214
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_534
timestamp 1
transform -1 0 7912 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_380
timestamp 1
transform 1 0 108008 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_50
timestamp 1
transform -1 0 118864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_215
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_535
timestamp 1
transform -1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_381
timestamp 1
transform 1 0 108008 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_51
timestamp 1
transform -1 0 118864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_216
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_536
timestamp 1
transform -1 0 7912 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_382
timestamp 1
transform 1 0 108008 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_52
timestamp 1
transform -1 0 118864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_217
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_537
timestamp 1
transform -1 0 7912 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_383
timestamp 1
transform 1 0 108008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_53
timestamp 1
transform -1 0 118864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_218
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_538
timestamp 1
transform -1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_384
timestamp 1
transform 1 0 108008 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_54
timestamp 1
transform -1 0 118864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_219
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_539
timestamp 1
transform -1 0 7912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_385
timestamp 1
transform 1 0 108008 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_55
timestamp 1
transform -1 0 118864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_220
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_540
timestamp 1
transform -1 0 7912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_386
timestamp 1
transform 1 0 108008 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_56
timestamp 1
transform -1 0 118864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_221
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_541
timestamp 1
transform -1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_387
timestamp 1
transform 1 0 108008 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_57
timestamp 1
transform -1 0 118864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_222
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_542
timestamp 1
transform -1 0 7912 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_388
timestamp 1
transform 1 0 108008 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_58
timestamp 1
transform -1 0 118864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_223
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_543
timestamp 1
transform -1 0 7912 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_389
timestamp 1
transform 1 0 108008 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_59
timestamp 1
transform -1 0 118864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_224
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_544
timestamp 1
transform -1 0 7912 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_390
timestamp 1
transform 1 0 108008 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_60
timestamp 1
transform -1 0 118864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_225
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_545
timestamp 1
transform -1 0 7912 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_391
timestamp 1
transform 1 0 108008 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_61
timestamp 1
transform -1 0 118864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_226
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_546
timestamp 1
transform -1 0 7912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_392
timestamp 1
transform 1 0 108008 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_62
timestamp 1
transform -1 0 118864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_227
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_547
timestamp 1
transform -1 0 7912 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_393
timestamp 1
transform 1 0 108008 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_63
timestamp 1
transform -1 0 118864 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_228
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_548
timestamp 1
transform -1 0 7912 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_394
timestamp 1
transform 1 0 108008 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_64
timestamp 1
transform -1 0 118864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_229
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_549
timestamp 1
transform -1 0 7912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_395
timestamp 1
transform 1 0 108008 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_65
timestamp 1
transform -1 0 118864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_230
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_550
timestamp 1
transform -1 0 7912 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_396
timestamp 1
transform 1 0 108008 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_66
timestamp 1
transform -1 0 118864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_231
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_551
timestamp 1
transform -1 0 7912 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_397
timestamp 1
transform 1 0 108008 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_67
timestamp 1
transform -1 0 118864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_232
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_552
timestamp 1
transform -1 0 7912 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_398
timestamp 1
transform 1 0 108008 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_68
timestamp 1
transform -1 0 118864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_233
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_553
timestamp 1
transform -1 0 7912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_399
timestamp 1
transform 1 0 108008 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_69
timestamp 1
transform -1 0 118864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_234
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_554
timestamp 1
transform -1 0 7912 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_400
timestamp 1
transform 1 0 108008 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_70
timestamp 1
transform -1 0 118864 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_235
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_555
timestamp 1
transform -1 0 7912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_401
timestamp 1
transform 1 0 108008 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_71
timestamp 1
transform -1 0 118864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_236
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_556
timestamp 1
transform -1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_402
timestamp 1
transform 1 0 108008 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_72
timestamp 1
transform -1 0 118864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_237
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_557
timestamp 1
transform -1 0 7912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_403
timestamp 1
transform 1 0 108008 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_73
timestamp 1
transform -1 0 118864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_238
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_558
timestamp 1
transform -1 0 7912 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_404
timestamp 1
transform 1 0 108008 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_74
timestamp 1
transform -1 0 118864 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_239
timestamp 1
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_559
timestamp 1
transform -1 0 7912 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_405
timestamp 1
transform 1 0 108008 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_75
timestamp 1
transform -1 0 118864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_240
timestamp 1
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_560
timestamp 1
transform -1 0 7912 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_406
timestamp 1
transform 1 0 108008 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_76
timestamp 1
transform -1 0 118864 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_241
timestamp 1
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_561
timestamp 1
transform -1 0 7912 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_407
timestamp 1
transform 1 0 108008 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_77
timestamp 1
transform -1 0 118864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_242
timestamp 1
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_562
timestamp 1
transform -1 0 7912 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_408
timestamp 1
transform 1 0 108008 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_78
timestamp 1
transform -1 0 118864 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_243
timestamp 1
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_563
timestamp 1
transform -1 0 7912 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_409
timestamp 1
transform 1 0 108008 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_79
timestamp 1
transform -1 0 118864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_244
timestamp 1
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_564
timestamp 1
transform -1 0 7912 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_410
timestamp 1
transform 1 0 108008 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_80
timestamp 1
transform -1 0 118864 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_245
timestamp 1
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_565
timestamp 1
transform -1 0 7912 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_411
timestamp 1
transform 1 0 108008 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_81
timestamp 1
transform -1 0 118864 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_246
timestamp 1
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_566
timestamp 1
transform -1 0 7912 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_412
timestamp 1
transform 1 0 108008 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_82
timestamp 1
transform -1 0 118864 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_247
timestamp 1
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_567
timestamp 1
transform -1 0 7912 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_413
timestamp 1
transform 1 0 108008 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_83
timestamp 1
transform -1 0 118864 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_248
timestamp 1
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_568
timestamp 1
transform -1 0 7912 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_414
timestamp 1
transform 1 0 108008 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_84
timestamp 1
transform -1 0 118864 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_249
timestamp 1
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_569
timestamp 1
transform -1 0 7912 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_415
timestamp 1
transform 1 0 108008 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_85
timestamp 1
transform -1 0 118864 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_250
timestamp 1
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_570
timestamp 1
transform -1 0 7912 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_416
timestamp 1
transform 1 0 108008 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_86
timestamp 1
transform -1 0 118864 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_251
timestamp 1
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_571
timestamp 1
transform -1 0 7912 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_417
timestamp 1
transform 1 0 108008 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_87
timestamp 1
transform -1 0 118864 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_252
timestamp 1
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_572
timestamp 1
transform -1 0 7912 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_418
timestamp 1
transform 1 0 108008 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_88
timestamp 1
transform -1 0 118864 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_253
timestamp 1
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_573
timestamp 1
transform -1 0 7912 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_419
timestamp 1
transform 1 0 108008 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_89
timestamp 1
transform -1 0 118864 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_254
timestamp 1
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_574
timestamp 1
transform -1 0 7912 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_420
timestamp 1
transform 1 0 108008 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_90
timestamp 1
transform -1 0 118864 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_255
timestamp 1
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_575
timestamp 1
transform -1 0 7912 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_421
timestamp 1
transform 1 0 108008 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_91
timestamp 1
transform -1 0 118864 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_256
timestamp 1
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_576
timestamp 1
transform -1 0 7912 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_422
timestamp 1
transform 1 0 108008 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_92
timestamp 1
transform -1 0 118864 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_257
timestamp 1
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_577
timestamp 1
transform -1 0 7912 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_423
timestamp 1
transform 1 0 108008 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_93
timestamp 1
transform -1 0 118864 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_258
timestamp 1
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_578
timestamp 1
transform -1 0 7912 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_424
timestamp 1
transform 1 0 108008 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_94
timestamp 1
transform -1 0 118864 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_259
timestamp 1
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_579
timestamp 1
transform -1 0 7912 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_425
timestamp 1
transform 1 0 108008 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_95
timestamp 1
transform -1 0 118864 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_260
timestamp 1
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_580
timestamp 1
transform -1 0 7912 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_426
timestamp 1
transform 1 0 108008 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_96
timestamp 1
transform -1 0 118864 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_261
timestamp 1
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_581
timestamp 1
transform -1 0 7912 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_427
timestamp 1
transform 1 0 108008 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_97
timestamp 1
transform -1 0 118864 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_262
timestamp 1
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_582
timestamp 1
transform -1 0 7912 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_428
timestamp 1
transform 1 0 108008 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_98
timestamp 1
transform -1 0 118864 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_263
timestamp 1
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_583
timestamp 1
transform -1 0 7912 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_429
timestamp 1
transform 1 0 108008 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_99
timestamp 1
transform -1 0 118864 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_264
timestamp 1
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_584
timestamp 1
transform -1 0 7912 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_430
timestamp 1
transform 1 0 108008 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_100
timestamp 1
transform -1 0 118864 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_265
timestamp 1
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_585
timestamp 1
transform -1 0 7912 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_431
timestamp 1
transform 1 0 108008 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_101
timestamp 1
transform -1 0 118864 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_266
timestamp 1
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_586
timestamp 1
transform -1 0 7912 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_432
timestamp 1
transform 1 0 108008 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_102
timestamp 1
transform -1 0 118864 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_267
timestamp 1
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_587
timestamp 1
transform -1 0 7912 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_433
timestamp 1
transform 1 0 108008 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_103
timestamp 1
transform -1 0 118864 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_268
timestamp 1
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_588
timestamp 1
transform -1 0 7912 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_434
timestamp 1
transform 1 0 108008 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_104
timestamp 1
transform -1 0 118864 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_269
timestamp 1
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_589
timestamp 1
transform -1 0 7912 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_435
timestamp 1
transform 1 0 108008 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_105
timestamp 1
transform -1 0 118864 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_270
timestamp 1
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_590
timestamp 1
transform -1 0 7912 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_436
timestamp 1
transform 1 0 108008 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_106
timestamp 1
transform -1 0 118864 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_271
timestamp 1
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_591
timestamp 1
transform -1 0 7912 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_437
timestamp 1
transform 1 0 108008 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_107
timestamp 1
transform -1 0 118864 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_272
timestamp 1
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_592
timestamp 1
transform -1 0 7912 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_438
timestamp 1
transform 1 0 108008 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_108
timestamp 1
transform -1 0 118864 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_273
timestamp 1
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_593
timestamp 1
transform -1 0 7912 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_439
timestamp 1
transform 1 0 108008 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_109
timestamp 1
transform -1 0 118864 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_274
timestamp 1
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_594
timestamp 1
transform -1 0 7912 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_440
timestamp 1
transform 1 0 108008 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_110
timestamp 1
transform -1 0 118864 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_275
timestamp 1
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_595
timestamp 1
transform -1 0 7912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_441
timestamp 1
transform 1 0 108008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_111
timestamp 1
transform -1 0 118864 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_276
timestamp 1
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_596
timestamp 1
transform -1 0 7912 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_442
timestamp 1
transform 1 0 108008 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_112
timestamp 1
transform -1 0 118864 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_277
timestamp 1
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_597
timestamp 1
transform -1 0 7912 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_443
timestamp 1
transform 1 0 108008 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_113
timestamp 1
transform -1 0 118864 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_278
timestamp 1
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_598
timestamp 1
transform -1 0 7912 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_444
timestamp 1
transform 1 0 108008 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_114
timestamp 1
transform -1 0 118864 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_279
timestamp 1
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_599
timestamp 1
transform -1 0 7912 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_445
timestamp 1
transform 1 0 108008 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_115
timestamp 1
transform -1 0 118864 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_280
timestamp 1
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_600
timestamp 1
transform -1 0 7912 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_446
timestamp 1
transform 1 0 108008 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_116
timestamp 1
transform -1 0 118864 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_281
timestamp 1
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_601
timestamp 1
transform -1 0 7912 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_447
timestamp 1
transform 1 0 108008 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_117
timestamp 1
transform -1 0 118864 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_282
timestamp 1
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_602
timestamp 1
transform -1 0 7912 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_448
timestamp 1
transform 1 0 108008 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_118
timestamp 1
transform -1 0 118864 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_283
timestamp 1
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_603
timestamp 1
transform -1 0 7912 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_449
timestamp 1
transform 1 0 108008 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_119
timestamp 1
transform -1 0 118864 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_284
timestamp 1
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_604
timestamp 1
transform -1 0 7912 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_450
timestamp 1
transform 1 0 108008 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_120
timestamp 1
transform -1 0 118864 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_285
timestamp 1
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_605
timestamp 1
transform -1 0 7912 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_451
timestamp 1
transform 1 0 108008 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_121
timestamp 1
transform -1 0 118864 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_286
timestamp 1
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_606
timestamp 1
transform -1 0 7912 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_452
timestamp 1
transform 1 0 108008 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_122
timestamp 1
transform -1 0 118864 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_287
timestamp 1
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_607
timestamp 1
transform -1 0 7912 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_453
timestamp 1
transform 1 0 108008 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_123
timestamp 1
transform -1 0 118864 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_288
timestamp 1
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_608
timestamp 1
transform -1 0 7912 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_454
timestamp 1
transform 1 0 108008 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_124
timestamp 1
transform -1 0 118864 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_289
timestamp 1
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_609
timestamp 1
transform -1 0 7912 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_455
timestamp 1
transform 1 0 108008 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_125
timestamp 1
transform -1 0 118864 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_290
timestamp 1
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_610
timestamp 1
transform -1 0 7912 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_456
timestamp 1
transform 1 0 108008 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_126
timestamp 1
transform -1 0 118864 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Left_291
timestamp 1
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Right_611
timestamp 1
transform -1 0 7912 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Left_457
timestamp 1
transform 1 0 108008 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Right_127
timestamp 1
transform -1 0 118864 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Left_292
timestamp 1
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Right_612
timestamp 1
transform -1 0 7912 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Left_458
timestamp 1
transform 1 0 108008 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Right_128
timestamp 1
transform -1 0 118864 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Left_293
timestamp 1
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Right_613
timestamp 1
transform -1 0 7912 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Left_459
timestamp 1
transform 1 0 108008 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Right_129
timestamp 1
transform -1 0 118864 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Left_294
timestamp 1
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Right_614
timestamp 1
transform -1 0 7912 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Left_460
timestamp 1
transform 1 0 108008 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Right_130
timestamp 1
transform -1 0 118864 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Left_295
timestamp 1
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Right_615
timestamp 1
transform -1 0 7912 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Left_461
timestamp 1
transform 1 0 108008 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Right_131
timestamp 1
transform -1 0 118864 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Left_296
timestamp 1
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Right_616
timestamp 1
transform -1 0 7912 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Left_462
timestamp 1
transform 1 0 108008 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Right_132
timestamp 1
transform -1 0 118864 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Left_297
timestamp 1
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Right_617
timestamp 1
transform -1 0 7912 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Left_463
timestamp 1
transform 1 0 108008 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Right_133
timestamp 1
transform -1 0 118864 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Left_298
timestamp 1
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Right_618
timestamp 1
transform -1 0 7912 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Left_464
timestamp 1
transform 1 0 108008 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Right_134
timestamp 1
transform -1 0 118864 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Left_299
timestamp 1
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Right_619
timestamp 1
transform -1 0 7912 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Left_465
timestamp 1
transform 1 0 108008 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Right_135
timestamp 1
transform -1 0 118864 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Left_300
timestamp 1
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Right_620
timestamp 1
transform -1 0 7912 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Left_466
timestamp 1
transform 1 0 108008 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Right_136
timestamp 1
transform -1 0 118864 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Left_301
timestamp 1
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Right_621
timestamp 1
transform -1 0 7912 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Left_467
timestamp 1
transform 1 0 108008 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Right_137
timestamp 1
transform -1 0 118864 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Left_302
timestamp 1
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Right_622
timestamp 1
transform -1 0 7912 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Left_468
timestamp 1
transform 1 0 108008 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Right_138
timestamp 1
transform -1 0 118864 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Left_303
timestamp 1
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Right_623
timestamp 1
transform -1 0 7912 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Left_469
timestamp 1
transform 1 0 108008 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Right_139
timestamp 1
transform -1 0 118864 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Left_304
timestamp 1
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Right_624
timestamp 1
transform -1 0 7912 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Left_470
timestamp 1
transform 1 0 108008 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Right_140
timestamp 1
transform -1 0 118864 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Left_305
timestamp 1
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Right_625
timestamp 1
transform -1 0 7912 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Left_471
timestamp 1
transform 1 0 108008 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Right_141
timestamp 1
transform -1 0 118864 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Left_306
timestamp 1
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Right_626
timestamp 1
transform -1 0 7912 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Left_472
timestamp 1
transform 1 0 108008 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Right_142
timestamp 1
transform -1 0 118864 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Left_307
timestamp 1
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Right_627
timestamp 1
transform -1 0 7912 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Left_473
timestamp 1
transform 1 0 108008 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Right_143
timestamp 1
transform -1 0 118864 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Left_308
timestamp 1
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Right_628
timestamp 1
transform -1 0 7912 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Left_474
timestamp 1
transform 1 0 108008 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Right_144
timestamp 1
transform -1 0 118864 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Left_309
timestamp 1
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Right_629
timestamp 1
transform -1 0 7912 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Left_475
timestamp 1
transform 1 0 108008 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Right_145
timestamp 1
transform -1 0 118864 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Left_310
timestamp 1
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Right_630
timestamp 1
transform -1 0 7912 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Left_476
timestamp 1
transform 1 0 108008 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Right_146
timestamp 1
transform -1 0 118864 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Left_311
timestamp 1
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Right_631
timestamp 1
transform -1 0 7912 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Left_477
timestamp 1
transform 1 0 108008 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Right_147
timestamp 1
transform -1 0 118864 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Left_312
timestamp 1
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Right_632
timestamp 1
transform -1 0 7912 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Left_478
timestamp 1
transform 1 0 108008 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Right_148
timestamp 1
transform -1 0 118864 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_313
timestamp 1
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_633
timestamp 1
transform -1 0 7912 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Left_479
timestamp 1
transform 1 0 108008 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Right_149
timestamp 1
transform -1 0 118864 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_314
timestamp 1
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_634
timestamp 1
transform -1 0 7912 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Left_480
timestamp 1
transform 1 0 108008 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Right_150
timestamp 1
transform -1 0 118864 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_315
timestamp 1
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_635
timestamp 1
transform -1 0 7912 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Left_481
timestamp 1
transform 1 0 108008 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Right_151
timestamp 1
transform -1 0 118864 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_316
timestamp 1
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_636
timestamp 1
transform -1 0 7912 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Left_482
timestamp 1
transform 1 0 108008 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Right_152
timestamp 1
transform -1 0 118864 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_317
timestamp 1
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_637
timestamp 1
transform -1 0 7912 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Left_483
timestamp 1
transform 1 0 108008 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Right_153
timestamp 1
transform -1 0 118864 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_318
timestamp 1
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_638
timestamp 1
transform -1 0 7912 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Left_484
timestamp 1
transform 1 0 108008 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Right_154
timestamp 1
transform -1 0 118864 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_319
timestamp 1
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_639
timestamp 1
transform -1 0 7912 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Left_485
timestamp 1
transform 1 0 108008 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Right_155
timestamp 1
transform -1 0 118864 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Left_320
timestamp 1
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Right_640
timestamp 1
transform -1 0 7912 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Left_486
timestamp 1
transform 1 0 108008 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Right_156
timestamp 1
transform -1 0 118864 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Left_321
timestamp 1
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Right_641
timestamp 1
transform -1 0 7912 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Left_487
timestamp 1
transform 1 0 108008 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Right_157
timestamp 1
transform -1 0 118864 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Left_322
timestamp 1
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Right_642
timestamp 1
transform -1 0 7912 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Left_488
timestamp 1
transform 1 0 108008 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Right_158
timestamp 1
transform -1 0 118864 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Left_323
timestamp 1
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Right_643
timestamp 1
transform -1 0 7912 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Left_489
timestamp 1
transform 1 0 108008 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Right_159
timestamp 1
transform -1 0 118864 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Left_324
timestamp 1
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Right_644
timestamp 1
transform -1 0 7912 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Left_490
timestamp 1
transform 1 0 108008 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Right_160
timestamp 1
transform -1 0 118864 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Left_325
timestamp 1
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Right_645
timestamp 1
transform -1 0 7912 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Left_491
timestamp 1
transform 1 0 108008 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Right_161
timestamp 1
transform -1 0 118864 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Left_326
timestamp 1
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Right_646
timestamp 1
transform -1 0 7912 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Left_492
timestamp 1
transform 1 0 108008 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Right_162
timestamp 1
transform -1 0 118864 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Left_327
timestamp 1
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Right_647
timestamp 1
transform -1 0 7912 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Left_493
timestamp 1
transform 1 0 108008 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Right_163
timestamp 1
transform -1 0 118864 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Left_328
timestamp 1
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Right_648
timestamp 1
transform -1 0 7912 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Left_494
timestamp 1
transform 1 0 108008 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Right_164
timestamp 1
transform -1 0 118864 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Left_329
timestamp 1
transform 1 0 1104 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Right_649
timestamp 1
transform -1 0 7912 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Left_495
timestamp 1
transform 1 0 108008 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Right_165
timestamp 1
transform -1 0 118864 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Left_330
timestamp 1
transform 1 0 1104 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Right_650
timestamp 1
transform -1 0 7912 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_2_Left_496
timestamp 1
transform 1 0 108008 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_2_Right_166
timestamp 1
transform -1 0 118864 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Left_331
timestamp 1
transform 1 0 1104 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Right_651
timestamp 1
transform -1 0 7912 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_2_Left_497
timestamp 1
transform 1 0 108008 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_2_Right_167
timestamp 1
transform -1 0 118864 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Left_332
timestamp 1
transform 1 0 1104 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Right_652
timestamp 1
transform -1 0 7912 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_2_Left_498
timestamp 1
transform 1 0 108008 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_2_Right_168
timestamp 1
transform -1 0 118864 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Left_333
timestamp 1
transform 1 0 1104 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Right_653
timestamp 1
transform -1 0 7912 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_2_Left_499
timestamp 1
transform 1 0 108008 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_2_Right_169
timestamp 1
transform -1 0 118864 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Left_334
timestamp 1
transform 1 0 1104 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Right_654
timestamp 1
transform -1 0 7912 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_2_Left_500
timestamp 1
transform 1 0 108008 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_2_Right_170
timestamp 1
transform -1 0 118864 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Left_335
timestamp 1
transform 1 0 1104 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Right_655
timestamp 1
transform -1 0 7912 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_2_Left_501
timestamp 1
transform 1 0 108008 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_2_Right_171
timestamp 1
transform -1 0 118864 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Left_336
timestamp 1
transform 1 0 1104 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Right_656
timestamp 1
transform -1 0 7912 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_2_Left_502
timestamp 1
transform 1 0 108008 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_2_Right_172
timestamp 1
transform -1 0 118864 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Left_337
timestamp 1
transform 1 0 1104 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Right_657
timestamp 1
transform -1 0 7912 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_2_Left_503
timestamp 1
transform 1 0 108008 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_2_Right_173
timestamp 1
transform -1 0 118864 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Left_338
timestamp 1
transform 1 0 1104 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Right_658
timestamp 1
transform -1 0 7912 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_2_Left_504
timestamp 1
transform 1 0 108008 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_2_Right_174
timestamp 1
transform -1 0 118864 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_Left_339
timestamp 1
transform 1 0 1104 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_Right_10
timestamp 1
transform -1 0 118864 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_Left_340
timestamp 1
transform 1 0 1104 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_Right_11
timestamp 1
transform -1 0 118864 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_Left_341
timestamp 1
transform 1 0 1104 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_Right_12
timestamp 1
transform -1 0 118864 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_Left_342
timestamp 1
transform 1 0 1104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_Right_13
timestamp 1
transform -1 0 118864 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_Left_343
timestamp 1
transform 1 0 1104 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_Right_14
timestamp 1
transform -1 0 118864 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_Left_344
timestamp 1
transform 1 0 1104 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_Right_15
timestamp 1
transform -1 0 118864 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_Left_345
timestamp 1
transform 1 0 1104 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_Right_16
timestamp 1
transform -1 0 118864 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_Left_346
timestamp 1
transform 1 0 1104 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_Right_17
timestamp 1
transform -1 0 118864 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_Left_347
timestamp 1
transform 1 0 1104 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_Right_18
timestamp 1
transform -1 0 118864 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_Left_348
timestamp 1
transform 1 0 1104 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_Right_19
timestamp 1
transform -1 0 118864 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 1
transform 1 0 109204 0 -1 46784
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer3
timestamp 1
transform -1 0 110400 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_660
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_661
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_662
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_663
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_664
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_665
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_666
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_667
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_668
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_669
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_670
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_671
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_672
timestamp 1
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_673
timestamp 1
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_674
timestamp 1
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_675
timestamp 1
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_676
timestamp 1
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_677
timestamp 1
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_678
timestamp 1
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_679
timestamp 1
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_680
timestamp 1
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_681
timestamp 1
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_682
timestamp 1
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_683
timestamp 1
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_684
timestamp 1
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_685
timestamp 1
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_686
timestamp 1
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_687
timestamp 1
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_688
timestamp 1
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_689
timestamp 1
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_690
timestamp 1
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_691
timestamp 1
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_692
timestamp 1
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_693
timestamp 1
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_694
timestamp 1
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_695
timestamp 1
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_696
timestamp 1
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_697
timestamp 1
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_698
timestamp 1
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_699
timestamp 1
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_700
timestamp 1
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_701
timestamp 1
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_702
timestamp 1
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_703
timestamp 1
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_704
timestamp 1
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_705
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_706
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_707
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_708
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_709
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_710
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_711
timestamp 1
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_712
timestamp 1
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_713
timestamp 1
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_714
timestamp 1
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_715
timestamp 1
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_716
timestamp 1
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_717
timestamp 1
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_718
timestamp 1
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_719
timestamp 1
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_720
timestamp 1
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_721
timestamp 1
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_722
timestamp 1
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_723
timestamp 1
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_724
timestamp 1
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_725
timestamp 1
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_726
timestamp 1
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_727
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_728
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_729
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_730
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_731
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_732
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_733
timestamp 1
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_734
timestamp 1
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_735
timestamp 1
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_736
timestamp 1
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_737
timestamp 1
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_738
timestamp 1
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_739
timestamp 1
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_740
timestamp 1
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_741
timestamp 1
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_742
timestamp 1
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_743
timestamp 1
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_744
timestamp 1
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_745
timestamp 1
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_746
timestamp 1
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_747
timestamp 1
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_748
timestamp 1
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_749
timestamp 1
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_750
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_751
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_752
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_753
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_754
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_755
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_756
timestamp 1
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_757
timestamp 1
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_758
timestamp 1
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_759
timestamp 1
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_760
timestamp 1
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_761
timestamp 1
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_762
timestamp 1
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_763
timestamp 1
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_764
timestamp 1
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_765
timestamp 1
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_766
timestamp 1
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_767
timestamp 1
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_768
timestamp 1
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_769
timestamp 1
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_770
timestamp 1
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_771
timestamp 1
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_772
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_773
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_774
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_775
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_776
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_777
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_778
timestamp 1
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_779
timestamp 1
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_780
timestamp 1
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_781
timestamp 1
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_782
timestamp 1
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_783
timestamp 1
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_784
timestamp 1
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_785
timestamp 1
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_786
timestamp 1
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_787
timestamp 1
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_788
timestamp 1
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_789
timestamp 1
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_790
timestamp 1
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_791
timestamp 1
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_792
timestamp 1
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_793
timestamp 1
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_794
timestamp 1
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_795
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_796
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_797
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_798
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_799
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_800
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_801
timestamp 1
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_802
timestamp 1
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_803
timestamp 1
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_804
timestamp 1
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_805
timestamp 1
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_806
timestamp 1
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_807
timestamp 1
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_808
timestamp 1
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_809
timestamp 1
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_810
timestamp 1
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_811
timestamp 1
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_812
timestamp 1
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_813
timestamp 1
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_814
timestamp 1
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_815
timestamp 1
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_816
timestamp 1
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_817
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_818
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_819
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_820
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_821
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_822
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_823
timestamp 1
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_824
timestamp 1
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_825
timestamp 1
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_826
timestamp 1
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_827
timestamp 1
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_828
timestamp 1
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_829
timestamp 1
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_830
timestamp 1
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_831
timestamp 1
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_832
timestamp 1
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_833
timestamp 1
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_834
timestamp 1
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_835
timestamp 1
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_836
timestamp 1
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_837
timestamp 1
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_838
timestamp 1
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_839
timestamp 1
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_840
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_841
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_842
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_843
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_844
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_845
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_846
timestamp 1
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_847
timestamp 1
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_848
timestamp 1
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_849
timestamp 1
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_850
timestamp 1
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_851
timestamp 1
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_852
timestamp 1
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_853
timestamp 1
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_854
timestamp 1
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_855
timestamp 1
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_856
timestamp 1
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_857
timestamp 1
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_858
timestamp 1
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_859
timestamp 1
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_860
timestamp 1
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_861
timestamp 1
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_862
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_863
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_864
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_865
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_866
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_867
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_868
timestamp 1
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_869
timestamp 1
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_870
timestamp 1
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_871
timestamp 1
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_872
timestamp 1
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_873
timestamp 1
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_874
timestamp 1
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_875
timestamp 1
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_876
timestamp 1
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_877
timestamp 1
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_878
timestamp 1
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_879
timestamp 1
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_880
timestamp 1
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_881
timestamp 1
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_882
timestamp 1
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_883
timestamp 1
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_884
timestamp 1
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_885
timestamp 1
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_886
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_887
timestamp 1
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_888
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_889
timestamp 1
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_890
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_891
timestamp 1
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_892
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_893
timestamp 1
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_894
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_895
timestamp 1
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_896
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_897
timestamp 1
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_898
timestamp 1
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_899
timestamp 1
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_900
timestamp 1
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_901
timestamp 1
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_902
timestamp 1
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_903
timestamp 1
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_904
timestamp 1
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_905
timestamp 1
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_906
timestamp 1
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_907
timestamp 1
transform 1 0 60352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_908
timestamp 1
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_909
timestamp 1
transform 1 0 65504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_910
timestamp 1
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_911
timestamp 1
transform 1 0 70656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_912
timestamp 1
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_913
timestamp 1
transform 1 0 75808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_914
timestamp 1
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_915
timestamp 1
transform 1 0 80960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_916
timestamp 1
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_917
timestamp 1
transform 1 0 86112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_918
timestamp 1
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_919
timestamp 1
transform 1 0 91264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_920
timestamp 1
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_921
timestamp 1
transform 1 0 96416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_922
timestamp 1
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_923
timestamp 1
transform 1 0 101568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_924
timestamp 1
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_925
timestamp 1
transform 1 0 106720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_926
timestamp 1
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_927
timestamp 1
transform 1 0 111872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_928
timestamp 1
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_929
timestamp 1
transform 1 0 117024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_1354
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_1355
timestamp 1
transform 1 0 110584 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_1356
timestamp 1
transform 1 0 115736 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_1_930
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_1357
timestamp 1
transform 1 0 113160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_1358
timestamp 1
transform 1 0 118312 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_931
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_1359
timestamp 1
transform 1 0 110584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_1360
timestamp 1
transform 1 0 115736 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_1_932
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_1361
timestamp 1
transform 1 0 113160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_1362
timestamp 1
transform 1 0 118312 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_933
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_1363
timestamp 1
transform 1 0 110584 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_1364
timestamp 1
transform 1 0 115736 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_1_934
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_2_1365
timestamp 1
transform 1 0 113160 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_2_1366
timestamp 1
transform 1 0 118312 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_935
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_1367
timestamp 1
transform 1 0 110584 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_1368
timestamp 1
transform 1 0 115736 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_1_936
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_2_1369
timestamp 1
transform 1 0 113160 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_2_1370
timestamp 1
transform 1 0 118312 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_937
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_1371
timestamp 1
transform 1 0 110584 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_1372
timestamp 1
transform 1 0 115736 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_1_938
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_2_1373
timestamp 1
transform 1 0 113160 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_2_1374
timestamp 1
transform 1 0 118312 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_939
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_1375
timestamp 1
transform 1 0 110584 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_1376
timestamp 1
transform 1 0 115736 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_1_940
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_2_1377
timestamp 1
transform 1 0 113160 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_2_1378
timestamp 1
transform 1 0 118312 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_941
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_1379
timestamp 1
transform 1 0 110584 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_1380
timestamp 1
transform 1 0 115736 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_1_942
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_2_1381
timestamp 1
transform 1 0 113160 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_2_1382
timestamp 1
transform 1 0 118312 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_943
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_1383
timestamp 1
transform 1 0 110584 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_1384
timestamp 1
transform 1 0 115736 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_1_944
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_2_1385
timestamp 1
transform 1 0 113160 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_2_1386
timestamp 1
transform 1 0 118312 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_945
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_1387
timestamp 1
transform 1 0 110584 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_1388
timestamp 1
transform 1 0 115736 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_1_946
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_2_1389
timestamp 1
transform 1 0 113160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_2_1390
timestamp 1
transform 1 0 118312 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_947
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_1391
timestamp 1
transform 1 0 110584 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_1392
timestamp 1
transform 1 0 115736 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_1_948
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_2_1393
timestamp 1
transform 1 0 113160 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_2_1394
timestamp 1
transform 1 0 118312 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_949
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_1395
timestamp 1
transform 1 0 110584 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_1396
timestamp 1
transform 1 0 115736 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_1_950
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_2_1397
timestamp 1
transform 1 0 113160 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_2_1398
timestamp 1
transform 1 0 118312 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_951
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_1399
timestamp 1
transform 1 0 110584 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_1400
timestamp 1
transform 1 0 115736 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_1_952
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_2_1401
timestamp 1
transform 1 0 113160 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_2_1402
timestamp 1
transform 1 0 118312 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_953
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_1403
timestamp 1
transform 1 0 110584 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_1404
timestamp 1
transform 1 0 115736 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_1_954
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_2_1405
timestamp 1
transform 1 0 113160 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_2_1406
timestamp 1
transform 1 0 118312 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_955
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_1407
timestamp 1
transform 1 0 110584 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_1408
timestamp 1
transform 1 0 115736 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_1_956
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_2_1409
timestamp 1
transform 1 0 113160 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_2_1410
timestamp 1
transform 1 0 118312 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_957
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_1411
timestamp 1
transform 1 0 110584 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_1412
timestamp 1
transform 1 0 115736 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_1_958
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_2_1413
timestamp 1
transform 1 0 113160 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_2_1414
timestamp 1
transform 1 0 118312 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_959
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_1415
timestamp 1
transform 1 0 110584 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_1416
timestamp 1
transform 1 0 115736 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_1_960
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_2_1417
timestamp 1
transform 1 0 113160 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_2_1418
timestamp 1
transform 1 0 118312 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_961
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_1419
timestamp 1
transform 1 0 110584 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_1420
timestamp 1
transform 1 0 115736 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_1_962
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_2_1421
timestamp 1
transform 1 0 113160 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_2_1422
timestamp 1
transform 1 0 118312 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_963
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_1423
timestamp 1
transform 1 0 110584 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_1424
timestamp 1
transform 1 0 115736 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_1_964
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_2_1425
timestamp 1
transform 1 0 113160 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_2_1426
timestamp 1
transform 1 0 118312 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_965
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_1427
timestamp 1
transform 1 0 110584 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_1428
timestamp 1
transform 1 0 115736 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_1_966
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_2_1429
timestamp 1
transform 1 0 113160 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_2_1430
timestamp 1
transform 1 0 118312 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_967
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_1431
timestamp 1
transform 1 0 110584 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_1432
timestamp 1
transform 1 0 115736 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1_968
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_2_1433
timestamp 1
transform 1 0 113160 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_2_1434
timestamp 1
transform 1 0 118312 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_969
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_1435
timestamp 1
transform 1 0 110584 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_1436
timestamp 1
transform 1 0 115736 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1_970
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_2_1437
timestamp 1
transform 1 0 113160 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_2_1438
timestamp 1
transform 1 0 118312 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_971
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_1439
timestamp 1
transform 1 0 110584 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_1440
timestamp 1
transform 1 0 115736 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1_972
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_2_1441
timestamp 1
transform 1 0 113160 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_2_1442
timestamp 1
transform 1 0 118312 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_973
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_1443
timestamp 1
transform 1 0 110584 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_1444
timestamp 1
transform 1 0 115736 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1_974
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_2_1445
timestamp 1
transform 1 0 113160 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_2_1446
timestamp 1
transform 1 0 118312 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_975
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_1447
timestamp 1
transform 1 0 110584 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_1448
timestamp 1
transform 1 0 115736 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1_976
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_2_1449
timestamp 1
transform 1 0 113160 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_2_1450
timestamp 1
transform 1 0 118312 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_977
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_1451
timestamp 1
transform 1 0 110584 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_1452
timestamp 1
transform 1 0 115736 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1_978
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_2_1453
timestamp 1
transform 1 0 113160 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_2_1454
timestamp 1
transform 1 0 118312 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_979
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_1455
timestamp 1
transform 1 0 110584 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_1456
timestamp 1
transform 1 0 115736 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1_980
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_2_1457
timestamp 1
transform 1 0 113160 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_2_1458
timestamp 1
transform 1 0 118312 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_981
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_1459
timestamp 1
transform 1 0 110584 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_1460
timestamp 1
transform 1 0 115736 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1_982
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_2_1461
timestamp 1
transform 1 0 113160 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_2_1462
timestamp 1
transform 1 0 118312 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_983
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_1463
timestamp 1
transform 1 0 110584 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_1464
timestamp 1
transform 1 0 115736 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1_984
timestamp 1
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_2_1465
timestamp 1
transform 1 0 113160 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_2_1466
timestamp 1
transform 1 0 118312 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_985
timestamp 1
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_1467
timestamp 1
transform 1 0 110584 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_1468
timestamp 1
transform 1 0 115736 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1_986
timestamp 1
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_2_1469
timestamp 1
transform 1 0 113160 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_2_1470
timestamp 1
transform 1 0 118312 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_987
timestamp 1
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_1471
timestamp 1
transform 1 0 110584 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_1472
timestamp 1
transform 1 0 115736 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1_988
timestamp 1
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_2_1473
timestamp 1
transform 1 0 113160 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_2_1474
timestamp 1
transform 1 0 118312 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_989
timestamp 1
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_1475
timestamp 1
transform 1 0 110584 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_1476
timestamp 1
transform 1 0 115736 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1_990
timestamp 1
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_2_1477
timestamp 1
transform 1 0 113160 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_2_1478
timestamp 1
transform 1 0 118312 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_991
timestamp 1
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_1479
timestamp 1
transform 1 0 110584 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_1480
timestamp 1
transform 1 0 115736 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1_992
timestamp 1
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_2_1481
timestamp 1
transform 1 0 113160 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_2_1482
timestamp 1
transform 1 0 118312 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_993
timestamp 1
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_1483
timestamp 1
transform 1 0 110584 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_1484
timestamp 1
transform 1 0 115736 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1_994
timestamp 1
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_2_1485
timestamp 1
transform 1 0 113160 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_2_1486
timestamp 1
transform 1 0 118312 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_995
timestamp 1
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_1487
timestamp 1
transform 1 0 110584 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_1488
timestamp 1
transform 1 0 115736 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1_996
timestamp 1
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_2_1489
timestamp 1
transform 1 0 113160 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_2_1490
timestamp 1
transform 1 0 118312 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_997
timestamp 1
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_1491
timestamp 1
transform 1 0 110584 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_1492
timestamp 1
transform 1 0 115736 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1_998
timestamp 1
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_2_1493
timestamp 1
transform 1 0 113160 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_2_1494
timestamp 1
transform 1 0 118312 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_999
timestamp 1
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_1495
timestamp 1
transform 1 0 110584 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_1496
timestamp 1
transform 1 0 115736 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1_1000
timestamp 1
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_2_1497
timestamp 1
transform 1 0 113160 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_2_1498
timestamp 1
transform 1 0 118312 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_1001
timestamp 1
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_1499
timestamp 1
transform 1 0 110584 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_1500
timestamp 1
transform 1 0 115736 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1_1002
timestamp 1
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_2_1501
timestamp 1
transform 1 0 113160 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_2_1502
timestamp 1
transform 1 0 118312 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_1003
timestamp 1
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_1503
timestamp 1
transform 1 0 110584 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_1504
timestamp 1
transform 1 0 115736 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1_1004
timestamp 1
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_2_1505
timestamp 1
transform 1 0 113160 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_2_1506
timestamp 1
transform 1 0 118312 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_1005
timestamp 1
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_1507
timestamp 1
transform 1 0 110584 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_1508
timestamp 1
transform 1 0 115736 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1_1006
timestamp 1
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_2_1509
timestamp 1
transform 1 0 113160 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_2_1510
timestamp 1
transform 1 0 118312 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_1007
timestamp 1
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_1511
timestamp 1
transform 1 0 110584 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_1512
timestamp 1
transform 1 0 115736 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1_1008
timestamp 1
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_2_1513
timestamp 1
transform 1 0 113160 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_2_1514
timestamp 1
transform 1 0 118312 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_1009
timestamp 1
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_1515
timestamp 1
transform 1 0 110584 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_1516
timestamp 1
transform 1 0 115736 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1_1010
timestamp 1
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_2_1517
timestamp 1
transform 1 0 113160 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_2_1518
timestamp 1
transform 1 0 118312 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_1011
timestamp 1
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_1519
timestamp 1
transform 1 0 110584 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_1520
timestamp 1
transform 1 0 115736 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1_1012
timestamp 1
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_2_1521
timestamp 1
transform 1 0 113160 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_2_1522
timestamp 1
transform 1 0 118312 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_1013
timestamp 1
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_1523
timestamp 1
transform 1 0 110584 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_1524
timestamp 1
transform 1 0 115736 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1_1014
timestamp 1
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_2_1525
timestamp 1
transform 1 0 113160 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_2_1526
timestamp 1
transform 1 0 118312 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_1015
timestamp 1
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_1527
timestamp 1
transform 1 0 110584 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_1528
timestamp 1
transform 1 0 115736 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1_1016
timestamp 1
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_2_1529
timestamp 1
transform 1 0 113160 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_2_1530
timestamp 1
transform 1 0 118312 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_1017
timestamp 1
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_1531
timestamp 1
transform 1 0 110584 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_1532
timestamp 1
transform 1 0 115736 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1_1018
timestamp 1
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_2_1533
timestamp 1
transform 1 0 113160 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_2_1534
timestamp 1
transform 1 0 118312 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_1019
timestamp 1
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_1535
timestamp 1
transform 1 0 110584 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_1536
timestamp 1
transform 1 0 115736 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1_1020
timestamp 1
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_2_1537
timestamp 1
transform 1 0 113160 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_2_1538
timestamp 1
transform 1 0 118312 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_1021
timestamp 1
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_1539
timestamp 1
transform 1 0 110584 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_1540
timestamp 1
transform 1 0 115736 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1_1022
timestamp 1
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_2_1541
timestamp 1
transform 1 0 113160 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_2_1542
timestamp 1
transform 1 0 118312 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_1023
timestamp 1
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_1543
timestamp 1
transform 1 0 110584 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_1544
timestamp 1
transform 1 0 115736 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1_1024
timestamp 1
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_2_1545
timestamp 1
transform 1 0 113160 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_2_1546
timestamp 1
transform 1 0 118312 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_1025
timestamp 1
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_1547
timestamp 1
transform 1 0 110584 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_1548
timestamp 1
transform 1 0 115736 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1_1026
timestamp 1
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_2_1549
timestamp 1
transform 1 0 113160 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_2_1550
timestamp 1
transform 1 0 118312 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_1027
timestamp 1
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_1551
timestamp 1
transform 1 0 110584 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_1552
timestamp 1
transform 1 0 115736 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1_1028
timestamp 1
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_2_1553
timestamp 1
transform 1 0 113160 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_2_1554
timestamp 1
transform 1 0 118312 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_1029
timestamp 1
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_1555
timestamp 1
transform 1 0 110584 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_1556
timestamp 1
transform 1 0 115736 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1_1030
timestamp 1
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_2_1557
timestamp 1
transform 1 0 113160 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_2_1558
timestamp 1
transform 1 0 118312 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_1031
timestamp 1
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_1559
timestamp 1
transform 1 0 110584 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_1560
timestamp 1
transform 1 0 115736 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1_1032
timestamp 1
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_2_1561
timestamp 1
transform 1 0 113160 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_2_1562
timestamp 1
transform 1 0 118312 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_1033
timestamp 1
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_1563
timestamp 1
transform 1 0 110584 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_1564
timestamp 1
transform 1 0 115736 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1_1034
timestamp 1
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_2_1565
timestamp 1
transform 1 0 113160 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_2_1566
timestamp 1
transform 1 0 118312 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_1035
timestamp 1
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_1567
timestamp 1
transform 1 0 110584 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_1568
timestamp 1
transform 1 0 115736 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1_1036
timestamp 1
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2_1569
timestamp 1
transform 1 0 113160 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2_1570
timestamp 1
transform 1 0 118312 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1_1037
timestamp 1
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_1571
timestamp 1
transform 1 0 110584 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_1572
timestamp 1
transform 1 0 115736 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1_1038
timestamp 1
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2_1573
timestamp 1
transform 1 0 113160 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2_1574
timestamp 1
transform 1 0 118312 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1_1039
timestamp 1
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_1575
timestamp 1
transform 1 0 110584 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_1576
timestamp 1
transform 1 0 115736 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1_1040
timestamp 1
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2_1577
timestamp 1
transform 1 0 113160 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2_1578
timestamp 1
transform 1 0 118312 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1_1041
timestamp 1
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_1579
timestamp 1
transform 1 0 110584 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_1580
timestamp 1
transform 1 0 115736 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1_1042
timestamp 1
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2_1581
timestamp 1
transform 1 0 113160 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2_1582
timestamp 1
transform 1 0 118312 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1_1043
timestamp 1
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_1583
timestamp 1
transform 1 0 110584 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_1584
timestamp 1
transform 1 0 115736 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1_1044
timestamp 1
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2_1585
timestamp 1
transform 1 0 113160 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2_1586
timestamp 1
transform 1 0 118312 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1_1045
timestamp 1
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_1587
timestamp 1
transform 1 0 110584 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_1588
timestamp 1
transform 1 0 115736 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1_1046
timestamp 1
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2_1589
timestamp 1
transform 1 0 113160 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2_1590
timestamp 1
transform 1 0 118312 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1_1047
timestamp 1
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_1591
timestamp 1
transform 1 0 110584 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_1592
timestamp 1
transform 1 0 115736 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1_1048
timestamp 1
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2_1593
timestamp 1
transform 1 0 113160 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2_1594
timestamp 1
transform 1 0 118312 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1_1049
timestamp 1
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_1595
timestamp 1
transform 1 0 110584 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_1596
timestamp 1
transform 1 0 115736 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1_1050
timestamp 1
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2_1597
timestamp 1
transform 1 0 113160 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2_1598
timestamp 1
transform 1 0 118312 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1_1051
timestamp 1
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_1599
timestamp 1
transform 1 0 110584 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_1600
timestamp 1
transform 1 0 115736 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1_1052
timestamp 1
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2_1601
timestamp 1
transform 1 0 113160 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2_1602
timestamp 1
transform 1 0 118312 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1_1053
timestamp 1
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_1603
timestamp 1
transform 1 0 110584 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_1604
timestamp 1
transform 1 0 115736 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1_1054
timestamp 1
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2_1605
timestamp 1
transform 1 0 113160 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2_1606
timestamp 1
transform 1 0 118312 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1_1055
timestamp 1
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_1607
timestamp 1
transform 1 0 110584 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_1608
timestamp 1
transform 1 0 115736 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1_1056
timestamp 1
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2_1609
timestamp 1
transform 1 0 113160 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2_1610
timestamp 1
transform 1 0 118312 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1_1057
timestamp 1
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_1611
timestamp 1
transform 1 0 110584 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_1612
timestamp 1
transform 1 0 115736 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1_1058
timestamp 1
transform 1 0 6256 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_2_1613
timestamp 1
transform 1 0 113160 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_2_1614
timestamp 1
transform 1 0 118312 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_1059
timestamp 1
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_1615
timestamp 1
transform 1 0 110584 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_1616
timestamp 1
transform 1 0 115736 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1_1060
timestamp 1
transform 1 0 6256 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_2_1617
timestamp 1
transform 1 0 113160 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_2_1618
timestamp 1
transform 1 0 118312 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_1061
timestamp 1
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_1619
timestamp 1
transform 1 0 110584 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_1620
timestamp 1
transform 1 0 115736 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1_1062
timestamp 1
transform 1 0 6256 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_2_1621
timestamp 1
transform 1 0 113160 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_2_1622
timestamp 1
transform 1 0 118312 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_1063
timestamp 1
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_1623
timestamp 1
transform 1 0 110584 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_1624
timestamp 1
transform 1 0 115736 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1_1064
timestamp 1
transform 1 0 6256 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_2_1625
timestamp 1
transform 1 0 113160 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_2_1626
timestamp 1
transform 1 0 118312 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1_1065
timestamp 1
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_1627
timestamp 1
transform 1 0 110584 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_1628
timestamp 1
transform 1 0 115736 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1_1066
timestamp 1
transform 1 0 6256 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_2_1629
timestamp 1
transform 1 0 113160 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_2_1630
timestamp 1
transform 1 0 118312 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1_1067
timestamp 1
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_1631
timestamp 1
transform 1 0 110584 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_1632
timestamp 1
transform 1 0 115736 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1_1068
timestamp 1
transform 1 0 6256 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_2_1633
timestamp 1
transform 1 0 113160 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_2_1634
timestamp 1
transform 1 0 118312 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1_1069
timestamp 1
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_1635
timestamp 1
transform 1 0 110584 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_1636
timestamp 1
transform 1 0 115736 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1_1070
timestamp 1
transform 1 0 6256 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_2_1637
timestamp 1
transform 1 0 113160 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_2_1638
timestamp 1
transform 1 0 118312 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1_1071
timestamp 1
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_1639
timestamp 1
transform 1 0 110584 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_1640
timestamp 1
transform 1 0 115736 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1_1072
timestamp 1
transform 1 0 6256 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_2_1641
timestamp 1
transform 1 0 113160 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_2_1642
timestamp 1
transform 1 0 118312 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1_1073
timestamp 1
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_1643
timestamp 1
transform 1 0 110584 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_1644
timestamp 1
transform 1 0 115736 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1_1074
timestamp 1
transform 1 0 6256 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_1645
timestamp 1
transform 1 0 113160 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_1646
timestamp 1
transform 1 0 118312 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1_1075
timestamp 1
transform 1 0 3680 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_2_1647
timestamp 1
transform 1 0 110584 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_2_1648
timestamp 1
transform 1 0 115736 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1_1076
timestamp 1
transform 1 0 6256 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_2_1649
timestamp 1
transform 1 0 113160 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_2_1650
timestamp 1
transform 1 0 118312 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1_1077
timestamp 1
transform 1 0 3680 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_2_1651
timestamp 1
transform 1 0 110584 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_2_1652
timestamp 1
transform 1 0 115736 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1_1078
timestamp 1
transform 1 0 6256 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_2_1653
timestamp 1
transform 1 0 113160 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_2_1654
timestamp 1
transform 1 0 118312 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1_1079
timestamp 1
transform 1 0 3680 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_2_1655
timestamp 1
transform 1 0 110584 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_2_1656
timestamp 1
transform 1 0 115736 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1_1080
timestamp 1
transform 1 0 6256 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_2_1657
timestamp 1
transform 1 0 113160 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_2_1658
timestamp 1
transform 1 0 118312 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1_1081
timestamp 1
transform 1 0 3680 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_2_1659
timestamp 1
transform 1 0 110584 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_2_1660
timestamp 1
transform 1 0 115736 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1_1082
timestamp 1
transform 1 0 6256 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_2_1661
timestamp 1
transform 1 0 113160 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_2_1662
timestamp 1
transform 1 0 118312 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1_1083
timestamp 1
transform 1 0 3680 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_2_1663
timestamp 1
transform 1 0 110584 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_2_1664
timestamp 1
transform 1 0 115736 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1084
timestamp 1
transform 1 0 3680 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1085
timestamp 1
transform 1 0 6256 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1086
timestamp 1
transform 1 0 8832 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1087
timestamp 1
transform 1 0 11408 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1088
timestamp 1
transform 1 0 13984 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1089
timestamp 1
transform 1 0 16560 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1090
timestamp 1
transform 1 0 19136 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1091
timestamp 1
transform 1 0 21712 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1092
timestamp 1
transform 1 0 24288 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1093
timestamp 1
transform 1 0 26864 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1094
timestamp 1
transform 1 0 29440 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1095
timestamp 1
transform 1 0 32016 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1096
timestamp 1
transform 1 0 34592 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1097
timestamp 1
transform 1 0 37168 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1098
timestamp 1
transform 1 0 39744 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1099
timestamp 1
transform 1 0 42320 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1100
timestamp 1
transform 1 0 44896 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1101
timestamp 1
transform 1 0 47472 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1102
timestamp 1
transform 1 0 50048 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1103
timestamp 1
transform 1 0 52624 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1104
timestamp 1
transform 1 0 55200 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1105
timestamp 1
transform 1 0 57776 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1106
timestamp 1
transform 1 0 60352 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1107
timestamp 1
transform 1 0 62928 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1108
timestamp 1
transform 1 0 65504 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1109
timestamp 1
transform 1 0 68080 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1110
timestamp 1
transform 1 0 70656 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1111
timestamp 1
transform 1 0 73232 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1112
timestamp 1
transform 1 0 75808 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1113
timestamp 1
transform 1 0 78384 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1114
timestamp 1
transform 1 0 80960 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1115
timestamp 1
transform 1 0 83536 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1116
timestamp 1
transform 1 0 86112 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1117
timestamp 1
transform 1 0 88688 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1118
timestamp 1
transform 1 0 91264 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1119
timestamp 1
transform 1 0 93840 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1120
timestamp 1
transform 1 0 96416 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1121
timestamp 1
transform 1 0 98992 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1122
timestamp 1
transform 1 0 101568 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1123
timestamp 1
transform 1 0 104144 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1124
timestamp 1
transform 1 0 106720 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1125
timestamp 1
transform 1 0 109296 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1126
timestamp 1
transform 1 0 111872 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1127
timestamp 1
transform 1 0 114448 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1128
timestamp 1
transform 1 0 117024 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1129
timestamp 1
transform 1 0 3680 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1130
timestamp 1
transform 1 0 8832 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1131
timestamp 1
transform 1 0 13984 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1132
timestamp 1
transform 1 0 19136 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1133
timestamp 1
transform 1 0 24288 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1134
timestamp 1
transform 1 0 29440 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1135
timestamp 1
transform 1 0 34592 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1136
timestamp 1
transform 1 0 39744 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1137
timestamp 1
transform 1 0 44896 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1138
timestamp 1
transform 1 0 50048 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1139
timestamp 1
transform 1 0 55200 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1140
timestamp 1
transform 1 0 60352 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1141
timestamp 1
transform 1 0 65504 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1142
timestamp 1
transform 1 0 70656 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1143
timestamp 1
transform 1 0 75808 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1144
timestamp 1
transform 1 0 80960 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1145
timestamp 1
transform 1 0 86112 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1146
timestamp 1
transform 1 0 91264 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1147
timestamp 1
transform 1 0 96416 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1148
timestamp 1
transform 1 0 101568 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1149
timestamp 1
transform 1 0 106720 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1150
timestamp 1
transform 1 0 111872 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1151
timestamp 1
transform 1 0 117024 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1152
timestamp 1
transform 1 0 6256 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1153
timestamp 1
transform 1 0 11408 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1154
timestamp 1
transform 1 0 16560 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1155
timestamp 1
transform 1 0 21712 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1156
timestamp 1
transform 1 0 26864 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1157
timestamp 1
transform 1 0 32016 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1158
timestamp 1
transform 1 0 37168 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1159
timestamp 1
transform 1 0 42320 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1160
timestamp 1
transform 1 0 47472 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1161
timestamp 1
transform 1 0 52624 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1162
timestamp 1
transform 1 0 57776 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1163
timestamp 1
transform 1 0 62928 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1164
timestamp 1
transform 1 0 68080 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1165
timestamp 1
transform 1 0 73232 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1166
timestamp 1
transform 1 0 78384 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1167
timestamp 1
transform 1 0 83536 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1168
timestamp 1
transform 1 0 88688 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1169
timestamp 1
transform 1 0 93840 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1170
timestamp 1
transform 1 0 98992 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1171
timestamp 1
transform 1 0 104144 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1172
timestamp 1
transform 1 0 109296 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1173
timestamp 1
transform 1 0 114448 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1174
timestamp 1
transform 1 0 3680 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1175
timestamp 1
transform 1 0 8832 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1176
timestamp 1
transform 1 0 13984 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1177
timestamp 1
transform 1 0 19136 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1178
timestamp 1
transform 1 0 24288 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1179
timestamp 1
transform 1 0 29440 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1180
timestamp 1
transform 1 0 34592 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1181
timestamp 1
transform 1 0 39744 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1182
timestamp 1
transform 1 0 44896 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1183
timestamp 1
transform 1 0 50048 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1184
timestamp 1
transform 1 0 55200 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1185
timestamp 1
transform 1 0 60352 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1186
timestamp 1
transform 1 0 65504 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1187
timestamp 1
transform 1 0 70656 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1188
timestamp 1
transform 1 0 75808 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1189
timestamp 1
transform 1 0 80960 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1190
timestamp 1
transform 1 0 86112 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1191
timestamp 1
transform 1 0 91264 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1192
timestamp 1
transform 1 0 96416 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1193
timestamp 1
transform 1 0 101568 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1194
timestamp 1
transform 1 0 106720 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1195
timestamp 1
transform 1 0 111872 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1196
timestamp 1
transform 1 0 117024 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1197
timestamp 1
transform 1 0 6256 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1198
timestamp 1
transform 1 0 11408 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1199
timestamp 1
transform 1 0 16560 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1200
timestamp 1
transform 1 0 21712 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1201
timestamp 1
transform 1 0 26864 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1202
timestamp 1
transform 1 0 32016 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1203
timestamp 1
transform 1 0 37168 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1204
timestamp 1
transform 1 0 42320 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1205
timestamp 1
transform 1 0 47472 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1206
timestamp 1
transform 1 0 52624 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1207
timestamp 1
transform 1 0 57776 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1208
timestamp 1
transform 1 0 62928 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1209
timestamp 1
transform 1 0 68080 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1210
timestamp 1
transform 1 0 73232 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1211
timestamp 1
transform 1 0 78384 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1212
timestamp 1
transform 1 0 83536 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1213
timestamp 1
transform 1 0 88688 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1214
timestamp 1
transform 1 0 93840 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1215
timestamp 1
transform 1 0 98992 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1216
timestamp 1
transform 1 0 104144 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1217
timestamp 1
transform 1 0 109296 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1218
timestamp 1
transform 1 0 114448 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1219
timestamp 1
transform 1 0 3680 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1220
timestamp 1
transform 1 0 8832 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1221
timestamp 1
transform 1 0 13984 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1222
timestamp 1
transform 1 0 19136 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1223
timestamp 1
transform 1 0 24288 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1224
timestamp 1
transform 1 0 29440 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1225
timestamp 1
transform 1 0 34592 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1226
timestamp 1
transform 1 0 39744 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1227
timestamp 1
transform 1 0 44896 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1228
timestamp 1
transform 1 0 50048 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1229
timestamp 1
transform 1 0 55200 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1230
timestamp 1
transform 1 0 60352 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1231
timestamp 1
transform 1 0 65504 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1232
timestamp 1
transform 1 0 70656 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1233
timestamp 1
transform 1 0 75808 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1234
timestamp 1
transform 1 0 80960 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1235
timestamp 1
transform 1 0 86112 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1236
timestamp 1
transform 1 0 91264 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1237
timestamp 1
transform 1 0 96416 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1238
timestamp 1
transform 1 0 101568 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1239
timestamp 1
transform 1 0 106720 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1240
timestamp 1
transform 1 0 111872 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1241
timestamp 1
transform 1 0 117024 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1242
timestamp 1
transform 1 0 6256 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1243
timestamp 1
transform 1 0 11408 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1244
timestamp 1
transform 1 0 16560 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1245
timestamp 1
transform 1 0 21712 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1246
timestamp 1
transform 1 0 26864 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1247
timestamp 1
transform 1 0 32016 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1248
timestamp 1
transform 1 0 37168 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1249
timestamp 1
transform 1 0 42320 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1250
timestamp 1
transform 1 0 47472 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1251
timestamp 1
transform 1 0 52624 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1252
timestamp 1
transform 1 0 57776 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1253
timestamp 1
transform 1 0 62928 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1254
timestamp 1
transform 1 0 68080 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1255
timestamp 1
transform 1 0 73232 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1256
timestamp 1
transform 1 0 78384 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1257
timestamp 1
transform 1 0 83536 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1258
timestamp 1
transform 1 0 88688 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1259
timestamp 1
transform 1 0 93840 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1260
timestamp 1
transform 1 0 98992 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1261
timestamp 1
transform 1 0 104144 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1262
timestamp 1
transform 1 0 109296 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1263
timestamp 1
transform 1 0 114448 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1264
timestamp 1
transform 1 0 3680 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1265
timestamp 1
transform 1 0 8832 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1266
timestamp 1
transform 1 0 13984 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1267
timestamp 1
transform 1 0 19136 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1268
timestamp 1
transform 1 0 24288 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1269
timestamp 1
transform 1 0 29440 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1270
timestamp 1
transform 1 0 34592 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1271
timestamp 1
transform 1 0 39744 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1272
timestamp 1
transform 1 0 44896 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1273
timestamp 1
transform 1 0 50048 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1274
timestamp 1
transform 1 0 55200 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1275
timestamp 1
transform 1 0 60352 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1276
timestamp 1
transform 1 0 65504 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1277
timestamp 1
transform 1 0 70656 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1278
timestamp 1
transform 1 0 75808 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1279
timestamp 1
transform 1 0 80960 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1280
timestamp 1
transform 1 0 86112 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1281
timestamp 1
transform 1 0 91264 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1282
timestamp 1
transform 1 0 96416 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1283
timestamp 1
transform 1 0 101568 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1284
timestamp 1
transform 1 0 106720 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1285
timestamp 1
transform 1 0 111872 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1286
timestamp 1
transform 1 0 117024 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1287
timestamp 1
transform 1 0 6256 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1288
timestamp 1
transform 1 0 11408 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1289
timestamp 1
transform 1 0 16560 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1290
timestamp 1
transform 1 0 21712 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1291
timestamp 1
transform 1 0 26864 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1292
timestamp 1
transform 1 0 32016 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1293
timestamp 1
transform 1 0 37168 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1294
timestamp 1
transform 1 0 42320 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1295
timestamp 1
transform 1 0 47472 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1296
timestamp 1
transform 1 0 52624 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1297
timestamp 1
transform 1 0 57776 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1298
timestamp 1
transform 1 0 62928 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1299
timestamp 1
transform 1 0 68080 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1300
timestamp 1
transform 1 0 73232 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1301
timestamp 1
transform 1 0 78384 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1302
timestamp 1
transform 1 0 83536 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1303
timestamp 1
transform 1 0 88688 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1304
timestamp 1
transform 1 0 93840 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1305
timestamp 1
transform 1 0 98992 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1306
timestamp 1
transform 1 0 104144 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1307
timestamp 1
transform 1 0 109296 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1308
timestamp 1
transform 1 0 114448 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1309
timestamp 1
transform 1 0 3680 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1310
timestamp 1
transform 1 0 6256 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1311
timestamp 1
transform 1 0 8832 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1312
timestamp 1
transform 1 0 11408 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1313
timestamp 1
transform 1 0 13984 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1314
timestamp 1
transform 1 0 16560 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1315
timestamp 1
transform 1 0 19136 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1316
timestamp 1
transform 1 0 21712 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1317
timestamp 1
transform 1 0 24288 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1318
timestamp 1
transform 1 0 26864 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1319
timestamp 1
transform 1 0 29440 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1320
timestamp 1
transform 1 0 32016 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1321
timestamp 1
transform 1 0 34592 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1322
timestamp 1
transform 1 0 37168 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1323
timestamp 1
transform 1 0 39744 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1324
timestamp 1
transform 1 0 42320 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1325
timestamp 1
transform 1 0 44896 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1326
timestamp 1
transform 1 0 47472 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1327
timestamp 1
transform 1 0 50048 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1328
timestamp 1
transform 1 0 52624 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1329
timestamp 1
transform 1 0 55200 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1330
timestamp 1
transform 1 0 57776 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1331
timestamp 1
transform 1 0 60352 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1332
timestamp 1
transform 1 0 62928 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1333
timestamp 1
transform 1 0 65504 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1334
timestamp 1
transform 1 0 68080 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1335
timestamp 1
transform 1 0 70656 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1336
timestamp 1
transform 1 0 73232 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1337
timestamp 1
transform 1 0 75808 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1338
timestamp 1
transform 1 0 78384 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1339
timestamp 1
transform 1 0 80960 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1340
timestamp 1
transform 1 0 83536 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1341
timestamp 1
transform 1 0 86112 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1342
timestamp 1
transform 1 0 88688 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1343
timestamp 1
transform 1 0 91264 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1344
timestamp 1
transform 1 0 93840 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1345
timestamp 1
transform 1 0 96416 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1346
timestamp 1
transform 1 0 98992 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1347
timestamp 1
transform 1 0 101568 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1348
timestamp 1
transform 1 0 104144 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1349
timestamp 1
transform 1 0 106720 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1350
timestamp 1
transform 1 0 109296 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1351
timestamp 1
transform 1 0 111872 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1352
timestamp 1
transform 1 0 114448 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1353
timestamp 1
transform 1 0 117024 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire73
timestamp 1
transform -1 0 111872 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  wire74
timestamp 1
transform 1 0 112332 0 1 30464
box -38 -48 406 592
<< labels >>
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 addr00[0]
port 0 nsew signal input
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 addr00[1]
port 1 nsew signal input
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 addr00[2]
port 2 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 addr00[3]
port 3 nsew signal input
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 addr00[4]
port 4 nsew signal input
flabel metal3 s 0 40808 800 40928 0 FreeSans 480 0 0 0 addr00[5]
port 5 nsew signal input
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 addr00[6]
port 6 nsew signal input
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 addr00[7]
port 7 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 addr01[0]
port 8 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 addr01[1]
port 9 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 addr01[2]
port 10 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 addr01[3]
port 11 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 addr01[4]
port 12 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 addr01[5]
port 13 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 addr01[6]
port 14 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 addr01[7]
port 15 nsew signal input
flabel metal2 s 108210 99200 108266 100000 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 csb00
port 17 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 csb01
port 18 nsew signal input
flabel metal3 s 119200 28568 120000 28688 0 FreeSans 480 0 0 0 denum[0]
port 19 nsew signal input
flabel metal3 s 119200 27888 120000 28008 0 FreeSans 480 0 0 0 denum[1]
port 20 nsew signal input
flabel metal3 s 119200 29928 120000 30048 0 FreeSans 480 0 0 0 denum[2]
port 21 nsew signal input
flabel metal3 s 119200 29248 120000 29368 0 FreeSans 480 0 0 0 denum[3]
port 22 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 din00[0]
port 23 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 din00[10]
port 24 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 din00[11]
port 25 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 din00[12]
port 26 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 din00[13]
port 27 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 din00[14]
port 28 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 din00[15]
port 29 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 din00[1]
port 30 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 din00[2]
port 31 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 din00[3]
port 32 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 din00[4]
port 33 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 din00[5]
port 34 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 din00[6]
port 35 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 din00[7]
port 36 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 din00[8]
port 37 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 din00[9]
port 38 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 din01[0]
port 39 nsew signal input
flabel metal2 s 61842 0 61898 800 0 FreeSans 224 90 0 0 din01[10]
port 40 nsew signal input
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 din01[11]
port 41 nsew signal input
flabel metal2 s 63774 0 63830 800 0 FreeSans 224 90 0 0 din01[12]
port 42 nsew signal input
flabel metal2 s 65062 0 65118 800 0 FreeSans 224 90 0 0 din01[13]
port 43 nsew signal input
flabel metal2 s 66350 0 66406 800 0 FreeSans 224 90 0 0 din01[14]
port 44 nsew signal input
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 din01[15]
port 45 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 din01[1]
port 46 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 din01[2]
port 47 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 din01[3]
port 48 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 din01[4]
port 49 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 din01[5]
port 50 nsew signal input
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 din01[6]
port 51 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 din01[7]
port 52 nsew signal input
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 din01[8]
port 53 nsew signal input
flabel metal2 s 60554 0 60610 800 0 FreeSans 224 90 0 0 din01[9]
port 54 nsew signal input
flabel metal3 s 119200 30608 120000 30728 0 FreeSans 480 0 0 0 num[0]
port 55 nsew signal input
flabel metal3 s 119200 31968 120000 32088 0 FreeSans 480 0 0 0 num[1]
port 56 nsew signal input
flabel metal3 s 119200 27208 120000 27328 0 FreeSans 480 0 0 0 num[2]
port 57 nsew signal input
flabel metal3 s 119200 31288 120000 31408 0 FreeSans 480 0 0 0 num[3]
port 58 nsew signal input
flabel metal2 s 107566 99200 107622 100000 0 FreeSans 224 90 0 0 rst
port 59 nsew signal input
flabel metal2 s 56046 99200 56102 100000 0 FreeSans 224 90 0 0 sine_out[0]
port 60 nsew signal output
flabel metal2 s 67638 99200 67694 100000 0 FreeSans 224 90 0 0 sine_out[10]
port 61 nsew signal output
flabel metal2 s 68926 99200 68982 100000 0 FreeSans 224 90 0 0 sine_out[11]
port 62 nsew signal output
flabel metal2 s 70214 99200 70270 100000 0 FreeSans 224 90 0 0 sine_out[12]
port 63 nsew signal output
flabel metal2 s 71502 99200 71558 100000 0 FreeSans 224 90 0 0 sine_out[13]
port 64 nsew signal output
flabel metal2 s 72146 99200 72202 100000 0 FreeSans 224 90 0 0 sine_out[14]
port 65 nsew signal output
flabel metal2 s 74078 99200 74134 100000 0 FreeSans 224 90 0 0 sine_out[15]
port 66 nsew signal output
flabel metal2 s 57334 99200 57390 100000 0 FreeSans 224 90 0 0 sine_out[1]
port 67 nsew signal output
flabel metal2 s 58622 99200 58678 100000 0 FreeSans 224 90 0 0 sine_out[2]
port 68 nsew signal output
flabel metal2 s 60554 99200 60610 100000 0 FreeSans 224 90 0 0 sine_out[3]
port 69 nsew signal output
flabel metal2 s 59910 99200 59966 100000 0 FreeSans 224 90 0 0 sine_out[4]
port 70 nsew signal output
flabel metal2 s 62486 99200 62542 100000 0 FreeSans 224 90 0 0 sine_out[5]
port 71 nsew signal output
flabel metal2 s 63130 99200 63186 100000 0 FreeSans 224 90 0 0 sine_out[6]
port 72 nsew signal output
flabel metal2 s 64418 99200 64474 100000 0 FreeSans 224 90 0 0 sine_out[7]
port 73 nsew signal output
flabel metal2 s 65062 99200 65118 100000 0 FreeSans 224 90 0 0 sine_out[8]
port 74 nsew signal output
flabel metal2 s 66994 99200 67050 100000 0 FreeSans 224 90 0 0 sine_out[9]
port 75 nsew signal output
flabel metal4 s 4208 2128 4528 97424 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 34928 2128 35248 7880 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 34928 91436 35248 97424 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 65648 2128 65968 7880 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 65648 91620 65968 97424 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 96368 2128 96688 8064 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 96368 91436 96688 97424 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 1056 5346 118912 5666 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 1056 35982 118912 36302 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 1056 66618 118912 66938 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 112908 7024 113228 92528 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 4208 94020 118912 94340 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 4868 2128 5188 97424 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 8064 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 35588 91436 35908 97424 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 66308 2128 66628 7880 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 66308 91436 66628 97424 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 97028 2128 97348 8064 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 97028 91436 97348 97424 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 1056 6006 118912 6326 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 1056 36642 118912 36962 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 1056 67278 118912 67598 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 113644 7024 113964 92528 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 4208 94700 118912 95020 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
rlabel via4 104830 66778 104830 66778 0 vccd1
rlabel via4 105510 67438 105510 67438 0 vssd1
rlabel metal1 55246 95574 55246 95574 0 _000_
rlabel metal1 65090 93704 65090 93704 0 _001_
rlabel metal1 66792 94010 66792 94010 0 _002_
rlabel metal1 67436 93194 67436 93194 0 _003_
rlabel metal1 69000 93126 69000 93126 0 _004_
rlabel metal2 69782 93976 69782 93976 0 _005_
rlabel metal1 71346 93126 71346 93126 0 _006_
rlabel metal1 56212 94554 56212 94554 0 _007_
rlabel metal1 58190 94792 58190 94792 0 _008_
rlabel metal1 57730 95506 57730 95506 0 _009_
rlabel metal1 59340 94350 59340 94350 0 _010_
rlabel metal2 60766 94690 60766 94690 0 _011_
rlabel metal1 61226 93704 61226 93704 0 _012_
rlabel metal1 62284 93670 62284 93670 0 _013_
rlabel metal1 63296 93670 63296 93670 0 _014_
rlabel metal2 64170 94384 64170 94384 0 _015_
rlabel metal1 108790 49402 108790 49402 0 _016_
rlabel metal1 109066 45356 109066 45356 0 _017_
rlabel metal1 110308 45866 110308 45866 0 _018_
rlabel metal1 110124 40698 110124 40698 0 _019_
rlabel metal2 108606 39202 108606 39202 0 _020_
rlabel metal1 109250 35768 109250 35768 0 _021_
rlabel metal1 109618 36346 109618 36346 0 _022_
rlabel metal1 109802 37434 109802 37434 0 _023_
rlabel metal1 109894 43962 109894 43962 0 _024_
rlabel metal1 58558 94486 58558 94486 0 _025_
rlabel metal1 58749 95914 58749 95914 0 _026_
rlabel metal2 61778 94690 61778 94690 0 _027_
rlabel metal1 62974 93806 62974 93806 0 _028_
rlabel metal2 63250 93908 63250 93908 0 _029_
rlabel metal1 65090 93806 65090 93806 0 _030_
rlabel metal1 65320 94554 65320 94554 0 _031_
rlabel metal1 66654 93670 66654 93670 0 _032_
rlabel metal2 67114 94690 67114 94690 0 _033_
rlabel metal1 67942 93670 67942 93670 0 _034_
rlabel metal2 69138 94860 69138 94860 0 _035_
rlabel metal1 69414 94010 69414 94010 0 _036_
rlabel metal2 70886 93568 70886 93568 0 _037_
rlabel metal1 72220 93466 72220 93466 0 _038_
rlabel metal2 73002 94146 73002 94146 0 _039_
rlabel metal2 74750 94690 74750 94690 0 _040_
rlabel metal1 108790 54570 108790 54570 0 _041_
rlabel metal2 108974 49402 108974 49402 0 _042_
rlabel metal1 108744 49130 108744 49130 0 _043_
rlabel metal2 108560 43860 108560 43860 0 _044_
rlabel metal1 108652 44234 108652 44234 0 _045_
rlabel metal1 108507 36822 108507 36822 0 _046_
rlabel metal1 108560 43690 108560 43690 0 _047_
rlabel metal1 108691 38250 108691 38250 0 _048_
rlabel metal1 108790 50218 108790 50218 0 _049_
rlabel metal1 116334 30226 116334 30226 0 _050_
rlabel metal1 116840 30838 116840 30838 0 _051_
rlabel metal2 115598 28220 115598 28220 0 _052_
rlabel metal1 115598 35632 115598 35632 0 _053_
rlabel metal1 114632 29546 114632 29546 0 _054_
rlabel metal1 114310 35088 114310 35088 0 _055_
rlabel metal1 109802 27506 109802 27506 0 _056_
rlabel metal2 117162 31008 117162 31008 0 _057_
rlabel metal2 116518 30396 116518 30396 0 _058_
rlabel metal1 115414 30294 115414 30294 0 _059_
rlabel metal1 115736 30022 115736 30022 0 _060_
rlabel metal1 116028 30294 116028 30294 0 _061_
rlabel metal2 115874 29818 115874 29818 0 _062_
rlabel metal2 116610 29818 116610 29818 0 _063_
rlabel metal1 116058 29172 116058 29172 0 _064_
rlabel metal1 115552 29614 115552 29614 0 _065_
rlabel metal2 115966 29308 115966 29308 0 _066_
rlabel metal2 114770 29036 114770 29036 0 _067_
rlabel metal1 117990 30260 117990 30260 0 _068_
rlabel metal1 117576 28186 117576 28186 0 _069_
rlabel metal1 117668 29206 117668 29206 0 _070_
rlabel metal2 117438 29648 117438 29648 0 _071_
rlabel metal1 118036 27438 118036 27438 0 _072_
rlabel metal2 117622 27948 117622 27948 0 _073_
rlabel metal1 115874 29172 115874 29172 0 _074_
rlabel metal1 115322 29206 115322 29206 0 _075_
rlabel metal1 115414 28730 115414 28730 0 _076_
rlabel metal1 114172 29002 114172 29002 0 _077_
rlabel metal2 114954 27914 114954 27914 0 _078_
rlabel metal2 116702 28492 116702 28492 0 _079_
rlabel metal2 116886 28492 116886 28492 0 _080_
rlabel metal1 117530 27948 117530 27948 0 _081_
rlabel metal1 117484 27574 117484 27574 0 _082_
rlabel metal1 115046 27982 115046 27982 0 _083_
rlabel metal2 115046 27642 115046 27642 0 _084_
rlabel metal1 114172 27574 114172 27574 0 _085_
rlabel metal1 116380 27370 116380 27370 0 _086_
rlabel metal1 116426 27438 116426 27438 0 _087_
rlabel metal2 115414 27234 115414 27234 0 _088_
rlabel metal2 115322 27302 115322 27302 0 _089_
rlabel metal1 115598 26554 115598 26554 0 _090_
rlabel metal1 114678 28084 114678 28084 0 _091_
rlabel metal1 115000 26350 115000 26350 0 _092_
rlabel metal1 114172 26894 114172 26894 0 _093_
rlabel metal2 114494 27846 114494 27846 0 _094_
rlabel metal1 113574 34544 113574 34544 0 _095_
rlabel metal1 111274 38930 111274 38930 0 _096_
rlabel metal1 113988 27098 113988 27098 0 _097_
rlabel metal1 113436 28186 113436 28186 0 _098_
rlabel metal1 111550 26962 111550 26962 0 _099_
rlabel metal1 114954 25738 114954 25738 0 _100_
rlabel metal1 114402 26554 114402 26554 0 _101_
rlabel metal2 109894 28016 109894 28016 0 _102_
rlabel metal2 112194 27166 112194 27166 0 _103_
rlabel metal2 111274 27234 111274 27234 0 _104_
rlabel metal1 113988 28458 113988 28458 0 _105_
rlabel metal2 113574 28356 113574 28356 0 _106_
rlabel metal1 110262 29172 110262 29172 0 _107_
rlabel metal1 112194 28560 112194 28560 0 _108_
rlabel metal1 112608 28458 112608 28458 0 _109_
rlabel metal2 112010 28900 112010 28900 0 _110_
rlabel metal2 112286 27642 112286 27642 0 _111_
rlabel metal1 111182 27404 111182 27404 0 _112_
rlabel metal1 111044 27982 111044 27982 0 _113_
rlabel metal2 114218 29988 114218 29988 0 _114_
rlabel via1 111734 28067 111734 28067 0 _115_
rlabel metal1 111182 34680 111182 34680 0 _116_
rlabel metal1 110124 31790 110124 31790 0 _117_
rlabel metal1 111826 27506 111826 27506 0 _118_
rlabel metal2 111918 29121 111918 29121 0 _119_
rlabel metal1 110216 27438 110216 27438 0 _120_
rlabel metal2 109986 27846 109986 27846 0 _121_
rlabel metal2 111090 27812 111090 27812 0 _122_
rlabel metal1 110170 28730 110170 28730 0 _123_
rlabel metal1 110584 28526 110584 28526 0 _124_
rlabel metal2 111734 29172 111734 29172 0 _125_
rlabel metal2 110630 30022 110630 30022 0 _126_
rlabel metal1 111964 30566 111964 30566 0 _127_
rlabel metal1 110722 29274 110722 29274 0 _128_
rlabel metal1 110446 29002 110446 29002 0 _129_
rlabel metal1 109526 29648 109526 29648 0 _130_
rlabel metal1 109526 29818 109526 29818 0 _131_
rlabel metal1 110170 30906 110170 30906 0 _132_
rlabel metal1 110078 30158 110078 30158 0 _133_
rlabel metal1 110814 30158 110814 30158 0 _134_
rlabel metal2 109250 30532 109250 30532 0 _135_
rlabel metal1 111320 32402 111320 32402 0 _136_
rlabel metal1 113298 29750 113298 29750 0 _137_
rlabel metal1 111734 30192 111734 30192 0 _138_
rlabel metal1 112378 30702 112378 30702 0 _139_
rlabel via1 114311 32402 114311 32402 0 _140_
rlabel metal1 109572 30906 109572 30906 0 _141_
rlabel metal1 113344 30634 113344 30634 0 _142_
rlabel metal2 113850 31008 113850 31008 0 _143_
rlabel metal1 111504 32334 111504 32334 0 _144_
rlabel metal1 111090 31450 111090 31450 0 _145_
rlabel metal2 110906 32028 110906 32028 0 _146_
rlabel metal2 112746 33184 112746 33184 0 _147_
rlabel metal2 113298 32045 113298 32045 0 _148_
rlabel metal1 113298 32436 113298 32436 0 _149_
rlabel metal1 113068 31790 113068 31790 0 _150_
rlabel metal1 112976 31926 112976 31926 0 _151_
rlabel metal1 113620 30362 113620 30362 0 _152_
rlabel metal1 114264 30566 114264 30566 0 _153_
rlabel metal1 112378 29716 112378 29716 0 _154_
rlabel metal1 112194 29478 112194 29478 0 _155_
rlabel metal1 113160 30226 113160 30226 0 _156_
rlabel metal1 114126 31280 114126 31280 0 _157_
rlabel metal1 113850 33422 113850 33422 0 _158_
rlabel metal1 114632 30770 114632 30770 0 _159_
rlabel metal1 114494 30906 114494 30906 0 _160_
rlabel metal1 114319 30294 114319 30294 0 _161_
rlabel metal1 113620 30294 113620 30294 0 _162_
rlabel metal1 113850 30192 113850 30192 0 _163_
rlabel metal1 115230 32878 115230 32878 0 _164_
rlabel metal1 112378 33388 112378 33388 0 _165_
rlabel metal1 113436 33626 113436 33626 0 _166_
rlabel metal1 114218 33592 114218 33592 0 _167_
rlabel metal2 117806 32844 117806 32844 0 _168_
rlabel metal1 116242 32266 116242 32266 0 _169_
rlabel metal1 114402 32538 114402 32538 0 _170_
rlabel metal1 112930 32334 112930 32334 0 _171_
rlabel metal1 113758 32334 113758 32334 0 _172_
rlabel metal2 115966 32062 115966 32062 0 _173_
rlabel metal2 117530 32351 117530 32351 0 _174_
rlabel metal1 116518 31994 116518 31994 0 _175_
rlabel metal1 115782 32368 115782 32368 0 _176_
rlabel metal2 117714 32708 117714 32708 0 _177_
rlabel metal2 116242 32708 116242 32708 0 _178_
rlabel metal1 114632 33490 114632 33490 0 _179_
rlabel metal1 117254 31994 117254 31994 0 _180_
rlabel metal1 117714 33898 117714 33898 0 _181_
rlabel metal2 117346 35632 117346 35632 0 _182_
rlabel metal1 117944 34170 117944 34170 0 _183_
rlabel metal1 117668 34918 117668 34918 0 _184_
rlabel metal2 116058 33524 116058 33524 0 _185_
rlabel metal2 115414 32198 115414 32198 0 _186_
rlabel metal2 115690 33014 115690 33014 0 _187_
rlabel metal2 115598 34068 115598 34068 0 _188_
rlabel metal1 117852 34510 117852 34510 0 _189_
rlabel metal1 116472 34034 116472 34034 0 _190_
rlabel metal1 117806 34442 117806 34442 0 _191_
rlabel via1 118266 35462 118266 35462 0 _192_
rlabel metal2 118174 32742 118174 32742 0 _193_
rlabel metal2 117714 33252 117714 33252 0 _194_
rlabel metal1 117622 33626 117622 33626 0 _195_
rlabel metal2 117070 34238 117070 34238 0 _196_
rlabel metal1 116104 34714 116104 34714 0 _197_
rlabel metal1 116564 35258 116564 35258 0 _198_
rlabel metal2 116978 35972 116978 35972 0 _199_
rlabel metal1 116748 36754 116748 36754 0 _200_
rlabel metal1 115644 36006 115644 36006 0 _201_
rlabel metal1 115000 33626 115000 33626 0 _202_
rlabel metal1 115138 33898 115138 33898 0 _203_
rlabel metal1 115322 34170 115322 34170 0 _204_
rlabel metal1 114678 34476 114678 34476 0 _205_
rlabel metal1 114770 35088 114770 35088 0 _206_
rlabel metal1 114356 34918 114356 34918 0 _207_
rlabel viali 114218 34580 114218 34580 0 _208_
rlabel metal1 115552 36142 115552 36142 0 _209_
rlabel metal2 116978 36550 116978 36550 0 _210_
rlabel metal1 115782 36652 115782 36652 0 _211_
rlabel metal1 117714 35666 117714 35666 0 _212_
rlabel metal2 117438 36006 117438 36006 0 _213_
rlabel metal1 115690 36278 115690 36278 0 _214_
rlabel metal1 115874 36074 115874 36074 0 _215_
rlabel metal1 115966 36822 115966 36822 0 _216_
rlabel metal1 114816 35802 114816 35802 0 _217_
rlabel metal1 115092 37230 115092 37230 0 _218_
rlabel via2 114034 36771 114034 36771 0 _219_
rlabel metal2 115230 35258 115230 35258 0 _220_
rlabel metal1 113528 34170 113528 34170 0 _221_
rlabel metal1 113390 34952 113390 34952 0 _222_
rlabel metal1 113344 35734 113344 35734 0 _223_
rlabel metal1 113574 36108 113574 36108 0 _224_
rlabel metal2 114402 36992 114402 36992 0 _225_
rlabel metal2 116242 36992 116242 36992 0 _226_
rlabel metal1 114770 37128 114770 37128 0 _227_
rlabel metal1 114356 36822 114356 36822 0 _228_
rlabel metal1 114816 36890 114816 36890 0 _229_
rlabel metal2 113482 39168 113482 39168 0 _230_
rlabel metal1 113712 35802 113712 35802 0 _231_
rlabel metal1 112378 35190 112378 35190 0 _232_
rlabel metal2 114126 35734 114126 35734 0 _233_
rlabel metal1 112145 36142 112145 36142 0 _234_
rlabel metal2 111642 35428 111642 35428 0 _235_
rlabel metal2 111918 36278 111918 36278 0 _236_
rlabel metal1 112516 36550 112516 36550 0 _237_
rlabel metal2 112470 35700 112470 35700 0 _238_
rlabel metal2 112562 36720 112562 36720 0 _239_
rlabel metal1 113758 36788 113758 36788 0 _240_
rlabel metal2 114678 36822 114678 36822 0 _241_
rlabel metal2 113942 36652 113942 36652 0 _242_
rlabel metal2 112470 36992 112470 36992 0 _243_
rlabel metal2 110906 39304 110906 39304 0 _244_
rlabel metal1 111918 37162 111918 37162 0 _245_
rlabel metal1 110630 32946 110630 32946 0 _246_
rlabel metal1 109618 34544 109618 34544 0 _247_
rlabel metal1 110262 33626 110262 33626 0 _248_
rlabel metal1 109273 31994 109273 31994 0 _249_
rlabel metal2 110354 33218 110354 33218 0 _250_
rlabel metal1 110354 33490 110354 33490 0 _251_
rlabel metal1 110078 33082 110078 33082 0 _252_
rlabel metal1 109480 32334 109480 32334 0 _253_
rlabel metal1 110308 34374 110308 34374 0 _254_
rlabel metal2 109618 33762 109618 33762 0 _255_
rlabel metal1 110906 35598 110906 35598 0 _256_
rlabel metal2 110814 36516 110814 36516 0 _257_
rlabel metal1 111638 34714 111638 34714 0 _258_
rlabel metal1 110630 35190 110630 35190 0 _259_
rlabel metal2 111274 37502 111274 37502 0 _260_
rlabel metal1 110952 37434 110952 37434 0 _261_
rlabel metal1 110768 41514 110768 41514 0 _262_
rlabel metal1 110814 40086 110814 40086 0 _263_
rlabel metal1 110630 40052 110630 40052 0 _264_
rlabel metal1 111108 36686 111108 36686 0 _265_
rlabel metal1 111136 36822 111136 36822 0 _266_
rlabel metal2 110722 35598 110722 35598 0 _267_
rlabel metal1 111036 34646 111036 34646 0 _268_
rlabel metal1 110492 34034 110492 34034 0 _269_
rlabel metal1 109940 33966 109940 33966 0 _270_
rlabel via1 110547 34442 110547 34442 0 _271_
rlabel metal1 109756 43690 109756 43690 0 _272_
rlabel metal1 109250 45288 109250 45288 0 _273_
rlabel metal1 109434 45050 109434 45050 0 _274_
rlabel metal1 109940 43418 109940 43418 0 _275_
rlabel metal2 109894 43248 109894 43248 0 _276_
rlabel metal1 109802 38794 109802 38794 0 _277_
rlabel metal2 110354 39882 110354 39882 0 _278_
rlabel metal1 110078 40154 110078 40154 0 _279_
rlabel metal1 109342 37672 109342 37672 0 _280_
rlabel metal2 109342 36856 109342 36856 0 _281_
rlabel metal1 109526 34544 109526 34544 0 _282_
rlabel metal1 109158 35258 109158 35258 0 _283_
rlabel via1 109066 35717 109066 35717 0 _284_
rlabel metal2 108514 34272 108514 34272 0 _285_
rlabel metal2 109434 35530 109434 35530 0 _286_
rlabel metal2 109250 35360 109250 35360 0 _287_
rlabel metal1 109296 41650 109296 41650 0 _288_
rlabel metal2 108882 35632 108882 35632 0 _289_
rlabel metal1 109894 41786 109894 41786 0 _290_
rlabel metal2 25806 1520 25806 1520 0 addr00[0]
rlabel metal1 1380 35666 1380 35666 0 addr00[1]
rlabel metal1 1380 37842 1380 37842 0 addr00[2]
rlabel metal1 1334 38318 1334 38318 0 addr00[3]
rlabel metal1 1380 40494 1380 40494 0 addr00[4]
rlabel metal1 1380 41106 1380 41106 0 addr00[5]
rlabel metal1 1380 43282 1380 43282 0 addr00[6]
rlabel metal1 1380 44370 1380 44370 0 addr00[7]
rlabel metal2 107870 98311 107870 98311 0 clk
rlabel metal1 57132 97002 57132 97002 0 clknet_0_clk
rlabel metal4 15886 9968 15886 9968 0 clknet_3_0__leaf_clk
rlabel metal1 55660 94418 55660 94418 0 clknet_3_1__leaf_clk
rlabel metal2 56258 96798 56258 96798 0 clknet_3_2__leaf_clk
rlabel metal2 67482 95982 67482 95982 0 clknet_3_3__leaf_clk
rlabel metal1 109158 57902 109158 57902 0 clknet_3_4__leaf_clk
rlabel metal2 109618 51102 109618 51102 0 clknet_3_5__leaf_clk
rlabel metal2 70794 93500 70794 93500 0 clknet_3_6__leaf_clk
rlabel metal4 100070 89775 100070 89775 0 clknet_3_7__leaf_clk
rlabel metal1 1380 16082 1380 16082 0 csb00
rlabel metal2 118542 28815 118542 28815 0 denum[0]
rlabel metal2 118266 27999 118266 27999 0 denum[1]
rlabel metal1 118588 28526 118588 28526 0 denum[2]
rlabel metal2 118266 28917 118266 28917 0 denum[3]
rlabel metal2 31602 1520 31602 1520 0 din00[0]
rlabel metal2 43194 1520 43194 1520 0 din00[10]
rlabel metal2 44482 1520 44482 1520 0 din00[11]
rlabel metal2 45770 1520 45770 1520 0 din00[12]
rlabel metal2 46414 1520 46414 1520 0 din00[13]
rlabel metal2 47702 1520 47702 1520 0 din00[14]
rlabel metal2 48990 1520 48990 1520 0 din00[15]
rlabel metal2 32890 1520 32890 1520 0 din00[1]
rlabel metal2 33534 1520 33534 1520 0 din00[2]
rlabel metal2 34822 1520 34822 1520 0 din00[3]
rlabel metal2 36110 1520 36110 1520 0 din00[4]
rlabel metal2 37398 1520 37398 1520 0 din00[5]
rlabel metal2 38042 1520 38042 1520 0 din00[6]
rlabel metal2 39974 1520 39974 1520 0 din00[7]
rlabel metal2 40618 1520 40618 1520 0 din00[8]
rlabel metal2 41906 1520 41906 1520 0 din00[9]
rlabel metal2 50278 1520 50278 1520 0 din01[0]
rlabel metal2 61870 1520 61870 1520 0 din01[10]
rlabel metal2 63158 1520 63158 1520 0 din01[11]
rlabel metal2 63802 1520 63802 1520 0 din01[12]
rlabel metal2 65090 1520 65090 1520 0 din01[13]
rlabel metal1 66562 2278 66562 2278 0 din01[14]
rlabel metal2 67666 1520 67666 1520 0 din01[15]
rlabel metal2 51566 1520 51566 1520 0 din01[1]
rlabel metal2 52210 1520 52210 1520 0 din01[2]
rlabel metal2 53498 1520 53498 1520 0 din01[3]
rlabel metal2 54786 1520 54786 1520 0 din01[4]
rlabel metal2 56074 1520 56074 1520 0 din01[5]
rlabel metal2 57362 1520 57362 1520 0 din01[6]
rlabel metal2 58006 1520 58006 1520 0 din01[7]
rlabel metal2 59294 1520 59294 1520 0 din01[8]
rlabel metal2 60582 1520 60582 1520 0 din01[9]
rlabel metal4 25542 9968 25542 9968 0 net1
rlabel metal1 117760 28050 117760 28050 0 net10
rlabel metal1 109342 43350 109342 43350 0 net100
rlabel metal4 89462 89571 89462 89571 0 net101
rlabel metal1 68770 93840 68770 93840 0 net102
rlabel metal1 72312 93398 72312 93398 0 net103
rlabel metal1 108468 44370 108468 44370 0 net104
rlabel metal1 117484 31382 117484 31382 0 net105
rlabel metal1 113482 36754 113482 36754 0 net106
rlabel metal1 116472 32878 116472 32878 0 net107
rlabel metal1 114908 31790 114908 31790 0 net108
rlabel metal1 116564 33966 116564 33966 0 net109
rlabel metal1 117300 28526 117300 28526 0 net11
rlabel metal1 116334 31926 116334 31926 0 net110
rlabel metal1 113252 28458 113252 28458 0 net111
rlabel metal1 114310 33830 114310 33830 0 net112
rlabel metal3 106068 86470 106068 86470 0 net113
rlabel metal3 9852 17246 9852 17246 0 net114
rlabel metal2 27002 8619 27002 8619 0 net115
rlabel metal1 27876 7514 27876 7514 0 net116
rlabel metal2 29578 8619 29578 8619 0 net117
rlabel metal2 30222 8619 30222 8619 0 net118
rlabel metal1 109848 43826 109848 43826 0 net119
rlabel metal1 117898 28492 117898 28492 0 net12
rlabel metal1 110032 45458 110032 45458 0 net120
rlabel metal2 109618 45050 109618 45050 0 net121
rlabel metal1 118082 29648 118082 29648 0 net13
rlabel metal4 31390 9968 31390 9968 0 net14
rlabel metal4 43086 9968 43086 9968 0 net15
rlabel metal4 44174 9968 44174 9968 0 net16
rlabel metal4 45534 9968 45534 9968 0 net17
rlabel metal4 46622 9968 46622 9968 0 net18
rlabel metal4 47710 9968 47710 9968 0 net19
rlabel metal1 4255 35802 4255 35802 0 net2
rlabel metal4 48934 9968 48934 9968 0 net20
rlabel metal4 32614 9968 32614 9968 0 net21
rlabel metal4 33702 9968 33702 9968 0 net22
rlabel metal1 34960 2618 34960 2618 0 net23
rlabel metal4 36150 9968 36150 9968 0 net24
rlabel metal4 37238 9968 37238 9968 0 net25
rlabel metal4 38326 9968 38326 9968 0 net26
rlabel via2 40066 2635 40066 2635 0 net27
rlabel metal4 40774 9968 40774 9968 0 net28
rlabel metal4 41862 9968 41862 9968 0 net29
rlabel metal2 9522 37608 9522 37608 0 net3
rlabel metal4 50294 9968 50294 9968 0 net30
rlabel metal4 61854 9868 61854 9868 0 net31
rlabel metal4 62942 9868 62942 9868 0 net32
rlabel metal4 64030 9868 64030 9868 0 net33
rlabel metal4 65254 9968 65254 9968 0 net34
rlabel metal1 66700 2618 66700 2618 0 net35
rlabel metal4 67702 9900 67702 9900 0 net36
rlabel metal4 51382 9900 51382 9900 0 net37
rlabel metal4 52470 9900 52470 9900 0 net38
rlabel metal4 53558 9900 53558 9900 0 net39
rlabel metal1 1610 38216 1610 38216 0 net4
rlabel metal4 54918 9900 54918 9900 0 net40
rlabel metal4 56006 9900 56006 9900 0 net41
rlabel metal4 57094 9900 57094 9900 0 net42
rlabel metal4 58318 9900 58318 9900 0 net43
rlabel metal4 59406 9900 59406 9900 0 net44
rlabel metal4 60766 9968 60766 9968 0 net45
rlabel metal2 117990 30940 117990 30940 0 net46
rlabel metal2 118358 31178 118358 31178 0 net47
rlabel metal1 116978 32266 116978 32266 0 net48
rlabel metal1 117162 31790 117162 31790 0 net49
rlabel metal1 1610 40392 1610 40392 0 net5
rlabel metal1 107962 96934 107962 96934 0 net50
rlabel metal2 57454 96356 57454 96356 0 net51
rlabel metal1 67942 96186 67942 96186 0 net52
rlabel metal1 69276 95098 69276 95098 0 net53
rlabel metal1 70012 95370 70012 95370 0 net54
rlabel metal1 71852 95642 71852 95642 0 net55
rlabel metal2 72542 96084 72542 96084 0 net56
rlabel metal1 73830 96186 73830 96186 0 net57
rlabel metal1 58374 96186 58374 96186 0 net58
rlabel metal1 59478 95098 59478 95098 0 net59
rlabel metal2 9706 41076 9706 41076 0 net6
rlabel metal1 60996 95642 60996 95642 0 net60
rlabel metal2 60582 95812 60582 95812 0 net61
rlabel metal2 62882 96356 62882 96356 0 net62
rlabel metal1 63664 95098 63664 95098 0 net63
rlabel metal2 64998 96356 64998 96356 0 net64
rlabel metal1 66792 95642 66792 95642 0 net65
rlabel metal2 67390 96084 67390 96084 0 net66
rlabel metal2 112838 37604 112838 37604 0 net67
rlabel metal2 114494 35326 114494 35326 0 net68
rlabel metal1 116426 35666 116426 35666 0 net69
rlabel metal2 9706 43048 9706 43048 0 net7
rlabel metal2 117622 32164 117622 32164 0 net70
rlabel metal1 116794 32436 116794 32436 0 net71
rlabel metal1 112194 32198 112194 32198 0 net72
rlabel metal1 111918 32198 111918 32198 0 net73
rlabel metal1 110814 31926 110814 31926 0 net74
rlabel metal2 115690 27132 115690 27132 0 net75
rlabel metal1 56488 94894 56488 94894 0 net76
rlabel metal1 65136 93874 65136 93874 0 net77
rlabel metal4 93380 9112 93380 9112 0 net78
rlabel metal1 109342 33864 109342 33864 0 net79
rlabel metal1 4255 44234 4255 44234 0 net8
rlabel metal2 93058 8704 93058 8704 0 net80
rlabel metal2 109158 33286 109158 33286 0 net81
rlabel metal1 109434 33558 109434 33558 0 net82
rlabel metal2 92874 8738 92874 8738 0 net83
rlabel metal1 108514 32232 108514 32232 0 net84
rlabel metal1 109986 32436 109986 32436 0 net85
rlabel metal2 93426 8772 93426 8772 0 net86
rlabel metal1 109572 32402 109572 32402 0 net87
rlabel metal1 109986 35598 109986 35598 0 net88
rlabel metal3 106789 23596 106789 23596 0 net89
rlabel metal2 9706 15780 9706 15780 0 net9
rlabel metal1 110308 36142 110308 36142 0 net90
rlabel metal3 106743 24956 106743 24956 0 net91
rlabel metal1 110722 37876 110722 37876 0 net92
rlabel metal1 110124 43146 110124 43146 0 net93
rlabel metal2 110170 42874 110170 42874 0 net94
rlabel metal3 106697 26588 106697 26588 0 net95
rlabel metal1 110538 39372 110538 39372 0 net96
rlabel metal1 109434 42636 109434 42636 0 net99
rlabel metal2 118542 30481 118542 30481 0 num[0]
rlabel metal2 118542 31909 118542 31909 0 num[1]
rlabel metal2 118542 27353 118542 27353 0 num[2]
rlabel via2 118542 31331 118542 31331 0 num[3]
rlabel metal2 107502 98277 107502 98277 0 rst
rlabel metal1 55706 97274 55706 97274 0 sine_out[0]
rlabel metal2 67850 98277 67850 98277 0 sine_out[10]
rlabel metal1 69000 96458 69000 96458 0 sine_out[11]
rlabel metal2 70334 98277 70334 98277 0 sine_out[12]
rlabel metal2 71714 98277 71714 98277 0 sine_out[13]
rlabel metal2 72358 98277 72358 98277 0 sine_out[14]
rlabel metal2 74382 98277 74382 98277 0 sine_out[15]
rlabel metal1 57868 97274 57868 97274 0 sine_out[1]
rlabel metal2 58834 98311 58834 98311 0 sine_out[2]
rlabel metal2 60674 98311 60674 98311 0 sine_out[3]
rlabel metal2 60122 98311 60122 98311 0 sine_out[4]
rlabel metal2 62698 98311 62698 98311 0 sine_out[5]
rlabel metal2 63342 98311 63342 98311 0 sine_out[6]
rlabel metal2 64630 98311 64630 98311 0 sine_out[7]
rlabel metal2 65274 98311 65274 98311 0 sine_out[8]
rlabel metal2 67206 98277 67206 98277 0 sine_out[9]
rlabel metal2 46966 93024 46966 93024 0 sine_out_reg0\[0\]
rlabel metal2 64722 92497 64722 92497 0 sine_out_reg0\[10\]
rlabel metal2 61318 92752 61318 92752 0 sine_out_reg0\[11\]
rlabel metal1 60306 92344 60306 92344 0 sine_out_reg0\[12\]
rlabel metal1 64998 92106 64998 92106 0 sine_out_reg0\[13\]
rlabel metal1 64124 92582 64124 92582 0 sine_out_reg0\[14\]
rlabel metal1 65826 92582 65826 92582 0 sine_out_reg0\[15\]
rlabel metal1 53728 94418 53728 94418 0 sine_out_reg0\[1\]
rlabel metal1 55798 94758 55798 94758 0 sine_out_reg0\[2\]
rlabel metal1 56718 93262 56718 93262 0 sine_out_reg0\[3\]
rlabel metal2 58466 94129 58466 94129 0 sine_out_reg0\[4\]
rlabel metal2 56258 93262 56258 93262 0 sine_out_reg0\[5\]
rlabel metal2 56350 93194 56350 93194 0 sine_out_reg0\[6\]
rlabel metal2 56074 92072 56074 92072 0 sine_out_reg0\[7\]
rlabel metal1 55338 92888 55338 92888 0 sine_out_reg0\[8\]
rlabel metal2 63802 94044 63802 94044 0 sine_out_reg0\[9\]
rlabel metal2 55798 93534 55798 93534 0 sine_out_reg1\[0\]
rlabel metal2 68586 92990 68586 92990 0 sine_out_reg1\[10\]
rlabel metal2 68310 92922 68310 92922 0 sine_out_reg1\[11\]
rlabel metal1 70702 92922 70702 92922 0 sine_out_reg1\[12\]
rlabel metal1 68770 93262 68770 93262 0 sine_out_reg1\[13\]
rlabel metal1 71760 92922 71760 92922 0 sine_out_reg1\[14\]
rlabel metal1 72726 92106 72726 92106 0 sine_out_reg1\[15\]
rlabel metal1 55982 92922 55982 92922 0 sine_out_reg1\[1\]
rlabel metal2 57822 94418 57822 94418 0 sine_out_reg1\[2\]
rlabel metal1 57270 93228 57270 93228 0 sine_out_reg1\[3\]
rlabel metal1 59202 94554 59202 94554 0 sine_out_reg1\[4\]
rlabel metal2 60674 93568 60674 93568 0 sine_out_reg1\[5\]
rlabel metal1 62514 93466 62514 93466 0 sine_out_reg1\[6\]
rlabel metal1 64170 93126 64170 93126 0 sine_out_reg1\[7\]
rlabel metal1 64630 92922 64630 92922 0 sine_out_reg1\[8\]
rlabel metal1 66424 92922 66424 92922 0 sine_out_reg1\[9\]
rlabel metal2 44206 92599 44206 92599 0 sine_out_temp0\[0\]
rlabel metal1 56380 92310 56380 92310 0 sine_out_temp0\[10\]
rlabel via2 58006 92803 58006 92803 0 sine_out_temp0\[11\]
rlabel via2 58742 92123 58742 92123 0 sine_out_temp0\[12\]
rlabel metal2 60582 90831 60582 90831 0 sine_out_temp0\[13\]
rlabel metal2 59294 91239 59294 91239 0 sine_out_temp0\[14\]
rlabel metal4 56948 91528 56948 91528 0 sine_out_temp0\[15\]
rlabel metal4 39652 91392 39652 91392 0 sine_out_temp0\[1\]
rlabel metal4 40638 89571 40638 89571 0 sine_out_temp0\[2\]
rlabel metal4 42044 91664 42044 91664 0 sine_out_temp0\[3\]
rlabel metal4 43332 91120 43332 91120 0 sine_out_temp0\[4\]
rlabel metal4 44620 91460 44620 91460 0 sine_out_temp0\[5\]
rlabel via1 52573 92650 52573 92650 0 sine_out_temp0\[6\]
rlabel via2 53222 92021 53222 92021 0 sine_out_temp0\[7\]
rlabel metal1 55361 92718 55361 92718 0 sine_out_temp0\[8\]
rlabel via2 55614 93925 55614 93925 0 sine_out_temp0\[9\]
rlabel metal4 58182 89707 58182 89707 0 sine_out_temp1\[0\]
rlabel metal4 70694 89575 70694 89575 0 sine_out_temp1\[10\]
rlabel metal4 71918 89571 71918 89571 0 sine_out_temp1\[11\]
rlabel metal4 73278 89575 73278 89575 0 sine_out_temp1\[12\]
rlabel metal4 74366 89575 74366 89575 0 sine_out_temp1\[13\]
rlabel metal4 75590 89571 75590 89571 0 sine_out_temp1\[14\]
rlabel metal3 76448 89692 76448 89692 0 sine_out_temp1\[15\]
rlabel metal4 59542 89707 59542 89707 0 sine_out_temp1\[1\]
rlabel metal4 60630 89571 60630 89571 0 sine_out_temp1\[2\]
rlabel metal2 59846 93007 59846 93007 0 sine_out_temp1\[3\]
rlabel metal4 63078 89575 63078 89575 0 sine_out_temp1\[4\]
rlabel metal4 64302 89575 64302 89575 0 sine_out_temp1\[5\]
rlabel metal3 65468 89692 65468 89692 0 sine_out_temp1\[6\]
rlabel metal4 66886 89571 66886 89571 0 sine_out_temp1\[7\]
rlabel metal4 68246 89571 68246 89571 0 sine_out_temp1\[8\]
rlabel metal4 69334 89575 69334 89575 0 sine_out_temp1\[9\]
rlabel metal1 109480 44846 109480 44846 0 tcout\[0\]
rlabel metal1 108698 45458 108698 45458 0 tcout\[1\]
rlabel metal1 109296 43282 109296 43282 0 tcout\[2\]
rlabel metal1 109066 41990 109066 41990 0 tcout\[3\]
rlabel metal1 110308 35054 110308 35054 0 tcout\[4\]
rlabel metal2 108330 35020 108330 35020 0 tcout\[5\]
rlabel metal2 109066 34272 109066 34272 0 tcout\[6\]
rlabel metal1 109526 34000 109526 34000 0 tcout\[7\]
rlabel metal1 109710 41616 109710 41616 0 tcout\[8\]
rlabel metal1 109158 67354 109158 67354 0 tcout_delay\[0\]
rlabel metal1 109628 67218 109628 67218 0 tcout_delay\[1\]
<< properties >>
string FIXED_BBOX 0 0 120000 100000
<< end >>
