magic
tech sky130A
magscale 1 2
timestamp 1741277098
<< viali >>
rect 85497 136969 85531 137003
rect 85046 136833 85080 136867
rect 85313 136833 85347 136867
rect 83657 136629 83691 136663
rect 83933 136629 83967 136663
rect 85681 136629 85715 136663
rect 34345 136221 34379 136255
rect 34161 136153 34195 136187
rect 34713 136153 34747 136187
rect 34989 136153 35023 136187
rect 35173 136153 35207 136187
rect 36185 136153 36219 136187
rect 43177 136153 43211 136187
rect 47777 136153 47811 136187
rect 50353 136153 50387 136187
rect 55413 136153 55447 136187
rect 57989 136153 58023 136187
rect 60565 136153 60599 136187
rect 60749 136153 60783 136187
rect 63141 136153 63175 136187
rect 72525 136153 72559 136187
rect 73445 136153 73479 136187
rect 77401 136153 77435 136187
rect 35357 136085 35391 136119
rect 36093 136085 36127 136119
rect 36369 136085 36403 136119
rect 43085 136085 43119 136119
rect 43361 136085 43395 136119
rect 46121 136085 46155 136119
rect 47685 136085 47719 136119
rect 47961 136085 47995 136119
rect 50261 136085 50295 136119
rect 50537 136085 50571 136119
rect 55505 136085 55539 136119
rect 55781 136085 55815 136119
rect 58081 136085 58115 136119
rect 58357 136085 58391 136119
rect 60933 136085 60967 136119
rect 63233 136085 63267 136119
rect 63509 136085 63543 136119
rect 63601 136085 63635 136119
rect 68569 136085 68603 136119
rect 72617 136085 72651 136119
rect 72893 136085 72927 136119
rect 73537 136085 73571 136119
rect 73813 136085 73847 136119
rect 77493 136085 77527 136119
rect 77769 136085 77803 136119
rect 86325 136085 86359 136119
rect 87337 136085 87371 136119
rect 95985 136085 96019 136119
rect 104357 129761 104391 129795
rect 7481 118473 7515 118507
rect 6193 117725 6227 117759
rect 6460 117657 6494 117691
rect 7573 117589 7607 117623
rect 7297 117045 7331 117079
rect 7481 117045 7515 117079
rect 106013 113577 106047 113611
rect 104357 113441 104391 113475
rect 104624 113373 104658 113407
rect 105737 113237 105771 113271
rect 105829 113237 105863 113271
rect 104449 113033 104483 113067
rect 1593 111333 1627 111367
rect 1409 111197 1443 111231
rect 1685 111197 1719 111231
rect 1409 109633 1443 109667
rect 1685 109633 1719 109667
rect 1593 109497 1627 109531
rect 1409 108545 1443 108579
rect 1685 108545 1719 108579
rect 1593 108409 1627 108443
rect 105645 107049 105679 107083
rect 106381 107049 106415 107083
rect 1593 106981 1627 107015
rect 1409 106845 1443 106879
rect 1685 106845 1719 106879
rect 104357 106777 104391 106811
rect 106289 106777 106323 106811
rect 1593 105893 1627 105927
rect 1409 105757 1443 105791
rect 1685 105757 1719 105791
rect 1409 104193 1443 104227
rect 1685 104193 1719 104227
rect 1593 104057 1627 104091
rect 7573 101065 7607 101099
rect 104624 100997 104658 101031
rect 104357 100861 104391 100895
rect 106013 100793 106047 100827
rect 105737 100725 105771 100759
rect 105829 100725 105863 100759
rect 104449 100521 104483 100555
rect 6193 100317 6227 100351
rect 6460 100249 6494 100283
rect 7573 100181 7607 100215
rect 7481 99977 7515 100011
rect 7297 99637 7331 99671
rect 104613 96577 104647 96611
rect 104357 96509 104391 96543
rect 106013 96441 106047 96475
rect 105737 96373 105771 96407
rect 105829 96373 105863 96407
rect 104357 96169 104391 96203
rect 7481 95625 7515 95659
rect 104357 95285 104391 95319
rect 7481 94945 7515 94979
rect 5733 94809 5767 94843
rect 5825 94809 5859 94843
rect 6561 94401 6595 94435
rect 6653 94401 6687 94435
rect 6193 93789 6227 93823
rect 6460 93721 6494 93755
rect 7573 93653 7607 93687
rect 104357 93653 104391 93687
rect 7389 93449 7423 93483
rect 7113 93109 7147 93143
rect 7481 93109 7515 93143
rect 104357 92565 104391 92599
rect 104357 91545 104391 91579
rect 105093 91545 105127 91579
rect 105369 91545 105403 91579
rect 104357 91069 104391 91103
rect 1501 88961 1535 88995
rect 1961 88961 1995 88995
rect 1685 88825 1719 88859
rect 1869 88825 1903 88859
rect 1501 87873 1535 87907
rect 1961 87873 1995 87907
rect 1685 87737 1719 87771
rect 1869 87737 1903 87771
rect 1501 87193 1535 87227
rect 1961 87193 1995 87227
rect 1593 87125 1627 87159
rect 1869 87125 1903 87159
rect 1501 86785 1535 86819
rect 1961 86785 1995 86819
rect 1685 86649 1719 86683
rect 1869 86649 1903 86683
rect 1409 86173 1443 86207
rect 1685 86173 1719 86207
rect 1593 86037 1627 86071
rect 1501 85017 1535 85051
rect 1961 85017 1995 85051
rect 1593 84949 1627 84983
rect 1869 84949 1903 84983
rect 1501 84609 1535 84643
rect 1961 84609 1995 84643
rect 1685 84473 1719 84507
rect 1777 84473 1811 84507
rect 1409 83997 1443 84031
rect 1961 83997 1995 84031
rect 1593 83861 1627 83895
rect 1869 83861 1903 83895
rect 1501 83521 1535 83555
rect 1961 83521 1995 83555
rect 1593 83317 1627 83351
rect 1869 83317 1903 83351
rect 1501 82433 1535 82467
rect 1961 82433 1995 82467
rect 4997 82433 5031 82467
rect 4261 82365 4295 82399
rect 5181 82365 5215 82399
rect 1593 82229 1627 82263
rect 1869 82229 1903 82263
rect 5365 82229 5399 82263
rect 1501 81753 1535 81787
rect 1961 81753 1995 81787
rect 1593 81685 1627 81719
rect 1869 81685 1903 81719
rect 1501 81345 1535 81379
rect 1961 81345 1995 81379
rect 1685 81209 1719 81243
rect 1869 81209 1903 81243
rect 1409 80733 1443 80767
rect 1685 80733 1719 80767
rect 108221 80733 108255 80767
rect 108497 80733 108531 80767
rect 2421 80597 2455 80631
rect 1409 80325 1443 80359
rect 108497 80325 108531 80359
rect 108221 79645 108255 79679
rect 1501 79577 1535 79611
rect 1685 79577 1719 79611
rect 1869 79577 1903 79611
rect 1961 79509 1995 79543
rect 108405 79509 108439 79543
rect 1501 79169 1535 79203
rect 1961 79169 1995 79203
rect 108221 79169 108255 79203
rect 1685 79033 1719 79067
rect 1869 79033 1903 79067
rect 108405 78965 108439 78999
rect 108221 78557 108255 78591
rect 1501 78489 1535 78523
rect 1685 78489 1719 78523
rect 1869 78489 1903 78523
rect 1961 78421 1995 78455
rect 108405 78421 108439 78455
rect 1501 78081 1535 78115
rect 1961 78081 1995 78115
rect 108221 78081 108255 78115
rect 1685 77945 1719 77979
rect 1869 77945 1903 77979
rect 108405 77877 108439 77911
rect 16681 77673 16715 77707
rect 26065 77673 26099 77707
rect 26985 77673 27019 77707
rect 28181 77673 28215 77707
rect 29561 77673 29595 77707
rect 30481 77673 30515 77707
rect 31769 77673 31803 77707
rect 32873 77673 32907 77707
rect 33977 77673 34011 77707
rect 35265 77673 35299 77707
rect 36369 77673 36403 77707
rect 37473 77673 37507 77707
rect 38669 77673 38703 77707
rect 39865 77673 39899 77707
rect 41061 77673 41095 77707
rect 42165 77673 42199 77707
rect 43361 77673 43395 77707
rect 94973 77673 95007 77707
rect 14749 77605 14783 77639
rect 25789 77605 25823 77639
rect 87245 77605 87279 77639
rect 89453 77605 89487 77639
rect 90465 77605 90499 77639
rect 91109 77605 91143 77639
rect 94145 77605 94179 77639
rect 98929 77605 98963 77639
rect 83749 77537 83783 77571
rect 85957 77537 85991 77571
rect 86417 77537 86451 77571
rect 86601 77537 86635 77571
rect 90649 77537 90683 77571
rect 94605 77537 94639 77571
rect 16497 77469 16531 77503
rect 24133 77469 24167 77503
rect 24409 77469 24443 77503
rect 24665 77469 24699 77503
rect 25881 77469 25915 77503
rect 54493 77469 54527 77503
rect 83933 77469 83967 77503
rect 84577 77469 84611 77503
rect 90005 77469 90039 77503
rect 93777 77469 93811 77503
rect 94053 77469 94087 77503
rect 94881 77469 94915 77503
rect 95157 77469 95191 77503
rect 97181 77469 97215 77503
rect 16221 77401 16255 77435
rect 55137 77401 55171 77435
rect 55321 77401 55355 77435
rect 89545 77401 89579 77435
rect 89729 77401 89763 77435
rect 91477 77401 91511 77435
rect 94697 77401 94731 77435
rect 97457 77401 97491 77435
rect 14657 77333 14691 77367
rect 23489 77333 23523 77367
rect 56609 77333 56643 77367
rect 57161 77333 57195 77367
rect 83381 77333 83415 77367
rect 84025 77333 84059 77367
rect 84393 77333 84427 77367
rect 86693 77333 86727 77367
rect 87061 77333 87095 77367
rect 89913 77333 89947 77367
rect 91569 77333 91603 77367
rect 91845 77333 91879 77367
rect 92489 77333 92523 77367
rect 94329 77333 94363 77367
rect 99113 77333 99147 77367
rect 1593 77129 1627 77163
rect 1869 77129 1903 77163
rect 88533 77129 88567 77163
rect 89545 77129 89579 77163
rect 90189 77129 90223 77163
rect 91753 77129 91787 77163
rect 97641 77129 97675 77163
rect 22385 77061 22419 77095
rect 24685 77061 24719 77095
rect 25881 77061 25915 77095
rect 89085 77061 89119 77095
rect 99481 77061 99515 77095
rect 1501 76993 1535 77027
rect 1961 76993 1995 77027
rect 22477 76993 22511 77027
rect 25789 76993 25823 77027
rect 89177 76993 89211 77027
rect 89729 76993 89763 77027
rect 90373 76993 90407 77027
rect 90557 76993 90591 77027
rect 91385 76993 91419 77027
rect 91937 76993 91971 77027
rect 92121 76993 92155 77027
rect 92673 76993 92707 77027
rect 93961 76993 93995 77027
rect 94237 76993 94271 77027
rect 95801 76993 95835 77027
rect 99113 76993 99147 77027
rect 99297 76993 99331 77027
rect 99573 76993 99607 77027
rect 100493 76993 100527 77027
rect 100677 76993 100711 77027
rect 108221 76993 108255 77027
rect 26065 76925 26099 76959
rect 88901 76925 88935 76959
rect 91109 76925 91143 76959
rect 91293 76925 91327 76959
rect 96077 76925 96111 76959
rect 25237 76857 25271 76891
rect 90833 76857 90867 76891
rect 97549 76857 97583 76891
rect 108405 76857 108439 76891
rect 22569 76789 22603 76823
rect 25421 76789 25455 76823
rect 26341 76789 26375 76823
rect 55045 76789 55079 76823
rect 90465 76789 90499 76823
rect 93133 76789 93167 76823
rect 94053 76789 94087 76823
rect 99205 76789 99239 76823
rect 100493 76789 100527 76823
rect 41337 76585 41371 76619
rect 46949 76585 46983 76619
rect 60473 76585 60507 76619
rect 67005 76585 67039 76619
rect 94513 76585 94547 76619
rect 23213 76517 23247 76551
rect 23029 76449 23063 76483
rect 23673 76449 23707 76483
rect 23857 76449 23891 76483
rect 24133 76449 24167 76483
rect 27353 76449 27387 76483
rect 29009 76449 29043 76483
rect 29101 76449 29135 76483
rect 60749 76449 60783 76483
rect 82829 76449 82863 76483
rect 93041 76449 93075 76483
rect 98101 76449 98135 76483
rect 100585 76449 100619 76483
rect 101045 76449 101079 76483
rect 1685 76381 1719 76415
rect 26525 76381 26559 76415
rect 27169 76381 27203 76415
rect 27629 76381 27663 76415
rect 41245 76381 41279 76415
rect 41613 76381 41647 76415
rect 44281 76381 44315 76415
rect 44649 76381 44683 76415
rect 46857 76381 46891 76415
rect 47133 76381 47167 76415
rect 62865 76381 62899 76415
rect 64337 76381 64371 76415
rect 65625 76381 65659 76415
rect 67189 76381 67223 76415
rect 67649 76381 67683 76415
rect 85129 76381 85163 76415
rect 85221 76381 85255 76415
rect 92765 76381 92799 76415
rect 98469 76381 98503 76415
rect 98653 76381 98687 76415
rect 99021 76381 99055 76415
rect 99665 76381 99699 76415
rect 99849 76381 99883 76415
rect 101137 76381 101171 76415
rect 108221 76381 108255 76415
rect 28917 76313 28951 76347
rect 40978 76313 41012 76347
rect 44014 76313 44048 76347
rect 44373 76313 44407 76347
rect 46612 76313 46646 76347
rect 60289 76313 60323 76347
rect 61016 76313 61050 76347
rect 62773 76313 62807 76347
rect 63132 76313 63166 76347
rect 65441 76313 65475 76347
rect 65892 76313 65926 76347
rect 67557 76313 67591 76347
rect 67916 76313 67950 76347
rect 69121 76313 69155 76347
rect 83013 76313 83047 76347
rect 84862 76313 84896 76347
rect 97825 76313 97859 76347
rect 99297 76313 99331 76347
rect 99389 76313 99423 76347
rect 100309 76313 100343 76347
rect 1501 76245 1535 76279
rect 23581 76245 23615 76279
rect 26709 76245 26743 76279
rect 27077 76245 27111 76279
rect 28549 76245 28583 76279
rect 29653 76245 29687 76279
rect 39865 76245 39899 76279
rect 42901 76245 42935 76279
rect 45477 76245 45511 76279
rect 62129 76245 62163 76279
rect 64245 76245 64279 76279
rect 69029 76245 69063 76279
rect 82553 76245 82587 76279
rect 83105 76245 83139 76279
rect 83473 76245 83507 76279
rect 83657 76245 83691 76279
rect 83749 76245 83783 76279
rect 92581 76245 92615 76279
rect 99941 76245 99975 76279
rect 100401 76245 100435 76279
rect 100769 76245 100803 76279
rect 108037 76245 108071 76279
rect 108405 76245 108439 76279
rect 14657 76041 14691 76075
rect 83749 76041 83783 76075
rect 90081 76041 90115 76075
rect 90833 76041 90867 76075
rect 96905 76041 96939 76075
rect 100769 76041 100803 76075
rect 108405 76041 108439 76075
rect 90281 75973 90315 76007
rect 99481 75973 99515 76007
rect 1685 75905 1719 75939
rect 16497 75905 16531 75939
rect 90741 75905 90775 75939
rect 91109 75905 91143 75939
rect 98285 75905 98319 75939
rect 98561 75905 98595 75939
rect 98653 75905 98687 75939
rect 98745 75905 98779 75939
rect 98929 75905 98963 75939
rect 99265 75905 99299 75939
rect 99389 75905 99423 75939
rect 99665 75905 99699 75939
rect 99757 75905 99791 75939
rect 100585 75905 100619 75939
rect 108221 75905 108255 75939
rect 14749 75837 14783 75871
rect 16221 75837 16255 75871
rect 95157 75837 95191 75871
rect 95433 75837 95467 75871
rect 97825 75837 97859 75871
rect 97917 75837 97951 75871
rect 100401 75837 100435 75871
rect 88165 75769 88199 75803
rect 88901 75769 88935 75803
rect 108037 75769 108071 75803
rect 1501 75701 1535 75735
rect 87981 75701 88015 75735
rect 89913 75701 89947 75735
rect 90097 75701 90131 75735
rect 94973 75701 95007 75735
rect 97641 75701 97675 75735
rect 98377 75701 98411 75735
rect 99113 75701 99147 75735
rect 22293 75497 22327 75531
rect 94881 75497 94915 75531
rect 99021 75497 99055 75531
rect 102885 75497 102919 75531
rect 103253 75497 103287 75531
rect 104633 75497 104667 75531
rect 108037 75497 108071 75531
rect 87705 75429 87739 75463
rect 88349 75429 88383 75463
rect 98101 75429 98135 75463
rect 100769 75429 100803 75463
rect 103529 75429 103563 75463
rect 105001 75429 105035 75463
rect 87981 75361 88015 75395
rect 93409 75361 93443 75395
rect 97181 75361 97215 75395
rect 101321 75361 101355 75395
rect 101965 75361 101999 75395
rect 1685 75293 1719 75327
rect 22385 75293 22419 75327
rect 25605 75293 25639 75327
rect 88717 75293 88751 75327
rect 93133 75293 93167 75327
rect 98285 75293 98319 75327
rect 98377 75293 98411 75327
rect 98929 75293 98963 75327
rect 99113 75293 99147 75327
rect 100309 75293 100343 75327
rect 100493 75293 100527 75327
rect 102057 75293 102091 75327
rect 102793 75293 102827 75327
rect 102977 75293 103011 75327
rect 103805 75293 103839 75327
rect 103897 75293 103931 75327
rect 103989 75293 104023 75327
rect 104173 75293 104207 75327
rect 105093 75293 105127 75327
rect 105185 75293 105219 75327
rect 105369 75293 105403 75327
rect 108221 75293 108255 75327
rect 25513 75225 25547 75259
rect 88165 75225 88199 75259
rect 88993 75225 89027 75259
rect 90741 75225 90775 75259
rect 98101 75225 98135 75259
rect 101137 75225 101171 75259
rect 103221 75225 103255 75259
rect 103437 75225 103471 75259
rect 103529 75225 103563 75259
rect 103713 75225 103747 75259
rect 104817 75225 104851 75259
rect 1501 75157 1535 75191
rect 22569 75157 22603 75191
rect 25697 75157 25731 75191
rect 87521 75157 87555 75191
rect 90925 75157 90959 75191
rect 92949 75157 92983 75191
rect 97365 75157 97399 75191
rect 97457 75157 97491 75191
rect 97825 75157 97859 75191
rect 100493 75157 100527 75191
rect 101229 75157 101263 75191
rect 101689 75157 101723 75191
rect 103069 75157 103103 75191
rect 104357 75157 104391 75191
rect 104449 75157 104483 75191
rect 104617 75157 104651 75191
rect 105277 75157 105311 75191
rect 108405 75157 108439 75191
rect 18061 74953 18095 74987
rect 88257 74953 88291 74987
rect 89637 74953 89671 74987
rect 90925 74953 90959 74987
rect 91661 74953 91695 74987
rect 92213 74953 92247 74987
rect 96997 74953 97031 74987
rect 100033 74953 100067 74987
rect 100959 74953 100993 74987
rect 104081 74953 104115 74987
rect 87797 74885 87831 74919
rect 88349 74885 88383 74919
rect 98285 74885 98319 74919
rect 101045 74885 101079 74919
rect 101597 74885 101631 74919
rect 104449 74885 104483 74919
rect 19901 74817 19935 74851
rect 88073 74817 88107 74851
rect 89545 74817 89579 74851
rect 89821 74817 89855 74851
rect 91201 74817 91235 74851
rect 91477 74817 91511 74851
rect 91753 74817 91787 74851
rect 91845 74817 91879 74851
rect 91937 74817 91971 74851
rect 92121 74817 92155 74851
rect 92397 74817 92431 74851
rect 94421 74817 94455 74851
rect 96629 74817 96663 74851
rect 97365 74817 97399 74851
rect 97457 74817 97491 74851
rect 97549 74817 97583 74851
rect 97733 74817 97767 74851
rect 98009 74817 98043 74851
rect 98469 74817 98503 74851
rect 98745 74817 98779 74851
rect 99297 74817 99331 74851
rect 99757 74817 99791 74851
rect 99941 74817 99975 74851
rect 100125 74817 100159 74851
rect 100217 74817 100251 74851
rect 100309 74817 100343 74851
rect 100493 74817 100527 74851
rect 100585 74817 100619 74851
rect 100861 74817 100895 74851
rect 101137 74817 101171 74851
rect 101413 74817 101447 74851
rect 101781 74817 101815 74851
rect 101965 74817 101999 74851
rect 102057 74817 102091 74851
rect 102149 74817 102183 74851
rect 102333 74817 102367 74851
rect 103069 74817 103103 74851
rect 103253 74817 103287 74851
rect 103345 74817 103379 74851
rect 103529 74817 103563 74851
rect 103713 74817 103747 74851
rect 105185 74817 105219 74851
rect 18153 74749 18187 74783
rect 19625 74749 19659 74783
rect 86049 74749 86083 74783
rect 89453 74749 89487 74783
rect 94513 74749 94547 74783
rect 96721 74749 96755 74783
rect 99481 74749 99515 74783
rect 99573 74749 99607 74783
rect 102241 74749 102275 74783
rect 103161 74749 103195 74783
rect 104909 74749 104943 74783
rect 105093 74749 105127 74783
rect 99389 74681 99423 74715
rect 101229 74681 101263 74715
rect 104725 74681 104759 74715
rect 88993 74613 89027 74647
rect 91293 74613 91327 74647
rect 91845 74613 91879 74647
rect 94145 74613 94179 74647
rect 97089 74613 97123 74647
rect 99113 74613 99147 74647
rect 100769 74613 100803 74647
rect 103621 74613 103655 74647
rect 103805 74613 103839 74647
rect 105461 74613 105495 74647
rect 21741 74409 21775 74443
rect 23323 74409 23357 74443
rect 74733 74409 74767 74443
rect 75101 74409 75135 74443
rect 85681 74409 85715 74443
rect 85957 74409 85991 74443
rect 87521 74409 87555 74443
rect 91569 74409 91603 74443
rect 96721 74409 96755 74443
rect 99941 74409 99975 74443
rect 101781 74409 101815 74443
rect 102885 74409 102919 74443
rect 1501 74341 1535 74375
rect 90097 74341 90131 74375
rect 90281 74341 90315 74375
rect 100401 74341 100435 74375
rect 101505 74341 101539 74375
rect 104449 74341 104483 74375
rect 21833 74273 21867 74307
rect 28181 74273 28215 74307
rect 88349 74273 88383 74307
rect 88625 74273 88659 74307
rect 96905 74273 96939 74307
rect 101965 74273 101999 74307
rect 102793 74273 102827 74307
rect 105369 74273 105403 74307
rect 105461 74273 105495 74307
rect 1685 74205 1719 74239
rect 1869 74205 1903 74239
rect 23581 74205 23615 74239
rect 24593 74205 24627 74239
rect 24777 74205 24811 74239
rect 28273 74205 28307 74239
rect 28457 74205 28491 74239
rect 29745 74205 29779 74239
rect 74917 74205 74951 74239
rect 85589 74205 85623 74239
rect 87153 74205 87187 74239
rect 91477 74205 91511 74239
rect 91753 74205 91787 74239
rect 96997 74205 97031 74239
rect 97912 74205 97946 74239
rect 98101 74205 98135 74239
rect 98284 74205 98318 74239
rect 98377 74205 98411 74239
rect 100125 74205 100159 74239
rect 100217 74205 100251 74239
rect 100389 74205 100423 74239
rect 100585 74205 100619 74239
rect 101321 74205 101355 74239
rect 102057 74205 102091 74239
rect 102885 74205 102919 74239
rect 103253 74205 103287 74239
rect 104449 74205 104483 74239
rect 104725 74205 104759 74239
rect 105277 74205 105311 74239
rect 108221 74205 108255 74239
rect 23949 74137 23983 74171
rect 87245 74137 87279 74171
rect 98009 74137 98043 74171
rect 104633 74137 104667 74171
rect 108037 74137 108071 74171
rect 23673 74069 23707 74103
rect 24501 74069 24535 74103
rect 29653 74069 29687 74103
rect 29929 74069 29963 74103
rect 90465 74069 90499 74103
rect 97733 74069 97767 74103
rect 102517 74069 102551 74103
rect 103069 74069 103103 74103
rect 104909 74069 104943 74103
rect 108405 74069 108439 74103
rect 35541 73865 35575 73899
rect 68477 73865 68511 73899
rect 68937 73865 68971 73899
rect 70133 73865 70167 73899
rect 74457 73865 74491 73899
rect 75101 73865 75135 73899
rect 84853 73865 84887 73899
rect 87429 73865 87463 73899
rect 87613 73865 87647 73899
rect 93317 73865 93351 73899
rect 98837 73865 98871 73899
rect 101965 73865 101999 73899
rect 104909 73865 104943 73899
rect 105277 73865 105311 73899
rect 108313 73865 108347 73899
rect 85957 73797 85991 73831
rect 90817 73797 90851 73831
rect 91017 73797 91051 73831
rect 91201 73797 91235 73831
rect 102517 73797 102551 73831
rect 104633 73797 104667 73831
rect 105645 73797 105679 73831
rect 1685 73729 1719 73763
rect 11621 73729 11655 73763
rect 18981 73729 19015 73763
rect 27997 73729 28031 73763
rect 28181 73729 28215 73763
rect 35449 73729 35483 73763
rect 55229 73729 55263 73763
rect 55321 73729 55355 73763
rect 68569 73729 68603 73763
rect 70225 73729 70259 73763
rect 73813 73729 73847 73763
rect 74549 73729 74583 73763
rect 84945 73729 84979 73763
rect 85129 73729 85163 73763
rect 88809 73729 88843 73763
rect 93501 73729 93535 73763
rect 93685 73729 93719 73763
rect 94145 73729 94179 73763
rect 94421 73729 94455 73763
rect 94605 73729 94639 73763
rect 98653 73729 98687 73763
rect 98929 73729 98963 73763
rect 99113 73729 99147 73763
rect 99297 73729 99331 73763
rect 100033 73729 100067 73763
rect 100493 73729 100527 73763
rect 100677 73729 100711 73763
rect 101873 73729 101907 73763
rect 102333 73729 102367 73763
rect 102977 73729 103011 73763
rect 103161 73729 103195 73763
rect 103437 73729 103471 73763
rect 104265 73729 104299 73763
rect 104358 73729 104392 73763
rect 104541 73729 104575 73763
rect 104730 73729 104764 73763
rect 105185 73729 105219 73763
rect 105369 73729 105403 73763
rect 105829 73729 105863 73763
rect 108221 73729 108255 73763
rect 108497 73729 108531 73763
rect 13369 73661 13403 73695
rect 18705 73661 18739 73695
rect 24777 73661 24811 73695
rect 25053 73661 25087 73695
rect 25421 73661 25455 73695
rect 35633 73661 35667 73695
rect 35909 73661 35943 73695
rect 68293 73661 68327 73695
rect 69121 73661 69155 73695
rect 69949 73661 69983 73695
rect 70685 73661 70719 73695
rect 73537 73661 73571 73695
rect 73905 73661 73939 73695
rect 74365 73661 74399 73695
rect 85681 73661 85715 73695
rect 89085 73661 89119 73695
rect 90557 73661 90591 73695
rect 99573 73661 99607 73695
rect 99849 73661 99883 73695
rect 100217 73661 100251 73695
rect 100309 73661 100343 73695
rect 100401 73661 100435 73695
rect 102701 73661 102735 73695
rect 105461 73661 105495 73695
rect 1501 73593 1535 73627
rect 13553 73593 13587 73627
rect 17141 73593 17175 73627
rect 74917 73593 74951 73627
rect 90649 73593 90683 73627
rect 98653 73593 98687 73627
rect 99481 73593 99515 73627
rect 1869 73525 1903 73559
rect 11253 73525 11287 73559
rect 17233 73525 17267 73559
rect 23305 73525 23339 73559
rect 25145 73525 25179 73559
rect 27905 73525 27939 73559
rect 35081 73525 35115 73559
rect 56793 73525 56827 73559
rect 57253 73525 57287 73559
rect 70593 73525 70627 73559
rect 85589 73525 85623 73559
rect 90833 73525 90867 73559
rect 91385 73525 91419 73559
rect 93593 73525 93627 73559
rect 93961 73525 93995 73559
rect 99389 73525 99423 73559
rect 103621 73525 103655 73559
rect 21465 73321 21499 73355
rect 23305 73321 23339 73355
rect 23581 73321 23615 73355
rect 88165 73321 88199 73355
rect 93777 73321 93811 73355
rect 98561 73321 98595 73355
rect 98745 73321 98779 73355
rect 99573 73321 99607 73355
rect 100585 73321 100619 73355
rect 100769 73321 100803 73355
rect 101689 73321 101723 73355
rect 102977 73321 103011 73355
rect 103345 73321 103379 73355
rect 103805 73321 103839 73355
rect 70501 73253 70535 73287
rect 78781 73253 78815 73287
rect 106197 73253 106231 73287
rect 1869 73185 1903 73219
rect 23213 73185 23247 73219
rect 37933 73185 37967 73219
rect 38209 73185 38243 73219
rect 40417 73185 40451 73219
rect 40693 73185 40727 73219
rect 72433 73185 72467 73219
rect 78689 73185 78723 73219
rect 80161 73185 80195 73219
rect 95525 73185 95559 73219
rect 95893 73185 95927 73219
rect 97365 73185 97399 73219
rect 97917 73185 97951 73219
rect 100401 73185 100435 73219
rect 102241 73185 102275 73219
rect 102793 73185 102827 73219
rect 103621 73185 103655 73219
rect 104541 73185 104575 73219
rect 1685 73117 1719 73151
rect 40325 73117 40359 73151
rect 72617 73117 72651 73151
rect 73169 73117 73203 73151
rect 87797 73117 87831 73151
rect 87889 73117 87923 73151
rect 95709 73117 95743 73151
rect 96997 73117 97031 73151
rect 97089 73117 97123 73151
rect 97181 73117 97215 73151
rect 97641 73117 97675 73151
rect 97733 73117 97767 73151
rect 97825 73117 97859 73151
rect 98101 73117 98135 73151
rect 98193 73117 98227 73151
rect 98377 73117 98411 73151
rect 98653 73117 98687 73151
rect 99481 73117 99515 73151
rect 99757 73117 99791 73151
rect 100309 73117 100343 73151
rect 100493 73117 100527 73151
rect 101045 73117 101079 73151
rect 102977 73117 103011 73151
rect 103897 73117 103931 73151
rect 104081 73117 104115 73151
rect 105645 73117 105679 73151
rect 106013 73117 106047 73151
rect 106289 73117 106323 73151
rect 108221 73117 108255 73151
rect 108497 73117 108531 73151
rect 22937 73049 22971 73083
rect 40233 73049 40267 73083
rect 70133 73049 70167 73083
rect 70225 73049 70259 73083
rect 72709 73049 72743 73083
rect 79916 73049 79950 73083
rect 100953 73049 100987 73083
rect 101229 73049 101263 73083
rect 101413 73049 101447 73083
rect 102057 73049 102091 73083
rect 102517 73049 102551 73083
rect 104173 73049 104207 73083
rect 1501 72981 1535 73015
rect 37381 72981 37415 73015
rect 37749 72981 37783 73015
rect 37841 72981 37875 73015
rect 39865 72981 39899 73015
rect 68845 72981 68879 73015
rect 73077 72981 73111 73015
rect 96813 72981 96847 73015
rect 97457 72981 97491 73015
rect 99205 72981 99239 73015
rect 100743 72981 100777 73015
rect 102149 72981 102183 73015
rect 103161 72981 103195 73015
rect 104265 72981 104299 73015
rect 105461 72981 105495 73015
rect 105829 72981 105863 73015
rect 108313 72981 108347 73015
rect 69121 72777 69155 72811
rect 86233 72777 86267 72811
rect 88165 72777 88199 72811
rect 97739 72777 97773 72811
rect 98377 72777 98411 72811
rect 100033 72777 100067 72811
rect 100861 72777 100895 72811
rect 104817 72777 104851 72811
rect 105369 72777 105403 72811
rect 88349 72709 88383 72743
rect 97641 72709 97675 72743
rect 98561 72709 98595 72743
rect 99113 72709 99147 72743
rect 102793 72709 102827 72743
rect 102977 72709 103011 72743
rect 105001 72709 105035 72743
rect 1685 72641 1719 72675
rect 1869 72641 1903 72675
rect 68845 72641 68879 72675
rect 96445 72641 96479 72675
rect 97825 72641 97859 72675
rect 97917 72641 97951 72675
rect 98285 72641 98319 72675
rect 98745 72641 98779 72675
rect 99297 72641 99331 72675
rect 100401 72641 100435 72675
rect 101045 72641 101079 72675
rect 101137 72641 101171 72675
rect 101597 72641 101631 72675
rect 101781 72641 101815 72675
rect 101873 72641 101907 72675
rect 103529 72641 103563 72675
rect 103713 72641 103747 72675
rect 103805 72641 103839 72675
rect 104357 72641 104391 72675
rect 104633 72641 104667 72675
rect 104909 72641 104943 72675
rect 105185 72641 105219 72675
rect 105461 72641 105495 72675
rect 105737 72641 105771 72675
rect 105921 72641 105955 72675
rect 106013 72641 106047 72675
rect 106289 72641 106323 72675
rect 108221 72641 108255 72675
rect 108497 72641 108531 72675
rect 86417 72573 86451 72607
rect 86693 72573 86727 72607
rect 96537 72573 96571 72607
rect 99481 72573 99515 72607
rect 100493 72573 100527 72607
rect 100585 72573 100619 72607
rect 104541 72573 104575 72607
rect 106105 72573 106139 72607
rect 96813 72505 96847 72539
rect 101597 72505 101631 72539
rect 104449 72505 104483 72539
rect 105599 72505 105633 72539
rect 1501 72437 1535 72471
rect 86049 72437 86083 72471
rect 98101 72437 98135 72471
rect 102609 72437 102643 72471
rect 103621 72437 103655 72471
rect 103989 72437 104023 72471
rect 105829 72437 105863 72471
rect 106013 72437 106047 72471
rect 106473 72437 106507 72471
rect 108313 72437 108347 72471
rect 82001 72233 82035 72267
rect 85497 72233 85531 72267
rect 88717 72233 88751 72267
rect 99021 72233 99055 72267
rect 101229 72233 101263 72267
rect 104357 72233 104391 72267
rect 85681 72165 85715 72199
rect 98469 72165 98503 72199
rect 96813 72097 96847 72131
rect 97089 72097 97123 72131
rect 97457 72097 97491 72131
rect 98377 72097 98411 72131
rect 99573 72097 99607 72131
rect 83125 72029 83159 72063
rect 83381 72029 83415 72063
rect 85405 72029 85439 72063
rect 88441 72029 88475 72063
rect 93409 72029 93443 72063
rect 93557 72029 93591 72063
rect 93915 72029 93949 72063
rect 96721 72029 96755 72063
rect 97549 72029 97583 72063
rect 97641 72029 97675 72063
rect 98101 72029 98135 72063
rect 98285 72029 98319 72063
rect 98561 72029 98595 72063
rect 99757 72029 99791 72063
rect 100033 72029 100067 72063
rect 100217 72029 100251 72063
rect 101137 72029 101171 72063
rect 101321 72029 101355 72063
rect 102241 72029 102275 72063
rect 103069 72029 103103 72063
rect 103161 72029 103195 72063
rect 103437 72029 103471 72063
rect 103529 72029 103563 72063
rect 104173 72029 104207 72063
rect 104541 72029 104575 72063
rect 104817 72029 104851 72063
rect 105277 72029 105311 72063
rect 105553 72029 105587 72063
rect 105645 72029 105679 72063
rect 105737 72029 105771 72063
rect 106197 72029 106231 72063
rect 88533 71961 88567 71995
rect 93685 71961 93719 71995
rect 93777 71961 93811 71995
rect 98745 71961 98779 71995
rect 99205 71961 99239 71995
rect 103253 71961 103287 71995
rect 105461 71961 105495 71995
rect 105921 71961 105955 71995
rect 83473 71893 83507 71927
rect 94053 71893 94087 71927
rect 98009 71893 98043 71927
rect 98837 71893 98871 71927
rect 99005 71893 99039 71927
rect 102333 71893 102367 71927
rect 102885 71893 102919 71927
rect 103897 71893 103931 71927
rect 105001 71893 105035 71927
rect 105093 71893 105127 71927
rect 105829 71893 105863 71927
rect 106013 71893 106047 71927
rect 91569 71689 91603 71723
rect 96905 71689 96939 71723
rect 98193 71689 98227 71723
rect 100493 71689 100527 71723
rect 101413 71689 101447 71723
rect 108313 71689 108347 71723
rect 89637 71621 89671 71655
rect 91385 71621 91419 71655
rect 96169 71621 96203 71655
rect 98561 71621 98595 71655
rect 102609 71621 102643 71655
rect 104357 71621 104391 71655
rect 1501 71553 1535 71587
rect 1961 71553 1995 71587
rect 97180 71553 97214 71587
rect 97273 71553 97307 71587
rect 97825 71553 97859 71587
rect 98009 71553 98043 71587
rect 98469 71553 98503 71587
rect 98745 71553 98779 71587
rect 99481 71553 99515 71587
rect 99573 71553 99607 71587
rect 99757 71553 99791 71587
rect 99849 71553 99883 71587
rect 100861 71553 100895 71587
rect 101321 71553 101355 71587
rect 101781 71553 101815 71587
rect 102241 71553 102275 71587
rect 102793 71553 102827 71587
rect 102977 71553 103011 71587
rect 103437 71553 103471 71587
rect 103529 71553 103563 71587
rect 103713 71553 103747 71587
rect 103805 71553 103839 71587
rect 104265 71553 104299 71587
rect 104449 71553 104483 71587
rect 104541 71553 104575 71587
rect 104725 71553 104759 71587
rect 105369 71553 105403 71587
rect 105645 71553 105679 71587
rect 107761 71553 107795 71587
rect 108497 71553 108531 71587
rect 89361 71485 89395 71519
rect 100769 71485 100803 71519
rect 101873 71485 101907 71519
rect 102885 71485 102919 71519
rect 105553 71485 105587 71519
rect 108221 71485 108255 71519
rect 1685 71417 1719 71451
rect 1869 71417 1903 71451
rect 95893 71417 95927 71451
rect 102149 71417 102183 71451
rect 104633 71417 104667 71451
rect 89177 71349 89211 71383
rect 95709 71349 95743 71383
rect 98929 71349 98963 71383
rect 99297 71349 99331 71383
rect 103989 71349 104023 71383
rect 105185 71349 105219 71383
rect 105829 71349 105863 71383
rect 107669 71349 107703 71383
rect 31585 71145 31619 71179
rect 33149 71145 33183 71179
rect 48605 71145 48639 71179
rect 74273 71145 74307 71179
rect 86325 71145 86359 71179
rect 92673 71145 92707 71179
rect 96537 71145 96571 71179
rect 99021 71145 99055 71179
rect 99573 71145 99607 71179
rect 100309 71145 100343 71179
rect 105829 71145 105863 71179
rect 108313 71145 108347 71179
rect 85681 71077 85715 71111
rect 92765 71077 92799 71111
rect 94145 71077 94179 71111
rect 97641 71077 97675 71111
rect 98561 71077 98595 71111
rect 106381 71077 106415 71111
rect 33057 71009 33091 71043
rect 48145 71009 48179 71043
rect 72617 71009 72651 71043
rect 72893 71009 72927 71043
rect 85957 71009 85991 71043
rect 88073 71009 88107 71043
rect 93133 71009 93167 71043
rect 94237 71009 94271 71043
rect 99941 71009 99975 71043
rect 103713 71009 103747 71043
rect 104265 71009 104299 71043
rect 104909 71009 104943 71043
rect 105093 71009 105127 71043
rect 105553 71009 105587 71043
rect 32873 70941 32907 70975
rect 47317 70941 47351 70975
rect 79241 70941 79275 70975
rect 79425 70941 79459 70975
rect 81081 70941 81115 70975
rect 85405 70941 85439 70975
rect 93225 70941 93259 70975
rect 93317 70941 93351 70975
rect 93409 70941 93443 70975
rect 93777 70941 93811 70975
rect 94421 70941 94455 70975
rect 96721 70941 96755 70975
rect 96997 70941 97031 70975
rect 97641 70941 97675 70975
rect 97825 70941 97859 70975
rect 98101 70941 98135 70975
rect 98469 70941 98503 70975
rect 98653 70941 98687 70975
rect 98929 70941 98963 70975
rect 99448 70941 99482 70975
rect 100033 70941 100067 70975
rect 101045 70941 101079 70975
rect 101873 70941 101907 70975
rect 102056 70941 102090 70975
rect 102149 70941 102183 70975
rect 102241 70941 102275 70975
rect 102425 70941 102459 70975
rect 104357 70941 104391 70975
rect 105185 70941 105219 70975
rect 106105 70941 106139 70975
rect 106381 70941 106415 70975
rect 108221 70941 108255 70975
rect 108497 70941 108531 70975
rect 48421 70873 48455 70907
rect 73138 70873 73172 70907
rect 79670 70873 79704 70907
rect 85497 70873 85531 70907
rect 87797 70873 87831 70907
rect 93961 70873 93995 70907
rect 102609 70873 102643 70907
rect 103529 70873 103563 70907
rect 106013 70873 106047 70907
rect 106197 70873 106231 70907
rect 72709 70805 72743 70839
rect 80805 70805 80839 70839
rect 92949 70805 92983 70839
rect 93593 70805 93627 70839
rect 93869 70805 93903 70839
rect 96905 70805 96939 70839
rect 98009 70805 98043 70839
rect 99389 70805 99423 70839
rect 101137 70805 101171 70839
rect 103161 70805 103195 70839
rect 103621 70805 103655 70839
rect 103989 70805 104023 70839
rect 105645 70805 105679 70839
rect 105813 70805 105847 70839
rect 30573 70601 30607 70635
rect 32137 70601 32171 70635
rect 34529 70601 34563 70635
rect 87981 70601 88015 70635
rect 93041 70601 93075 70635
rect 97089 70601 97123 70635
rect 99481 70601 99515 70635
rect 103621 70601 103655 70635
rect 106197 70601 106231 70635
rect 108313 70601 108347 70635
rect 34345 70533 34379 70567
rect 90189 70533 90223 70567
rect 91201 70533 91235 70567
rect 97641 70533 97675 70567
rect 98745 70533 98779 70567
rect 105829 70533 105863 70567
rect 106013 70533 106047 70567
rect 31686 70465 31720 70499
rect 31953 70465 31987 70499
rect 33261 70465 33295 70499
rect 33517 70465 33551 70499
rect 35653 70465 35687 70499
rect 35909 70465 35943 70499
rect 88165 70465 88199 70499
rect 90925 70465 90959 70499
rect 91109 70465 91143 70499
rect 96077 70465 96111 70499
rect 97273 70465 97307 70499
rect 97733 70465 97767 70499
rect 98193 70465 98227 70499
rect 98285 70465 98319 70499
rect 98469 70465 98503 70499
rect 98561 70465 98595 70499
rect 99297 70465 99331 70499
rect 99389 70465 99423 70499
rect 99573 70465 99607 70499
rect 100217 70465 100251 70499
rect 101965 70465 101999 70499
rect 103805 70465 103839 70499
rect 105185 70465 105219 70499
rect 106105 70465 106139 70499
rect 106289 70465 106323 70499
rect 108221 70465 108255 70499
rect 108497 70465 108531 70499
rect 88349 70397 88383 70431
rect 96169 70397 96203 70431
rect 97549 70397 97583 70431
rect 102057 70397 102091 70431
rect 103989 70397 104023 70431
rect 105277 70397 105311 70431
rect 105369 70397 105403 70431
rect 105461 70397 105495 70431
rect 96445 70329 96479 70363
rect 98101 70329 98135 70363
rect 99113 70329 99147 70363
rect 102333 70329 102367 70363
rect 93317 70261 93351 70295
rect 100033 70261 100067 70295
rect 105001 70261 105035 70295
rect 105645 70261 105679 70295
rect 32045 70057 32079 70091
rect 32229 70057 32263 70091
rect 35541 70057 35575 70091
rect 73353 70057 73387 70091
rect 75101 70057 75135 70091
rect 81173 70057 81207 70091
rect 89729 70057 89763 70091
rect 91569 70057 91603 70091
rect 97733 70057 97767 70091
rect 98469 70057 98503 70091
rect 99297 70057 99331 70091
rect 99941 70057 99975 70091
rect 100309 70057 100343 70091
rect 108313 70057 108347 70091
rect 35725 69989 35759 70023
rect 80897 69989 80931 70023
rect 91385 69989 91419 70023
rect 96353 69989 96387 70023
rect 97089 69989 97123 70023
rect 100861 69989 100895 70023
rect 37105 69921 37139 69955
rect 73721 69921 73755 69955
rect 79149 69921 79183 69955
rect 79517 69921 79551 69955
rect 89545 69921 89579 69955
rect 90097 69921 90131 69955
rect 90649 69921 90683 69955
rect 95065 69921 95099 69955
rect 96813 69921 96847 69955
rect 99849 69921 99883 69955
rect 101965 69921 101999 69955
rect 104633 69921 104667 69955
rect 77585 69853 77619 69887
rect 79333 69853 79367 69887
rect 90373 69853 90407 69887
rect 90465 69853 90499 69887
rect 91017 69853 91051 69887
rect 94053 69853 94087 69887
rect 94697 69853 94731 69887
rect 95157 69853 95191 69887
rect 96077 69853 96111 69887
rect 96721 69853 96755 69887
rect 97733 69853 97767 69887
rect 97917 69853 97951 69887
rect 98469 69853 98503 69887
rect 98653 69853 98687 69887
rect 99021 69853 99055 69887
rect 99113 69853 99147 69887
rect 99757 69853 99791 69887
rect 100217 69853 100251 69887
rect 100401 69853 100435 69887
rect 100493 69853 100527 69887
rect 100861 69853 100895 69887
rect 100953 69853 100987 69887
rect 101321 69853 101355 69887
rect 101505 69853 101539 69887
rect 101873 69853 101907 69887
rect 104449 69853 104483 69887
rect 105093 69853 105127 69887
rect 105185 69853 105219 69887
rect 105277 69853 105311 69887
rect 108221 69853 108255 69887
rect 108497 69853 108531 69887
rect 36860 69785 36894 69819
rect 73966 69785 74000 69819
rect 77493 69785 77527 69819
rect 77852 69785 77886 69819
rect 79784 69785 79818 69819
rect 94237 69785 94271 69819
rect 94421 69785 94455 69819
rect 96353 69785 96387 69819
rect 100769 69785 100803 69819
rect 101137 69785 101171 69819
rect 104541 69785 104575 69819
rect 30665 69717 30699 69751
rect 66729 69717 66763 69751
rect 73537 69717 73571 69751
rect 78965 69717 78999 69751
rect 94789 69717 94823 69751
rect 96169 69717 96203 69751
rect 99573 69717 99607 69751
rect 100033 69717 100067 69751
rect 100125 69717 100159 69751
rect 100677 69717 100711 69751
rect 101321 69717 101355 69751
rect 102241 69717 102275 69751
rect 104081 69717 104115 69751
rect 104909 69717 104943 69751
rect 42441 69513 42475 69547
rect 62865 69513 62899 69547
rect 68293 69513 68327 69547
rect 79517 69513 79551 69547
rect 88809 69513 88843 69547
rect 92105 69513 92139 69547
rect 97825 69513 97859 69547
rect 98009 69513 98043 69547
rect 100309 69513 100343 69547
rect 102609 69513 102643 69547
rect 63141 69445 63175 69479
rect 89545 69445 89579 69479
rect 91569 69445 91603 69479
rect 92305 69445 92339 69479
rect 100493 69445 100527 69479
rect 43565 69377 43599 69411
rect 61485 69377 61519 69411
rect 61741 69377 61775 69411
rect 66637 69377 66671 69411
rect 66893 69377 66927 69411
rect 89177 69377 89211 69411
rect 89453 69377 89487 69411
rect 91845 69377 91879 69411
rect 92581 69377 92615 69411
rect 98006 69377 98040 69411
rect 98377 69377 98411 69411
rect 98836 69377 98870 69411
rect 98929 69377 98963 69411
rect 99113 69377 99147 69411
rect 99297 69377 99331 69411
rect 99481 69377 99515 69411
rect 99665 69377 99699 69411
rect 99941 69377 99975 69411
rect 100217 69377 100251 69411
rect 101689 69377 101723 69411
rect 101873 69377 101907 69411
rect 102609 69377 102643 69411
rect 103345 69377 103379 69411
rect 103529 69377 103563 69411
rect 103805 69377 103839 69411
rect 103989 69377 104023 69411
rect 104817 69377 104851 69411
rect 105001 69377 105035 69411
rect 43821 69309 43855 69343
rect 66453 69309 66487 69343
rect 89085 69309 89119 69343
rect 89821 69309 89855 69343
rect 92857 69309 92891 69343
rect 98469 69309 98503 69343
rect 98561 69309 98595 69343
rect 102425 69309 102459 69343
rect 102977 69309 103011 69343
rect 99573 69241 99607 69275
rect 42165 69173 42199 69207
rect 61393 69173 61427 69207
rect 68017 69173 68051 69207
rect 91937 69173 91971 69207
rect 92121 69173 92155 69207
rect 92489 69173 92523 69207
rect 92765 69173 92799 69207
rect 99297 69173 99331 69207
rect 99757 69173 99791 69207
rect 100493 69173 100527 69207
rect 101781 69173 101815 69207
rect 103161 69173 103195 69207
rect 103621 69173 103655 69207
rect 104633 69173 104667 69207
rect 44741 68969 44775 69003
rect 58633 68969 58667 69003
rect 60289 68969 60323 69003
rect 67373 68969 67407 69003
rect 87061 68969 87095 69003
rect 90097 68969 90131 69003
rect 93593 68969 93627 69003
rect 98285 68969 98319 69003
rect 100585 68969 100619 69003
rect 103253 68969 103287 69003
rect 105093 68969 105127 69003
rect 105277 68969 105311 69003
rect 45017 68901 45051 68935
rect 67005 68901 67039 68935
rect 100769 68901 100803 68935
rect 46397 68833 46431 68867
rect 58909 68833 58943 68867
rect 65625 68833 65659 68867
rect 91661 68833 91695 68867
rect 94881 68833 94915 68867
rect 95525 68833 95559 68867
rect 95985 68833 96019 68867
rect 99941 68833 99975 68867
rect 102149 68833 102183 68867
rect 102241 68833 102275 68867
rect 102977 68833 103011 68867
rect 86693 68765 86727 68799
rect 89821 68765 89855 68799
rect 91385 68765 91419 68799
rect 93409 68765 93443 68799
rect 94789 68765 94823 68799
rect 95893 68765 95927 68799
rect 97089 68765 97123 68799
rect 97457 68765 97491 68799
rect 98377 68765 98411 68799
rect 99570 68765 99604 68799
rect 100033 68765 100067 68799
rect 100861 68765 100895 68799
rect 101045 68765 101079 68799
rect 103069 68765 103103 68799
rect 103345 68765 103379 68799
rect 103437 68765 103471 68799
rect 103621 68765 103655 68799
rect 103713 68765 103747 68799
rect 104541 68765 104575 68799
rect 104817 68765 104851 68799
rect 105001 68765 105035 68799
rect 42533 68697 42567 68731
rect 46152 68697 46186 68731
rect 58725 68697 58759 68731
rect 59154 68697 59188 68731
rect 65892 68697 65926 68731
rect 67097 68697 67131 68731
rect 91109 68697 91143 68731
rect 97181 68697 97215 68731
rect 97273 68697 97307 68731
rect 100401 68697 100435 68731
rect 100617 68697 100651 68731
rect 105245 68697 105279 68731
rect 105461 68697 105495 68731
rect 46489 68629 46523 68663
rect 61485 68629 61519 68663
rect 86785 68629 86819 68663
rect 89913 68629 89947 68663
rect 94513 68629 94547 68663
rect 95157 68629 95191 68663
rect 96905 68629 96939 68663
rect 99389 68629 99423 68663
rect 99573 68629 99607 68663
rect 101689 68629 101723 68663
rect 102057 68629 102091 68663
rect 102609 68629 102643 68663
rect 103897 68629 103931 68663
rect 104357 68629 104391 68663
rect 38669 68425 38703 68459
rect 38853 68425 38887 68459
rect 91569 68425 91603 68459
rect 91737 68425 91771 68459
rect 96261 68425 96295 68459
rect 96353 68425 96387 68459
rect 98193 68425 98227 68459
rect 100217 68425 100251 68459
rect 101781 68425 101815 68459
rect 101965 68425 101999 68459
rect 102977 68425 103011 68459
rect 103345 68425 103379 68459
rect 105093 68425 105127 68459
rect 91937 68357 91971 68391
rect 94973 68357 95007 68391
rect 100585 68357 100619 68391
rect 101413 68357 101447 68391
rect 39966 68289 40000 68323
rect 40233 68289 40267 68323
rect 95249 68289 95283 68323
rect 95801 68289 95835 68323
rect 95985 68289 96019 68323
rect 96169 68289 96203 68323
rect 96537 68289 96571 68323
rect 97089 68289 97123 68323
rect 97825 68289 97859 68323
rect 99113 68289 99147 68323
rect 99297 68289 99331 68323
rect 99573 68289 99607 68323
rect 99849 68289 99883 68323
rect 100401 68289 100435 68323
rect 100677 68289 100711 68323
rect 100769 68289 100803 68323
rect 101137 68289 101171 68323
rect 101597 68289 101631 68323
rect 101873 68289 101907 68323
rect 102149 68289 102183 68323
rect 103161 68289 103195 68323
rect 103437 68289 103471 68323
rect 103897 68289 103931 68323
rect 104081 68289 104115 68323
rect 104633 68289 104667 68323
rect 104909 68289 104943 68323
rect 105185 68289 105219 68323
rect 95065 68221 95099 68255
rect 96813 68221 96847 68255
rect 96905 68221 96939 68255
rect 96997 68221 97031 68255
rect 97549 68221 97583 68255
rect 97733 68221 97767 68255
rect 99941 68221 99975 68255
rect 100125 68221 100159 68255
rect 101321 68221 101355 68255
rect 104541 68221 104575 68255
rect 96261 68153 96295 68187
rect 100861 68153 100895 68187
rect 102149 68153 102183 68187
rect 104265 68153 104299 68187
rect 104909 68153 104943 68187
rect 91753 68085 91787 68119
rect 95157 68085 95191 68119
rect 95433 68085 95467 68119
rect 95893 68085 95927 68119
rect 96629 68085 96663 68119
rect 103989 68085 104023 68119
rect 89269 67881 89303 67915
rect 89729 67881 89763 67915
rect 94697 67881 94731 67915
rect 98929 67881 98963 67915
rect 100309 67881 100343 67915
rect 101689 67881 101723 67915
rect 107945 67881 107979 67915
rect 108313 67881 108347 67915
rect 89545 67813 89579 67847
rect 95065 67813 95099 67847
rect 102977 67813 103011 67847
rect 88717 67745 88751 67779
rect 94973 67745 95007 67779
rect 95194 67745 95228 67779
rect 95893 67745 95927 67779
rect 98561 67745 98595 67779
rect 99665 67745 99699 67779
rect 101321 67745 101355 67779
rect 102333 67745 102367 67779
rect 84761 67677 84795 67711
rect 84945 67677 84979 67711
rect 86877 67677 86911 67711
rect 88993 67677 89027 67711
rect 95341 67677 95375 67711
rect 95801 67677 95835 67711
rect 98009 67677 98043 67711
rect 98193 67677 98227 67711
rect 98745 67677 98779 67711
rect 98837 67677 98871 67711
rect 99021 67677 99055 67711
rect 100953 67677 100987 67711
rect 101137 67677 101171 67711
rect 101873 67677 101907 67711
rect 101965 67677 101999 67711
rect 102149 67677 102183 67711
rect 102241 67671 102275 67705
rect 102517 67677 102551 67711
rect 102609 67677 102643 67711
rect 102793 67677 102827 67711
rect 102885 67677 102919 67711
rect 103253 67677 103287 67711
rect 108221 67677 108255 67711
rect 108497 67677 108531 67711
rect 82829 67609 82863 67643
rect 83013 67609 83047 67643
rect 86969 67609 87003 67643
rect 89453 67609 89487 67643
rect 89713 67609 89747 67643
rect 89913 67609 89947 67643
rect 99941 67609 99975 67643
rect 102977 67609 103011 67643
rect 89085 67541 89119 67575
rect 89253 67541 89287 67575
rect 95433 67541 95467 67575
rect 99849 67541 99883 67575
rect 103161 67541 103195 67575
rect 86969 67337 87003 67371
rect 89085 67337 89119 67371
rect 89545 67337 89579 67371
rect 90833 67337 90867 67371
rect 92949 67337 92983 67371
rect 93409 67337 93443 67371
rect 95433 67337 95467 67371
rect 96797 67337 96831 67371
rect 97273 67337 97307 67371
rect 103069 67337 103103 67371
rect 89913 67269 89947 67303
rect 91017 67269 91051 67303
rect 93317 67269 93351 67303
rect 96997 67269 97031 67303
rect 99941 67269 99975 67303
rect 100033 67269 100067 67303
rect 100125 67269 100159 67303
rect 100769 67269 100803 67303
rect 102517 67269 102551 67303
rect 102885 67269 102919 67303
rect 103221 67269 103255 67303
rect 103437 67269 103471 67303
rect 86693 67201 86727 67235
rect 89453 67201 89487 67235
rect 89729 67201 89763 67235
rect 90465 67201 90499 67235
rect 91201 67201 91235 67235
rect 91293 67201 91327 67235
rect 92857 67201 92891 67235
rect 93133 67201 93167 67235
rect 93409 67201 93443 67235
rect 93593 67201 93627 67235
rect 95341 67201 95375 67235
rect 95801 67201 95835 67235
rect 97089 67201 97123 67235
rect 97365 67201 97399 67235
rect 99481 67201 99515 67235
rect 99665 67201 99699 67235
rect 100309 67201 100343 67235
rect 100401 67201 100435 67235
rect 100585 67201 100619 67235
rect 101505 67201 101539 67235
rect 101689 67201 101723 67235
rect 101781 67201 101815 67235
rect 101873 67201 101907 67235
rect 102701 67201 102735 67235
rect 102977 67201 103011 67235
rect 103713 67201 103747 67235
rect 93777 67133 93811 67167
rect 95709 67133 95743 67167
rect 102149 67133 102183 67167
rect 103897 67133 103931 67167
rect 103529 67065 103563 67099
rect 86785 66997 86819 67031
rect 90373 66997 90407 67031
rect 96629 66997 96663 67031
rect 96813 66997 96847 67031
rect 97089 66997 97123 67031
rect 100953 66997 100987 67031
rect 103253 66997 103287 67031
rect 89453 66793 89487 66827
rect 89821 66793 89855 66827
rect 92397 66793 92431 66827
rect 92581 66793 92615 66827
rect 95801 66793 95835 66827
rect 95985 66793 96019 66827
rect 99757 66793 99791 66827
rect 100217 66793 100251 66827
rect 102609 66793 102643 66827
rect 103805 66793 103839 66827
rect 90189 66725 90223 66759
rect 92121 66725 92155 66759
rect 97641 66725 97675 66759
rect 101873 66725 101907 66759
rect 87245 66657 87279 66691
rect 95065 66657 95099 66691
rect 96169 66657 96203 66691
rect 97365 66657 97399 66691
rect 99389 66657 99423 66691
rect 99481 66657 99515 66691
rect 100769 66657 100803 66691
rect 101689 66657 101723 66691
rect 102149 66657 102183 66691
rect 103253 66657 103287 66691
rect 84945 66589 84979 66623
rect 85221 66589 85255 66623
rect 89269 66589 89303 66623
rect 89361 66589 89395 66623
rect 89545 66589 89579 66623
rect 95985 66589 96019 66623
rect 96261 66589 96295 66623
rect 97273 66589 97307 66623
rect 98377 66589 98411 66623
rect 98745 66589 98779 66623
rect 99113 66589 99147 66623
rect 99665 66589 99699 66623
rect 99849 66589 99883 66623
rect 99941 66589 99975 66623
rect 100125 66589 100159 66623
rect 102793 66589 102827 66623
rect 102885 66589 102919 66623
rect 102977 66589 103011 66623
rect 103345 66589 103379 66623
rect 103989 66589 104023 66623
rect 104081 66589 104115 66623
rect 104357 66589 104391 66623
rect 104817 66589 104851 66623
rect 85037 66521 85071 66555
rect 88993 66521 89027 66555
rect 90005 66521 90039 66555
rect 92305 66521 92339 66555
rect 92765 66521 92799 66555
rect 94513 66521 94547 66555
rect 104173 66521 104207 66555
rect 104449 66521 104483 66555
rect 104633 66521 104667 66555
rect 87153 66453 87187 66487
rect 89637 66453 89671 66487
rect 89805 66453 89839 66487
rect 92565 66453 92599 66487
rect 99941 66453 99975 66487
rect 100585 66453 100619 66487
rect 100677 66453 100711 66487
rect 103713 66453 103747 66487
rect 88625 66249 88659 66283
rect 89269 66249 89303 66283
rect 92029 66249 92063 66283
rect 92305 66249 92339 66283
rect 95449 66249 95483 66283
rect 95617 66249 95651 66283
rect 95801 66249 95835 66283
rect 97181 66249 97215 66283
rect 104081 66249 104115 66283
rect 68661 66181 68695 66215
rect 73169 66181 73203 66215
rect 73353 66181 73387 66215
rect 74181 66181 74215 66215
rect 74365 66181 74399 66215
rect 86049 66181 86083 66215
rect 87981 66181 88015 66215
rect 90281 66181 90315 66215
rect 90649 66181 90683 66215
rect 91661 66181 91695 66215
rect 95249 66181 95283 66215
rect 101321 66181 101355 66215
rect 88257 66113 88291 66147
rect 90189 66113 90223 66147
rect 90465 66113 90499 66147
rect 90741 66113 90775 66147
rect 90925 66113 90959 66147
rect 91845 66113 91879 66147
rect 92121 66113 92155 66147
rect 93777 66113 93811 66147
rect 94145 66113 94179 66147
rect 94789 66113 94823 66147
rect 95709 66113 95743 66147
rect 95985 66113 96019 66147
rect 96905 66113 96939 66147
rect 97549 66113 97583 66147
rect 98561 66113 98595 66147
rect 99297 66113 99331 66147
rect 100401 66113 100435 66147
rect 101413 66113 101447 66147
rect 101689 66113 101723 66147
rect 101873 66113 101907 66147
rect 102241 66113 102275 66147
rect 102425 66113 102459 66147
rect 102609 66113 102643 66147
rect 103897 66113 103931 66147
rect 104081 66113 104115 66147
rect 86233 66045 86267 66079
rect 90833 66045 90867 66079
rect 91477 66045 91511 66079
rect 94237 66045 94271 66079
rect 94881 66045 94915 66079
rect 96997 66045 97031 66079
rect 97641 66045 97675 66079
rect 98377 66045 98411 66079
rect 99205 66045 99239 66079
rect 100309 66045 100343 66079
rect 102057 66045 102091 66079
rect 102149 66045 102183 66079
rect 96261 65977 96295 66011
rect 96537 65977 96571 66011
rect 98745 65977 98779 66011
rect 99665 65977 99699 66011
rect 88349 65909 88383 65943
rect 91017 65909 91051 65943
rect 94421 65909 94455 65943
rect 95065 65909 95099 65943
rect 95433 65909 95467 65943
rect 95985 65909 96019 65943
rect 96169 65909 96203 65943
rect 100677 65909 100711 65943
rect 104357 60061 104391 60095
rect 7573 41429 7607 41463
rect 7481 39797 7515 39831
rect 7573 38709 7607 38743
rect 7573 36601 7607 36635
rect 7481 35445 7515 35479
rect 7573 33881 7607 33915
rect 104357 25109 104391 25143
rect 104357 23477 104391 23511
rect 104357 22729 104391 22763
rect 7481 15317 7515 15351
rect 1593 14025 1627 14059
rect 1869 14025 1903 14059
rect 1501 13889 1535 13923
rect 1961 13889 1995 13923
rect 1593 13481 1627 13515
rect 1869 13481 1903 13515
rect 1501 13209 1535 13243
rect 1961 13209 1995 13243
rect 1593 12937 1627 12971
rect 1869 12937 1903 12971
rect 1501 12801 1535 12835
rect 1961 12801 1995 12835
rect 1593 11849 1627 11883
rect 1777 11849 1811 11883
rect 1501 11713 1535 11747
rect 1961 11713 1995 11747
rect 1593 11305 1627 11339
rect 1869 11305 1903 11339
rect 1501 11033 1535 11067
rect 1961 11033 1995 11067
rect 1593 10761 1627 10795
rect 1777 10761 1811 10795
rect 1501 10625 1535 10659
rect 1961 10625 1995 10659
rect 1501 9945 1535 9979
rect 1685 9945 1719 9979
rect 1869 9945 1903 9979
rect 1961 9877 1995 9911
rect 1501 8857 1535 8891
rect 1685 8857 1719 8891
rect 1869 8857 1903 8891
rect 1961 8789 1995 8823
rect 1961 8381 1995 8415
rect 2237 8381 2271 8415
rect 2421 8313 2455 8347
rect 1961 8041 1995 8075
rect 2145 7837 2179 7871
rect 1501 7769 1535 7803
rect 1685 7769 1719 7803
rect 1869 7769 1903 7803
rect 16129 7497 16163 7531
rect 23489 7497 23523 7531
rect 24685 7497 24719 7531
rect 25881 7497 25915 7531
rect 26985 7497 27019 7531
rect 28181 7497 28215 7531
rect 29561 7497 29595 7531
rect 30481 7497 30515 7531
rect 90557 7497 90591 7531
rect 90741 7497 90775 7531
rect 90925 7497 90959 7531
rect 1501 7361 1535 7395
rect 1961 7361 1995 7395
rect 1685 7225 1719 7259
rect 1869 7225 1903 7259
rect 1501 6273 1535 6307
rect 1961 6273 1995 6307
rect 1685 6137 1719 6171
rect 1869 6137 1903 6171
rect 1593 5865 1627 5899
rect 1777 5865 1811 5899
rect 1409 5661 1443 5695
rect 1869 5661 1903 5695
rect 1501 5185 1535 5219
rect 1961 5185 1995 5219
rect 1685 5049 1719 5083
rect 1869 5049 1903 5083
rect 31677 2601 31711 2635
rect 32965 2601 32999 2635
rect 34253 2601 34287 2635
rect 35541 2601 35575 2635
rect 36369 2601 36403 2635
rect 37473 2601 37507 2635
rect 38761 2601 38795 2635
rect 40049 2601 40083 2635
rect 41337 2601 41371 2635
rect 42165 2601 42199 2635
rect 43453 2601 43487 2635
rect 31861 2397 31895 2431
rect 33149 2397 33183 2431
rect 34437 2397 34471 2431
rect 35725 2397 35759 2431
rect 36185 2397 36219 2431
rect 37657 2397 37691 2431
rect 38945 2397 38979 2431
rect 40233 2397 40267 2431
rect 41521 2397 41555 2431
rect 41981 2397 42015 2431
rect 43269 2397 43303 2431
rect 31585 2261 31619 2295
rect 32873 2261 32907 2295
rect 34161 2261 34195 2295
rect 35449 2261 35483 2295
rect 36093 2261 36127 2295
rect 37381 2261 37415 2295
rect 38669 2261 38703 2295
rect 39957 2261 39991 2295
rect 41245 2261 41279 2295
rect 41889 2261 41923 2295
rect 43177 2261 43211 2295
<< metal1 >>
rect 1104 147450 108836 147472
rect 1104 147398 4214 147450
rect 4266 147398 4278 147450
rect 4330 147398 4342 147450
rect 4394 147398 4406 147450
rect 4458 147398 4470 147450
rect 4522 147398 34934 147450
rect 34986 147398 34998 147450
rect 35050 147398 35062 147450
rect 35114 147398 35126 147450
rect 35178 147398 35190 147450
rect 35242 147398 65654 147450
rect 65706 147398 65718 147450
rect 65770 147398 65782 147450
rect 65834 147398 65846 147450
rect 65898 147398 65910 147450
rect 65962 147398 96374 147450
rect 96426 147398 96438 147450
rect 96490 147398 96502 147450
rect 96554 147398 96566 147450
rect 96618 147398 96630 147450
rect 96682 147398 108836 147450
rect 1104 147376 108836 147398
rect 1104 146906 108836 146928
rect 1104 146854 4874 146906
rect 4926 146854 4938 146906
rect 4990 146854 5002 146906
rect 5054 146854 5066 146906
rect 5118 146854 5130 146906
rect 5182 146854 35594 146906
rect 35646 146854 35658 146906
rect 35710 146854 35722 146906
rect 35774 146854 35786 146906
rect 35838 146854 35850 146906
rect 35902 146854 66314 146906
rect 66366 146854 66378 146906
rect 66430 146854 66442 146906
rect 66494 146854 66506 146906
rect 66558 146854 66570 146906
rect 66622 146854 97034 146906
rect 97086 146854 97098 146906
rect 97150 146854 97162 146906
rect 97214 146854 97226 146906
rect 97278 146854 97290 146906
rect 97342 146854 108836 146906
rect 1104 146832 108836 146854
rect 1104 146362 108836 146384
rect 1104 146310 4214 146362
rect 4266 146310 4278 146362
rect 4330 146310 4342 146362
rect 4394 146310 4406 146362
rect 4458 146310 4470 146362
rect 4522 146310 34934 146362
rect 34986 146310 34998 146362
rect 35050 146310 35062 146362
rect 35114 146310 35126 146362
rect 35178 146310 35190 146362
rect 35242 146310 65654 146362
rect 65706 146310 65718 146362
rect 65770 146310 65782 146362
rect 65834 146310 65846 146362
rect 65898 146310 65910 146362
rect 65962 146310 96374 146362
rect 96426 146310 96438 146362
rect 96490 146310 96502 146362
rect 96554 146310 96566 146362
rect 96618 146310 96630 146362
rect 96682 146310 108836 146362
rect 1104 146288 108836 146310
rect 1104 145818 108836 145840
rect 1104 145766 4874 145818
rect 4926 145766 4938 145818
rect 4990 145766 5002 145818
rect 5054 145766 5066 145818
rect 5118 145766 5130 145818
rect 5182 145766 35594 145818
rect 35646 145766 35658 145818
rect 35710 145766 35722 145818
rect 35774 145766 35786 145818
rect 35838 145766 35850 145818
rect 35902 145766 66314 145818
rect 66366 145766 66378 145818
rect 66430 145766 66442 145818
rect 66494 145766 66506 145818
rect 66558 145766 66570 145818
rect 66622 145766 97034 145818
rect 97086 145766 97098 145818
rect 97150 145766 97162 145818
rect 97214 145766 97226 145818
rect 97278 145766 97290 145818
rect 97342 145766 108836 145818
rect 1104 145744 108836 145766
rect 1104 145274 108836 145296
rect 1104 145222 4214 145274
rect 4266 145222 4278 145274
rect 4330 145222 4342 145274
rect 4394 145222 4406 145274
rect 4458 145222 4470 145274
rect 4522 145222 34934 145274
rect 34986 145222 34998 145274
rect 35050 145222 35062 145274
rect 35114 145222 35126 145274
rect 35178 145222 35190 145274
rect 35242 145222 65654 145274
rect 65706 145222 65718 145274
rect 65770 145222 65782 145274
rect 65834 145222 65846 145274
rect 65898 145222 65910 145274
rect 65962 145222 96374 145274
rect 96426 145222 96438 145274
rect 96490 145222 96502 145274
rect 96554 145222 96566 145274
rect 96618 145222 96630 145274
rect 96682 145222 108836 145274
rect 1104 145200 108836 145222
rect 1104 144730 108836 144752
rect 1104 144678 4874 144730
rect 4926 144678 4938 144730
rect 4990 144678 5002 144730
rect 5054 144678 5066 144730
rect 5118 144678 5130 144730
rect 5182 144678 35594 144730
rect 35646 144678 35658 144730
rect 35710 144678 35722 144730
rect 35774 144678 35786 144730
rect 35838 144678 35850 144730
rect 35902 144678 66314 144730
rect 66366 144678 66378 144730
rect 66430 144678 66442 144730
rect 66494 144678 66506 144730
rect 66558 144678 66570 144730
rect 66622 144678 97034 144730
rect 97086 144678 97098 144730
rect 97150 144678 97162 144730
rect 97214 144678 97226 144730
rect 97278 144678 97290 144730
rect 97342 144678 108836 144730
rect 1104 144656 108836 144678
rect 1104 144186 108836 144208
rect 1104 144134 4214 144186
rect 4266 144134 4278 144186
rect 4330 144134 4342 144186
rect 4394 144134 4406 144186
rect 4458 144134 4470 144186
rect 4522 144134 34934 144186
rect 34986 144134 34998 144186
rect 35050 144134 35062 144186
rect 35114 144134 35126 144186
rect 35178 144134 35190 144186
rect 35242 144134 65654 144186
rect 65706 144134 65718 144186
rect 65770 144134 65782 144186
rect 65834 144134 65846 144186
rect 65898 144134 65910 144186
rect 65962 144134 96374 144186
rect 96426 144134 96438 144186
rect 96490 144134 96502 144186
rect 96554 144134 96566 144186
rect 96618 144134 96630 144186
rect 96682 144134 108836 144186
rect 1104 144112 108836 144134
rect 1104 143642 108836 143664
rect 1104 143590 4874 143642
rect 4926 143590 4938 143642
rect 4990 143590 5002 143642
rect 5054 143590 5066 143642
rect 5118 143590 5130 143642
rect 5182 143590 35594 143642
rect 35646 143590 35658 143642
rect 35710 143590 35722 143642
rect 35774 143590 35786 143642
rect 35838 143590 35850 143642
rect 35902 143590 66314 143642
rect 66366 143590 66378 143642
rect 66430 143590 66442 143642
rect 66494 143590 66506 143642
rect 66558 143590 66570 143642
rect 66622 143590 97034 143642
rect 97086 143590 97098 143642
rect 97150 143590 97162 143642
rect 97214 143590 97226 143642
rect 97278 143590 97290 143642
rect 97342 143590 108836 143642
rect 1104 143568 108836 143590
rect 1104 143098 108836 143120
rect 1104 143046 4214 143098
rect 4266 143046 4278 143098
rect 4330 143046 4342 143098
rect 4394 143046 4406 143098
rect 4458 143046 4470 143098
rect 4522 143046 34934 143098
rect 34986 143046 34998 143098
rect 35050 143046 35062 143098
rect 35114 143046 35126 143098
rect 35178 143046 35190 143098
rect 35242 143046 65654 143098
rect 65706 143046 65718 143098
rect 65770 143046 65782 143098
rect 65834 143046 65846 143098
rect 65898 143046 65910 143098
rect 65962 143046 96374 143098
rect 96426 143046 96438 143098
rect 96490 143046 96502 143098
rect 96554 143046 96566 143098
rect 96618 143046 96630 143098
rect 96682 143046 108836 143098
rect 1104 143024 108836 143046
rect 1104 142554 108836 142576
rect 1104 142502 4874 142554
rect 4926 142502 4938 142554
rect 4990 142502 5002 142554
rect 5054 142502 5066 142554
rect 5118 142502 5130 142554
rect 5182 142502 35594 142554
rect 35646 142502 35658 142554
rect 35710 142502 35722 142554
rect 35774 142502 35786 142554
rect 35838 142502 35850 142554
rect 35902 142502 66314 142554
rect 66366 142502 66378 142554
rect 66430 142502 66442 142554
rect 66494 142502 66506 142554
rect 66558 142502 66570 142554
rect 66622 142502 97034 142554
rect 97086 142502 97098 142554
rect 97150 142502 97162 142554
rect 97214 142502 97226 142554
rect 97278 142502 97290 142554
rect 97342 142502 108836 142554
rect 1104 142480 108836 142502
rect 1104 142010 108836 142032
rect 1104 141958 4214 142010
rect 4266 141958 4278 142010
rect 4330 141958 4342 142010
rect 4394 141958 4406 142010
rect 4458 141958 4470 142010
rect 4522 141958 34934 142010
rect 34986 141958 34998 142010
rect 35050 141958 35062 142010
rect 35114 141958 35126 142010
rect 35178 141958 35190 142010
rect 35242 141958 65654 142010
rect 65706 141958 65718 142010
rect 65770 141958 65782 142010
rect 65834 141958 65846 142010
rect 65898 141958 65910 142010
rect 65962 141958 96374 142010
rect 96426 141958 96438 142010
rect 96490 141958 96502 142010
rect 96554 141958 96566 142010
rect 96618 141958 96630 142010
rect 96682 141958 108836 142010
rect 1104 141936 108836 141958
rect 1104 141466 108836 141488
rect 1104 141414 4874 141466
rect 4926 141414 4938 141466
rect 4990 141414 5002 141466
rect 5054 141414 5066 141466
rect 5118 141414 5130 141466
rect 5182 141414 35594 141466
rect 35646 141414 35658 141466
rect 35710 141414 35722 141466
rect 35774 141414 35786 141466
rect 35838 141414 35850 141466
rect 35902 141414 66314 141466
rect 66366 141414 66378 141466
rect 66430 141414 66442 141466
rect 66494 141414 66506 141466
rect 66558 141414 66570 141466
rect 66622 141414 97034 141466
rect 97086 141414 97098 141466
rect 97150 141414 97162 141466
rect 97214 141414 97226 141466
rect 97278 141414 97290 141466
rect 97342 141414 108836 141466
rect 1104 141392 108836 141414
rect 1104 140922 108836 140944
rect 1104 140870 4214 140922
rect 4266 140870 4278 140922
rect 4330 140870 4342 140922
rect 4394 140870 4406 140922
rect 4458 140870 4470 140922
rect 4522 140870 34934 140922
rect 34986 140870 34998 140922
rect 35050 140870 35062 140922
rect 35114 140870 35126 140922
rect 35178 140870 35190 140922
rect 35242 140870 65654 140922
rect 65706 140870 65718 140922
rect 65770 140870 65782 140922
rect 65834 140870 65846 140922
rect 65898 140870 65910 140922
rect 65962 140870 96374 140922
rect 96426 140870 96438 140922
rect 96490 140870 96502 140922
rect 96554 140870 96566 140922
rect 96618 140870 96630 140922
rect 96682 140870 108836 140922
rect 1104 140848 108836 140870
rect 1104 140378 108836 140400
rect 1104 140326 4874 140378
rect 4926 140326 4938 140378
rect 4990 140326 5002 140378
rect 5054 140326 5066 140378
rect 5118 140326 5130 140378
rect 5182 140326 35594 140378
rect 35646 140326 35658 140378
rect 35710 140326 35722 140378
rect 35774 140326 35786 140378
rect 35838 140326 35850 140378
rect 35902 140326 66314 140378
rect 66366 140326 66378 140378
rect 66430 140326 66442 140378
rect 66494 140326 66506 140378
rect 66558 140326 66570 140378
rect 66622 140326 97034 140378
rect 97086 140326 97098 140378
rect 97150 140326 97162 140378
rect 97214 140326 97226 140378
rect 97278 140326 97290 140378
rect 97342 140326 108836 140378
rect 1104 140304 108836 140326
rect 1104 139834 108836 139856
rect 1104 139782 4214 139834
rect 4266 139782 4278 139834
rect 4330 139782 4342 139834
rect 4394 139782 4406 139834
rect 4458 139782 4470 139834
rect 4522 139782 34934 139834
rect 34986 139782 34998 139834
rect 35050 139782 35062 139834
rect 35114 139782 35126 139834
rect 35178 139782 35190 139834
rect 35242 139782 65654 139834
rect 65706 139782 65718 139834
rect 65770 139782 65782 139834
rect 65834 139782 65846 139834
rect 65898 139782 65910 139834
rect 65962 139782 96374 139834
rect 96426 139782 96438 139834
rect 96490 139782 96502 139834
rect 96554 139782 96566 139834
rect 96618 139782 96630 139834
rect 96682 139782 108836 139834
rect 1104 139760 108836 139782
rect 1104 139290 108836 139312
rect 1104 139238 4874 139290
rect 4926 139238 4938 139290
rect 4990 139238 5002 139290
rect 5054 139238 5066 139290
rect 5118 139238 5130 139290
rect 5182 139238 35594 139290
rect 35646 139238 35658 139290
rect 35710 139238 35722 139290
rect 35774 139238 35786 139290
rect 35838 139238 35850 139290
rect 35902 139238 66314 139290
rect 66366 139238 66378 139290
rect 66430 139238 66442 139290
rect 66494 139238 66506 139290
rect 66558 139238 66570 139290
rect 66622 139238 97034 139290
rect 97086 139238 97098 139290
rect 97150 139238 97162 139290
rect 97214 139238 97226 139290
rect 97278 139238 97290 139290
rect 97342 139238 108836 139290
rect 1104 139216 108836 139238
rect 1104 138746 108836 138768
rect 1104 138694 4214 138746
rect 4266 138694 4278 138746
rect 4330 138694 4342 138746
rect 4394 138694 4406 138746
rect 4458 138694 4470 138746
rect 4522 138694 34934 138746
rect 34986 138694 34998 138746
rect 35050 138694 35062 138746
rect 35114 138694 35126 138746
rect 35178 138694 35190 138746
rect 35242 138694 65654 138746
rect 65706 138694 65718 138746
rect 65770 138694 65782 138746
rect 65834 138694 65846 138746
rect 65898 138694 65910 138746
rect 65962 138694 96374 138746
rect 96426 138694 96438 138746
rect 96490 138694 96502 138746
rect 96554 138694 96566 138746
rect 96618 138694 96630 138746
rect 96682 138694 108836 138746
rect 1104 138672 108836 138694
rect 1104 138202 108836 138224
rect 1104 138150 4874 138202
rect 4926 138150 4938 138202
rect 4990 138150 5002 138202
rect 5054 138150 5066 138202
rect 5118 138150 5130 138202
rect 5182 138150 35594 138202
rect 35646 138150 35658 138202
rect 35710 138150 35722 138202
rect 35774 138150 35786 138202
rect 35838 138150 35850 138202
rect 35902 138150 66314 138202
rect 66366 138150 66378 138202
rect 66430 138150 66442 138202
rect 66494 138150 66506 138202
rect 66558 138150 66570 138202
rect 66622 138150 97034 138202
rect 97086 138150 97098 138202
rect 97150 138150 97162 138202
rect 97214 138150 97226 138202
rect 97278 138150 97290 138202
rect 97342 138150 108836 138202
rect 1104 138128 108836 138150
rect 1104 137658 108836 137680
rect 1104 137606 4214 137658
rect 4266 137606 4278 137658
rect 4330 137606 4342 137658
rect 4394 137606 4406 137658
rect 4458 137606 4470 137658
rect 4522 137606 34934 137658
rect 34986 137606 34998 137658
rect 35050 137606 35062 137658
rect 35114 137606 35126 137658
rect 35178 137606 35190 137658
rect 35242 137606 65654 137658
rect 65706 137606 65718 137658
rect 65770 137606 65782 137658
rect 65834 137606 65846 137658
rect 65898 137606 65910 137658
rect 65962 137606 96374 137658
rect 96426 137606 96438 137658
rect 96490 137606 96502 137658
rect 96554 137606 96566 137658
rect 96618 137606 96630 137658
rect 96682 137606 108836 137658
rect 1104 137584 108836 137606
rect 1104 137114 108836 137136
rect 1104 137062 4874 137114
rect 4926 137062 4938 137114
rect 4990 137062 5002 137114
rect 5054 137062 5066 137114
rect 5118 137062 5130 137114
rect 5182 137062 35594 137114
rect 35646 137062 35658 137114
rect 35710 137062 35722 137114
rect 35774 137062 35786 137114
rect 35838 137062 35850 137114
rect 35902 137062 66314 137114
rect 66366 137062 66378 137114
rect 66430 137062 66442 137114
rect 66494 137062 66506 137114
rect 66558 137062 66570 137114
rect 66622 137062 97034 137114
rect 97086 137062 97098 137114
rect 97150 137062 97162 137114
rect 97214 137062 97226 137114
rect 97278 137062 97290 137114
rect 97342 137062 108836 137114
rect 1104 137040 108836 137062
rect 85485 137003 85543 137009
rect 85485 137000 85497 137003
rect 85224 136972 85497 137000
rect 85034 136867 85092 136873
rect 85034 136864 85046 136867
rect 83660 136836 85046 136864
rect 63586 136620 63592 136672
rect 63644 136660 63650 136672
rect 83660 136669 83688 136836
rect 85034 136833 85046 136836
rect 85080 136833 85092 136867
rect 85034 136827 85092 136833
rect 85224 136796 85252 136972
rect 85485 136969 85497 136972
rect 85531 137000 85543 137003
rect 85531 136972 93854 137000
rect 85531 136969 85543 136972
rect 85485 136963 85543 136969
rect 85316 136904 85712 136932
rect 85316 136873 85344 136904
rect 85301 136867 85359 136873
rect 85301 136833 85313 136867
rect 85347 136833 85359 136867
rect 85301 136827 85359 136833
rect 85224 136768 85344 136796
rect 83645 136663 83703 136669
rect 83645 136660 83657 136663
rect 63644 136632 83657 136660
rect 63644 136620 63650 136632
rect 83645 136629 83657 136632
rect 83691 136629 83703 136663
rect 83645 136623 83703 136629
rect 83921 136663 83979 136669
rect 83921 136629 83933 136663
rect 83967 136660 83979 136663
rect 85316 136660 85344 136768
rect 85684 136669 85712 136904
rect 93826 136864 93854 136972
rect 102134 136864 102140 136876
rect 93826 136836 102140 136864
rect 102134 136824 102140 136836
rect 102192 136824 102198 136876
rect 83967 136632 85344 136660
rect 85669 136663 85727 136669
rect 83967 136629 83979 136632
rect 83921 136623 83979 136629
rect 85669 136629 85681 136663
rect 85715 136660 85727 136663
rect 95970 136660 95976 136672
rect 85715 136632 95976 136660
rect 85715 136629 85727 136632
rect 85669 136623 85727 136629
rect 95970 136620 95976 136632
rect 96028 136620 96034 136672
rect 1104 136570 108836 136592
rect 1104 136518 4214 136570
rect 4266 136518 4278 136570
rect 4330 136518 4342 136570
rect 4394 136518 4406 136570
rect 4458 136518 4470 136570
rect 4522 136518 34934 136570
rect 34986 136518 34998 136570
rect 35050 136518 35062 136570
rect 35114 136518 35126 136570
rect 35178 136518 35190 136570
rect 35242 136518 65654 136570
rect 65706 136518 65718 136570
rect 65770 136518 65782 136570
rect 65834 136518 65846 136570
rect 65898 136518 65910 136570
rect 65962 136518 96374 136570
rect 96426 136518 96438 136570
rect 96490 136518 96502 136570
rect 96554 136518 96566 136570
rect 96618 136518 96630 136570
rect 96682 136518 105922 136570
rect 105974 136518 105986 136570
rect 106038 136518 106050 136570
rect 106102 136518 106114 136570
rect 106166 136518 106178 136570
rect 106230 136518 108836 136570
rect 1104 136496 108836 136518
rect 34333 136255 34391 136261
rect 34333 136221 34345 136255
rect 34379 136252 34391 136255
rect 35986 136252 35992 136264
rect 34379 136224 35992 136252
rect 34379 136221 34391 136224
rect 34333 136215 34391 136221
rect 35986 136212 35992 136224
rect 36044 136212 36050 136264
rect 38562 136252 38568 136264
rect 36096 136224 38568 136252
rect 34146 136144 34152 136196
rect 34204 136184 34210 136196
rect 34701 136187 34759 136193
rect 34701 136184 34713 136187
rect 34204 136156 34713 136184
rect 34204 136144 34210 136156
rect 34701 136153 34713 136156
rect 34747 136153 34759 136187
rect 34701 136147 34759 136153
rect 34974 136144 34980 136196
rect 35032 136144 35038 136196
rect 35161 136187 35219 136193
rect 35161 136153 35173 136187
rect 35207 136184 35219 136187
rect 36096 136184 36124 136224
rect 38562 136212 38568 136224
rect 38620 136212 38626 136264
rect 35207 136156 36124 136184
rect 36173 136187 36231 136193
rect 35207 136153 35219 136156
rect 35161 136147 35219 136153
rect 36173 136153 36185 136187
rect 36219 136184 36231 136187
rect 38746 136184 38752 136196
rect 36219 136156 38752 136184
rect 36219 136153 36231 136156
rect 36173 136147 36231 136153
rect 38746 136144 38752 136156
rect 38804 136144 38810 136196
rect 43162 136144 43168 136196
rect 43220 136144 43226 136196
rect 47765 136187 47823 136193
rect 47765 136153 47777 136187
rect 47811 136184 47823 136187
rect 48498 136184 48504 136196
rect 47811 136156 48504 136184
rect 47811 136153 47823 136156
rect 47765 136147 47823 136153
rect 48498 136144 48504 136156
rect 48556 136144 48562 136196
rect 50341 136187 50399 136193
rect 50341 136153 50353 136187
rect 50387 136184 50399 136187
rect 51074 136184 51080 136196
rect 50387 136156 51080 136184
rect 50387 136153 50399 136156
rect 50341 136147 50399 136153
rect 51074 136144 51080 136156
rect 51132 136144 51138 136196
rect 55398 136144 55404 136196
rect 55456 136144 55462 136196
rect 57974 136144 57980 136196
rect 58032 136144 58038 136196
rect 60550 136144 60556 136196
rect 60608 136144 60614 136196
rect 60737 136187 60795 136193
rect 60737 136153 60749 136187
rect 60783 136153 60795 136187
rect 60737 136147 60795 136153
rect 34992 136116 35020 136144
rect 35345 136119 35403 136125
rect 35345 136116 35357 136119
rect 34992 136088 35357 136116
rect 35345 136085 35357 136088
rect 35391 136085 35403 136119
rect 35345 136079 35403 136085
rect 36078 136076 36084 136128
rect 36136 136116 36142 136128
rect 36357 136119 36415 136125
rect 36357 136116 36369 136119
rect 36136 136088 36369 136116
rect 36136 136076 36142 136088
rect 36357 136085 36369 136088
rect 36403 136085 36415 136119
rect 36357 136079 36415 136085
rect 43070 136076 43076 136128
rect 43128 136116 43134 136128
rect 43349 136119 43407 136125
rect 43349 136116 43361 136119
rect 43128 136088 43361 136116
rect 43128 136076 43134 136088
rect 43349 136085 43361 136088
rect 43395 136085 43407 136119
rect 43349 136079 43407 136085
rect 46106 136076 46112 136128
rect 46164 136076 46170 136128
rect 47670 136076 47676 136128
rect 47728 136116 47734 136128
rect 47949 136119 48007 136125
rect 47949 136116 47961 136119
rect 47728 136088 47961 136116
rect 47728 136076 47734 136088
rect 47949 136085 47961 136088
rect 47995 136085 48007 136119
rect 47949 136079 48007 136085
rect 50246 136076 50252 136128
rect 50304 136116 50310 136128
rect 50525 136119 50583 136125
rect 50525 136116 50537 136119
rect 50304 136088 50537 136116
rect 50304 136076 50310 136088
rect 50525 136085 50537 136088
rect 50571 136085 50583 136119
rect 50525 136079 50583 136085
rect 55493 136119 55551 136125
rect 55493 136085 55505 136119
rect 55539 136116 55551 136119
rect 55766 136116 55772 136128
rect 55539 136088 55772 136116
rect 55539 136085 55551 136088
rect 55493 136079 55551 136085
rect 55766 136076 55772 136088
rect 55824 136076 55830 136128
rect 58069 136119 58127 136125
rect 58069 136085 58081 136119
rect 58115 136116 58127 136119
rect 58342 136116 58348 136128
rect 58115 136088 58348 136116
rect 58115 136085 58127 136088
rect 58069 136079 58127 136085
rect 58342 136076 58348 136088
rect 58400 136076 58406 136128
rect 60752 136116 60780 136147
rect 63126 136144 63132 136196
rect 63184 136144 63190 136196
rect 72510 136144 72516 136196
rect 72568 136144 72574 136196
rect 72694 136144 72700 136196
rect 72752 136184 72758 136196
rect 73433 136187 73491 136193
rect 73433 136184 73445 136187
rect 72752 136156 73445 136184
rect 72752 136144 72758 136156
rect 73433 136153 73445 136156
rect 73479 136153 73491 136187
rect 73433 136147 73491 136153
rect 77386 136144 77392 136196
rect 77444 136144 77450 136196
rect 60918 136116 60924 136128
rect 60752 136088 60924 136116
rect 60918 136076 60924 136088
rect 60976 136076 60982 136128
rect 63221 136119 63279 136125
rect 63221 136085 63233 136119
rect 63267 136116 63279 136119
rect 63494 136116 63500 136128
rect 63267 136088 63500 136116
rect 63267 136085 63279 136088
rect 63221 136079 63279 136085
rect 63494 136076 63500 136088
rect 63552 136076 63558 136128
rect 63586 136076 63592 136128
rect 63644 136076 63650 136128
rect 68554 136076 68560 136128
rect 68612 136076 68618 136128
rect 72605 136119 72663 136125
rect 72605 136085 72617 136119
rect 72651 136116 72663 136119
rect 72878 136116 72884 136128
rect 72651 136088 72884 136116
rect 72651 136085 72663 136088
rect 72605 136079 72663 136085
rect 72878 136076 72884 136088
rect 72936 136076 72942 136128
rect 73525 136119 73583 136125
rect 73525 136085 73537 136119
rect 73571 136116 73583 136119
rect 73798 136116 73804 136128
rect 73571 136088 73804 136116
rect 73571 136085 73583 136088
rect 73525 136079 73583 136085
rect 73798 136076 73804 136088
rect 73856 136076 73862 136128
rect 77481 136119 77539 136125
rect 77481 136085 77493 136119
rect 77527 136116 77539 136119
rect 77754 136116 77760 136128
rect 77527 136088 77760 136116
rect 77527 136085 77539 136088
rect 77481 136079 77539 136085
rect 77754 136076 77760 136088
rect 77812 136076 77818 136128
rect 86310 136076 86316 136128
rect 86368 136076 86374 136128
rect 87322 136076 87328 136128
rect 87380 136076 87386 136128
rect 95970 136076 95976 136128
rect 96028 136116 96034 136128
rect 104342 136116 104348 136128
rect 96028 136088 104348 136116
rect 96028 136076 96034 136088
rect 104342 136076 104348 136088
rect 104400 136076 104406 136128
rect 1104 136026 108836 136048
rect 1104 135974 4874 136026
rect 4926 135974 4938 136026
rect 4990 135974 5002 136026
rect 5054 135974 5066 136026
rect 5118 135974 5130 136026
rect 5182 135974 35594 136026
rect 35646 135974 35658 136026
rect 35710 135974 35722 136026
rect 35774 135974 35786 136026
rect 35838 135974 35850 136026
rect 35902 135974 66314 136026
rect 66366 135974 66378 136026
rect 66430 135974 66442 136026
rect 66494 135974 66506 136026
rect 66558 135974 66570 136026
rect 66622 135974 97034 136026
rect 97086 135974 97098 136026
rect 97150 135974 97162 136026
rect 97214 135974 97226 136026
rect 97278 135974 97290 136026
rect 97342 135974 106658 136026
rect 106710 135974 106722 136026
rect 106774 135974 106786 136026
rect 106838 135974 106850 136026
rect 106902 135974 106914 136026
rect 106966 135974 108836 136026
rect 1104 135952 108836 135974
rect 9582 135872 9588 135924
rect 9640 135912 9646 135924
rect 47670 135912 47676 135924
rect 9640 135884 47676 135912
rect 9640 135872 9646 135884
rect 47670 135872 47676 135884
rect 47728 135872 47734 135924
rect 55766 135872 55772 135924
rect 55824 135912 55830 135924
rect 103698 135912 103704 135924
rect 55824 135884 103704 135912
rect 55824 135872 55830 135884
rect 103698 135872 103704 135884
rect 103756 135872 103762 135924
rect 8202 135804 8208 135856
rect 8260 135844 8266 135856
rect 43070 135844 43076 135856
rect 8260 135816 43076 135844
rect 8260 135804 8266 135816
rect 43070 135804 43076 135816
rect 43128 135804 43134 135856
rect 58342 135804 58348 135856
rect 58400 135844 58406 135856
rect 102226 135844 102232 135856
rect 58400 135816 102232 135844
rect 58400 135804 58406 135816
rect 102226 135804 102232 135816
rect 102284 135804 102290 135856
rect 8018 135736 8024 135788
rect 8076 135776 8082 135788
rect 36078 135776 36084 135788
rect 8076 135748 36084 135776
rect 8076 135736 8082 135748
rect 36078 135736 36084 135748
rect 36136 135736 36142 135788
rect 60918 135736 60924 135788
rect 60976 135776 60982 135788
rect 103790 135776 103796 135788
rect 60976 135748 103796 135776
rect 60976 135736 60982 135748
rect 103790 135736 103796 135748
rect 103848 135736 103854 135788
rect 63494 135668 63500 135720
rect 63552 135708 63558 135720
rect 103606 135708 103612 135720
rect 63552 135680 103612 135708
rect 63552 135668 63558 135680
rect 103606 135668 103612 135680
rect 103664 135668 103670 135720
rect 72878 135600 72884 135652
rect 72936 135640 72942 135652
rect 103514 135640 103520 135652
rect 72936 135612 103520 135640
rect 72936 135600 72942 135612
rect 103514 135600 103520 135612
rect 103572 135600 103578 135652
rect 8110 135532 8116 135584
rect 8168 135572 8174 135584
rect 50246 135572 50252 135584
rect 8168 135544 50252 135572
rect 8168 135532 8174 135544
rect 50246 135532 50252 135544
rect 50304 135532 50310 135584
rect 73798 135532 73804 135584
rect 73856 135572 73862 135584
rect 104618 135572 104624 135584
rect 73856 135544 104624 135572
rect 73856 135532 73862 135544
rect 104618 135532 104624 135544
rect 104676 135532 104682 135584
rect 1104 135482 7912 135504
rect 1104 135430 4214 135482
rect 4266 135430 4278 135482
rect 4330 135430 4342 135482
rect 4394 135430 4406 135482
rect 4458 135430 4470 135482
rect 4522 135430 7912 135482
rect 77754 135464 77760 135516
rect 77812 135504 77818 135516
rect 102778 135504 102784 135516
rect 77812 135476 102784 135504
rect 77812 135464 77818 135476
rect 102778 135464 102784 135476
rect 102836 135464 102842 135516
rect 104052 135482 108836 135504
rect 1104 135408 7912 135430
rect 86310 135396 86316 135448
rect 86368 135436 86374 135448
rect 102318 135436 102324 135448
rect 86368 135408 102324 135436
rect 86368 135396 86374 135408
rect 102318 135396 102324 135408
rect 102376 135396 102382 135448
rect 104052 135430 105922 135482
rect 105974 135430 105986 135482
rect 106038 135430 106050 135482
rect 106102 135430 106114 135482
rect 106166 135430 106178 135482
rect 106230 135430 108836 135482
rect 104052 135408 108836 135430
rect 1104 134938 7912 134960
rect 1104 134886 4874 134938
rect 4926 134886 4938 134938
rect 4990 134886 5002 134938
rect 5054 134886 5066 134938
rect 5118 134886 5130 134938
rect 5182 134886 7912 134938
rect 1104 134864 7912 134886
rect 104052 134938 108836 134960
rect 104052 134886 106658 134938
rect 106710 134886 106722 134938
rect 106774 134886 106786 134938
rect 106838 134886 106850 134938
rect 106902 134886 106914 134938
rect 106966 134886 108836 134938
rect 104052 134864 108836 134886
rect 8938 134580 8944 134632
rect 8996 134620 9002 134632
rect 34146 134620 34152 134632
rect 8996 134592 34152 134620
rect 8996 134580 9002 134592
rect 34146 134580 34152 134592
rect 34204 134580 34210 134632
rect 9030 134512 9036 134564
rect 9088 134552 9094 134564
rect 34974 134552 34980 134564
rect 9088 134524 34980 134552
rect 9088 134512 9094 134524
rect 34974 134512 34980 134524
rect 35032 134512 35038 134564
rect 1104 134394 7912 134416
rect 1104 134342 4214 134394
rect 4266 134342 4278 134394
rect 4330 134342 4342 134394
rect 4394 134342 4406 134394
rect 4458 134342 4470 134394
rect 4522 134342 7912 134394
rect 1104 134320 7912 134342
rect 104052 134394 108836 134416
rect 104052 134342 105922 134394
rect 105974 134342 105986 134394
rect 106038 134342 106050 134394
rect 106102 134342 106114 134394
rect 106166 134342 106178 134394
rect 106230 134342 108836 134394
rect 104052 134320 108836 134342
rect 87322 133900 87328 133952
rect 87380 133940 87386 133952
rect 104066 133940 104072 133952
rect 87380 133912 104072 133940
rect 87380 133900 87386 133912
rect 104066 133900 104072 133912
rect 104124 133900 104130 133952
rect 1104 133850 7912 133872
rect 1104 133798 4874 133850
rect 4926 133798 4938 133850
rect 4990 133798 5002 133850
rect 5054 133798 5066 133850
rect 5118 133798 5130 133850
rect 5182 133798 7912 133850
rect 1104 133776 7912 133798
rect 104052 133850 108836 133872
rect 104052 133798 106658 133850
rect 106710 133798 106722 133850
rect 106774 133798 106786 133850
rect 106838 133798 106850 133850
rect 106902 133798 106914 133850
rect 106966 133798 108836 133850
rect 104052 133776 108836 133798
rect 7374 133696 7380 133748
rect 7432 133736 7438 133748
rect 46106 133736 46112 133748
rect 7432 133708 46112 133736
rect 7432 133696 7438 133708
rect 46106 133696 46112 133708
rect 46164 133696 46170 133748
rect 68554 133696 68560 133748
rect 68612 133736 68618 133748
rect 104526 133736 104532 133748
rect 68612 133708 104532 133736
rect 68612 133696 68618 133708
rect 104526 133696 104532 133708
rect 104584 133696 104590 133748
rect 1104 133306 7912 133328
rect 1104 133254 4214 133306
rect 4266 133254 4278 133306
rect 4330 133254 4342 133306
rect 4394 133254 4406 133306
rect 4458 133254 4470 133306
rect 4522 133254 7912 133306
rect 1104 133232 7912 133254
rect 104052 133306 108836 133328
rect 104052 133254 105922 133306
rect 105974 133254 105986 133306
rect 106038 133254 106050 133306
rect 106102 133254 106114 133306
rect 106166 133254 106178 133306
rect 106230 133254 108836 133306
rect 104052 133232 108836 133254
rect 1104 132762 7912 132784
rect 1104 132710 4874 132762
rect 4926 132710 4938 132762
rect 4990 132710 5002 132762
rect 5054 132710 5066 132762
rect 5118 132710 5130 132762
rect 5182 132710 7912 132762
rect 1104 132688 7912 132710
rect 104052 132762 108836 132784
rect 104052 132710 106658 132762
rect 106710 132710 106722 132762
rect 106774 132710 106786 132762
rect 106838 132710 106850 132762
rect 106902 132710 106914 132762
rect 106966 132710 108836 132762
rect 104052 132688 108836 132710
rect 1104 132218 7912 132240
rect 1104 132166 4214 132218
rect 4266 132166 4278 132218
rect 4330 132166 4342 132218
rect 4394 132166 4406 132218
rect 4458 132166 4470 132218
rect 4522 132166 7912 132218
rect 1104 132144 7912 132166
rect 104052 132218 108836 132240
rect 104052 132166 105922 132218
rect 105974 132166 105986 132218
rect 106038 132166 106050 132218
rect 106102 132166 106114 132218
rect 106166 132166 106178 132218
rect 106230 132166 108836 132218
rect 104052 132144 108836 132166
rect 1104 131674 7912 131696
rect 1104 131622 4874 131674
rect 4926 131622 4938 131674
rect 4990 131622 5002 131674
rect 5054 131622 5066 131674
rect 5118 131622 5130 131674
rect 5182 131622 7912 131674
rect 1104 131600 7912 131622
rect 104052 131674 108836 131696
rect 104052 131622 106658 131674
rect 106710 131622 106722 131674
rect 106774 131622 106786 131674
rect 106838 131622 106850 131674
rect 106902 131622 106914 131674
rect 106966 131622 108836 131674
rect 104052 131600 108836 131622
rect 1104 131130 7912 131152
rect 1104 131078 4214 131130
rect 4266 131078 4278 131130
rect 4330 131078 4342 131130
rect 4394 131078 4406 131130
rect 4458 131078 4470 131130
rect 4522 131078 7912 131130
rect 1104 131056 7912 131078
rect 104052 131130 108836 131152
rect 104052 131078 105922 131130
rect 105974 131078 105986 131130
rect 106038 131078 106050 131130
rect 106102 131078 106114 131130
rect 106166 131078 106178 131130
rect 106230 131078 108836 131130
rect 104052 131056 108836 131078
rect 1104 130586 7912 130608
rect 1104 130534 4874 130586
rect 4926 130534 4938 130586
rect 4990 130534 5002 130586
rect 5054 130534 5066 130586
rect 5118 130534 5130 130586
rect 5182 130534 7912 130586
rect 1104 130512 7912 130534
rect 104052 130586 108836 130608
rect 104052 130534 106658 130586
rect 106710 130534 106722 130586
rect 106774 130534 106786 130586
rect 106838 130534 106850 130586
rect 106902 130534 106914 130586
rect 106966 130534 108836 130586
rect 104052 130512 108836 130534
rect 1104 130042 7912 130064
rect 1104 129990 4214 130042
rect 4266 129990 4278 130042
rect 4330 129990 4342 130042
rect 4394 129990 4406 130042
rect 4458 129990 4470 130042
rect 4522 129990 7912 130042
rect 1104 129968 7912 129990
rect 104052 130042 108836 130064
rect 104052 129990 105922 130042
rect 105974 129990 105986 130042
rect 106038 129990 106050 130042
rect 106102 129990 106114 130042
rect 106166 129990 106178 130042
rect 106230 129990 108836 130042
rect 104052 129968 108836 129990
rect 103882 129752 103888 129804
rect 103940 129792 103946 129804
rect 104345 129795 104403 129801
rect 104345 129792 104357 129795
rect 103940 129764 104357 129792
rect 103940 129752 103946 129764
rect 104345 129761 104357 129764
rect 104391 129761 104403 129795
rect 104345 129755 104403 129761
rect 1104 129498 7912 129520
rect 1104 129446 4874 129498
rect 4926 129446 4938 129498
rect 4990 129446 5002 129498
rect 5054 129446 5066 129498
rect 5118 129446 5130 129498
rect 5182 129446 7912 129498
rect 1104 129424 7912 129446
rect 104052 129498 108836 129520
rect 104052 129446 106658 129498
rect 106710 129446 106722 129498
rect 106774 129446 106786 129498
rect 106838 129446 106850 129498
rect 106902 129446 106914 129498
rect 106966 129446 108836 129498
rect 104052 129424 108836 129446
rect 1104 128954 7912 128976
rect 1104 128902 4214 128954
rect 4266 128902 4278 128954
rect 4330 128902 4342 128954
rect 4394 128902 4406 128954
rect 4458 128902 4470 128954
rect 4522 128902 7912 128954
rect 1104 128880 7912 128902
rect 104052 128954 108836 128976
rect 104052 128902 105922 128954
rect 105974 128902 105986 128954
rect 106038 128902 106050 128954
rect 106102 128902 106114 128954
rect 106166 128902 106178 128954
rect 106230 128902 108836 128954
rect 104052 128880 108836 128902
rect 1104 128410 7912 128432
rect 1104 128358 4874 128410
rect 4926 128358 4938 128410
rect 4990 128358 5002 128410
rect 5054 128358 5066 128410
rect 5118 128358 5130 128410
rect 5182 128358 7912 128410
rect 1104 128336 7912 128358
rect 104052 128410 108836 128432
rect 104052 128358 106658 128410
rect 106710 128358 106722 128410
rect 106774 128358 106786 128410
rect 106838 128358 106850 128410
rect 106902 128358 106914 128410
rect 106966 128358 108836 128410
rect 104052 128336 108836 128358
rect 1104 127866 7912 127888
rect 1104 127814 4214 127866
rect 4266 127814 4278 127866
rect 4330 127814 4342 127866
rect 4394 127814 4406 127866
rect 4458 127814 4470 127866
rect 4522 127814 7912 127866
rect 1104 127792 7912 127814
rect 104052 127866 108836 127888
rect 104052 127814 105922 127866
rect 105974 127814 105986 127866
rect 106038 127814 106050 127866
rect 106102 127814 106114 127866
rect 106166 127814 106178 127866
rect 106230 127814 108836 127866
rect 104052 127792 108836 127814
rect 1104 127322 7912 127344
rect 1104 127270 4874 127322
rect 4926 127270 4938 127322
rect 4990 127270 5002 127322
rect 5054 127270 5066 127322
rect 5118 127270 5130 127322
rect 5182 127270 7912 127322
rect 1104 127248 7912 127270
rect 104052 127322 108836 127344
rect 104052 127270 106658 127322
rect 106710 127270 106722 127322
rect 106774 127270 106786 127322
rect 106838 127270 106850 127322
rect 106902 127270 106914 127322
rect 106966 127270 108836 127322
rect 104052 127248 108836 127270
rect 1104 126778 7912 126800
rect 1104 126726 4214 126778
rect 4266 126726 4278 126778
rect 4330 126726 4342 126778
rect 4394 126726 4406 126778
rect 4458 126726 4470 126778
rect 4522 126726 7912 126778
rect 1104 126704 7912 126726
rect 104052 126778 108836 126800
rect 104052 126726 105922 126778
rect 105974 126726 105986 126778
rect 106038 126726 106050 126778
rect 106102 126726 106114 126778
rect 106166 126726 106178 126778
rect 106230 126726 108836 126778
rect 104052 126704 108836 126726
rect 1104 126234 7912 126256
rect 1104 126182 4874 126234
rect 4926 126182 4938 126234
rect 4990 126182 5002 126234
rect 5054 126182 5066 126234
rect 5118 126182 5130 126234
rect 5182 126182 7912 126234
rect 1104 126160 7912 126182
rect 104052 126234 108836 126256
rect 104052 126182 106658 126234
rect 106710 126182 106722 126234
rect 106774 126182 106786 126234
rect 106838 126182 106850 126234
rect 106902 126182 106914 126234
rect 106966 126182 108836 126234
rect 104052 126160 108836 126182
rect 1104 125690 7912 125712
rect 1104 125638 4214 125690
rect 4266 125638 4278 125690
rect 4330 125638 4342 125690
rect 4394 125638 4406 125690
rect 4458 125638 4470 125690
rect 4522 125638 7912 125690
rect 1104 125616 7912 125638
rect 104052 125690 108836 125712
rect 104052 125638 105922 125690
rect 105974 125638 105986 125690
rect 106038 125638 106050 125690
rect 106102 125638 106114 125690
rect 106166 125638 106178 125690
rect 106230 125638 108836 125690
rect 104052 125616 108836 125638
rect 1104 125146 7912 125168
rect 1104 125094 4874 125146
rect 4926 125094 4938 125146
rect 4990 125094 5002 125146
rect 5054 125094 5066 125146
rect 5118 125094 5130 125146
rect 5182 125094 7912 125146
rect 1104 125072 7912 125094
rect 104052 125146 108836 125168
rect 104052 125094 106658 125146
rect 106710 125094 106722 125146
rect 106774 125094 106786 125146
rect 106838 125094 106850 125146
rect 106902 125094 106914 125146
rect 106966 125094 108836 125146
rect 104052 125072 108836 125094
rect 1104 124602 7912 124624
rect 1104 124550 4214 124602
rect 4266 124550 4278 124602
rect 4330 124550 4342 124602
rect 4394 124550 4406 124602
rect 4458 124550 4470 124602
rect 4522 124550 7912 124602
rect 1104 124528 7912 124550
rect 104052 124602 108836 124624
rect 104052 124550 105922 124602
rect 105974 124550 105986 124602
rect 106038 124550 106050 124602
rect 106102 124550 106114 124602
rect 106166 124550 106178 124602
rect 106230 124550 108836 124602
rect 104052 124528 108836 124550
rect 1104 124058 7912 124080
rect 1104 124006 4874 124058
rect 4926 124006 4938 124058
rect 4990 124006 5002 124058
rect 5054 124006 5066 124058
rect 5118 124006 5130 124058
rect 5182 124006 7912 124058
rect 1104 123984 7912 124006
rect 104052 124058 108836 124080
rect 104052 124006 106658 124058
rect 106710 124006 106722 124058
rect 106774 124006 106786 124058
rect 106838 124006 106850 124058
rect 106902 124006 106914 124058
rect 106966 124006 108836 124058
rect 104052 123984 108836 124006
rect 1104 123514 7912 123536
rect 1104 123462 4214 123514
rect 4266 123462 4278 123514
rect 4330 123462 4342 123514
rect 4394 123462 4406 123514
rect 4458 123462 4470 123514
rect 4522 123462 7912 123514
rect 1104 123440 7912 123462
rect 104052 123514 108836 123536
rect 104052 123462 105922 123514
rect 105974 123462 105986 123514
rect 106038 123462 106050 123514
rect 106102 123462 106114 123514
rect 106166 123462 106178 123514
rect 106230 123462 108836 123514
rect 104052 123440 108836 123462
rect 1104 122970 7912 122992
rect 1104 122918 4874 122970
rect 4926 122918 4938 122970
rect 4990 122918 5002 122970
rect 5054 122918 5066 122970
rect 5118 122918 5130 122970
rect 5182 122918 7912 122970
rect 1104 122896 7912 122918
rect 104052 122970 108836 122992
rect 104052 122918 106658 122970
rect 106710 122918 106722 122970
rect 106774 122918 106786 122970
rect 106838 122918 106850 122970
rect 106902 122918 106914 122970
rect 106966 122918 108836 122970
rect 104052 122896 108836 122918
rect 1104 122426 7912 122448
rect 1104 122374 4214 122426
rect 4266 122374 4278 122426
rect 4330 122374 4342 122426
rect 4394 122374 4406 122426
rect 4458 122374 4470 122426
rect 4522 122374 7912 122426
rect 1104 122352 7912 122374
rect 104052 122426 108836 122448
rect 104052 122374 105922 122426
rect 105974 122374 105986 122426
rect 106038 122374 106050 122426
rect 106102 122374 106114 122426
rect 106166 122374 106178 122426
rect 106230 122374 108836 122426
rect 104052 122352 108836 122374
rect 1104 121882 7912 121904
rect 1104 121830 4874 121882
rect 4926 121830 4938 121882
rect 4990 121830 5002 121882
rect 5054 121830 5066 121882
rect 5118 121830 5130 121882
rect 5182 121830 7912 121882
rect 1104 121808 7912 121830
rect 104052 121882 108836 121904
rect 104052 121830 106658 121882
rect 106710 121830 106722 121882
rect 106774 121830 106786 121882
rect 106838 121830 106850 121882
rect 106902 121830 106914 121882
rect 106966 121830 108836 121882
rect 104052 121808 108836 121830
rect 1104 121338 7912 121360
rect 1104 121286 4214 121338
rect 4266 121286 4278 121338
rect 4330 121286 4342 121338
rect 4394 121286 4406 121338
rect 4458 121286 4470 121338
rect 4522 121286 7912 121338
rect 1104 121264 7912 121286
rect 104052 121338 108836 121360
rect 104052 121286 105922 121338
rect 105974 121286 105986 121338
rect 106038 121286 106050 121338
rect 106102 121286 106114 121338
rect 106166 121286 106178 121338
rect 106230 121286 108836 121338
rect 104052 121264 108836 121286
rect 1104 120794 7912 120816
rect 1104 120742 4874 120794
rect 4926 120742 4938 120794
rect 4990 120742 5002 120794
rect 5054 120742 5066 120794
rect 5118 120742 5130 120794
rect 5182 120742 7912 120794
rect 1104 120720 7912 120742
rect 104052 120794 108836 120816
rect 104052 120742 106658 120794
rect 106710 120742 106722 120794
rect 106774 120742 106786 120794
rect 106838 120742 106850 120794
rect 106902 120742 106914 120794
rect 106966 120742 108836 120794
rect 104052 120720 108836 120742
rect 1104 120250 7912 120272
rect 1104 120198 4214 120250
rect 4266 120198 4278 120250
rect 4330 120198 4342 120250
rect 4394 120198 4406 120250
rect 4458 120198 4470 120250
rect 4522 120198 7912 120250
rect 1104 120176 7912 120198
rect 104052 120250 108836 120272
rect 104052 120198 105922 120250
rect 105974 120198 105986 120250
rect 106038 120198 106050 120250
rect 106102 120198 106114 120250
rect 106166 120198 106178 120250
rect 106230 120198 108836 120250
rect 104052 120176 108836 120198
rect 1104 119706 7912 119728
rect 1104 119654 4874 119706
rect 4926 119654 4938 119706
rect 4990 119654 5002 119706
rect 5054 119654 5066 119706
rect 5118 119654 5130 119706
rect 5182 119654 7912 119706
rect 1104 119632 7912 119654
rect 104052 119706 108836 119728
rect 104052 119654 106658 119706
rect 106710 119654 106722 119706
rect 106774 119654 106786 119706
rect 106838 119654 106850 119706
rect 106902 119654 106914 119706
rect 106966 119654 108836 119706
rect 104052 119632 108836 119654
rect 1104 119162 7912 119184
rect 1104 119110 4214 119162
rect 4266 119110 4278 119162
rect 4330 119110 4342 119162
rect 4394 119110 4406 119162
rect 4458 119110 4470 119162
rect 4522 119110 7912 119162
rect 1104 119088 7912 119110
rect 104052 119162 108836 119184
rect 104052 119110 105922 119162
rect 105974 119110 105986 119162
rect 106038 119110 106050 119162
rect 106102 119110 106114 119162
rect 106166 119110 106178 119162
rect 106230 119110 108836 119162
rect 104052 119088 108836 119110
rect 1104 118618 7912 118640
rect 1104 118566 4874 118618
rect 4926 118566 4938 118618
rect 4990 118566 5002 118618
rect 5054 118566 5066 118618
rect 5118 118566 5130 118618
rect 5182 118566 7912 118618
rect 1104 118544 7912 118566
rect 104052 118618 108836 118640
rect 104052 118566 106658 118618
rect 106710 118566 106722 118618
rect 106774 118566 106786 118618
rect 106838 118566 106850 118618
rect 106902 118566 106914 118618
rect 106966 118566 108836 118618
rect 104052 118544 108836 118566
rect 7374 118464 7380 118516
rect 7432 118504 7438 118516
rect 7469 118507 7527 118513
rect 7469 118504 7481 118507
rect 7432 118476 7481 118504
rect 7432 118464 7438 118476
rect 7469 118473 7481 118476
rect 7515 118473 7527 118507
rect 7469 118467 7527 118473
rect 1104 118074 7912 118096
rect 1104 118022 4214 118074
rect 4266 118022 4278 118074
rect 4330 118022 4342 118074
rect 4394 118022 4406 118074
rect 4458 118022 4470 118074
rect 4522 118022 7912 118074
rect 1104 118000 7912 118022
rect 104052 118074 108836 118096
rect 104052 118022 105922 118074
rect 105974 118022 105986 118074
rect 106038 118022 106050 118074
rect 106102 118022 106114 118074
rect 106166 118022 106178 118074
rect 106230 118022 108836 118074
rect 104052 118000 108836 118022
rect 6181 117759 6239 117765
rect 6181 117725 6193 117759
rect 6227 117756 6239 117759
rect 7466 117756 7472 117768
rect 6227 117728 7472 117756
rect 6227 117725 6239 117728
rect 6181 117719 6239 117725
rect 7466 117716 7472 117728
rect 7524 117716 7530 117768
rect 6448 117691 6506 117697
rect 6448 117657 6460 117691
rect 6494 117688 6506 117691
rect 7374 117688 7380 117700
rect 6494 117660 7380 117688
rect 6494 117657 6506 117660
rect 6448 117651 6506 117657
rect 7374 117648 7380 117660
rect 7432 117648 7438 117700
rect 7282 117580 7288 117632
rect 7340 117620 7346 117632
rect 7561 117623 7619 117629
rect 7561 117620 7573 117623
rect 7340 117592 7573 117620
rect 7340 117580 7346 117592
rect 7561 117589 7573 117592
rect 7607 117589 7619 117623
rect 7561 117583 7619 117589
rect 1104 117530 7912 117552
rect 1104 117478 4874 117530
rect 4926 117478 4938 117530
rect 4990 117478 5002 117530
rect 5054 117478 5066 117530
rect 5118 117478 5130 117530
rect 5182 117478 7912 117530
rect 1104 117456 7912 117478
rect 104052 117530 108836 117552
rect 104052 117478 106658 117530
rect 106710 117478 106722 117530
rect 106774 117478 106786 117530
rect 106838 117478 106850 117530
rect 106902 117478 106914 117530
rect 106966 117478 108836 117530
rect 104052 117456 108836 117478
rect 7282 117036 7288 117088
rect 7340 117036 7346 117088
rect 7466 117036 7472 117088
rect 7524 117036 7530 117088
rect 1104 116986 7912 117008
rect 1104 116934 4214 116986
rect 4266 116934 4278 116986
rect 4330 116934 4342 116986
rect 4394 116934 4406 116986
rect 4458 116934 4470 116986
rect 4522 116934 7912 116986
rect 1104 116912 7912 116934
rect 104052 116986 108836 117008
rect 104052 116934 105922 116986
rect 105974 116934 105986 116986
rect 106038 116934 106050 116986
rect 106102 116934 106114 116986
rect 106166 116934 106178 116986
rect 106230 116934 108836 116986
rect 104052 116912 108836 116934
rect 1104 116442 7912 116464
rect 1104 116390 4874 116442
rect 4926 116390 4938 116442
rect 4990 116390 5002 116442
rect 5054 116390 5066 116442
rect 5118 116390 5130 116442
rect 5182 116390 7912 116442
rect 1104 116368 7912 116390
rect 104052 116442 108836 116464
rect 104052 116390 106658 116442
rect 106710 116390 106722 116442
rect 106774 116390 106786 116442
rect 106838 116390 106850 116442
rect 106902 116390 106914 116442
rect 106966 116390 108836 116442
rect 104052 116368 108836 116390
rect 1104 115898 7912 115920
rect 1104 115846 4214 115898
rect 4266 115846 4278 115898
rect 4330 115846 4342 115898
rect 4394 115846 4406 115898
rect 4458 115846 4470 115898
rect 4522 115846 7912 115898
rect 1104 115824 7912 115846
rect 104052 115898 108836 115920
rect 104052 115846 105922 115898
rect 105974 115846 105986 115898
rect 106038 115846 106050 115898
rect 106102 115846 106114 115898
rect 106166 115846 106178 115898
rect 106230 115846 108836 115898
rect 104052 115824 108836 115846
rect 1104 115354 7912 115376
rect 1104 115302 4874 115354
rect 4926 115302 4938 115354
rect 4990 115302 5002 115354
rect 5054 115302 5066 115354
rect 5118 115302 5130 115354
rect 5182 115302 7912 115354
rect 1104 115280 7912 115302
rect 104052 115354 108836 115376
rect 104052 115302 106658 115354
rect 106710 115302 106722 115354
rect 106774 115302 106786 115354
rect 106838 115302 106850 115354
rect 106902 115302 106914 115354
rect 106966 115302 108836 115354
rect 104052 115280 108836 115302
rect 1104 114810 7912 114832
rect 1104 114758 4214 114810
rect 4266 114758 4278 114810
rect 4330 114758 4342 114810
rect 4394 114758 4406 114810
rect 4458 114758 4470 114810
rect 4522 114758 7912 114810
rect 1104 114736 7912 114758
rect 104052 114810 108836 114832
rect 104052 114758 105922 114810
rect 105974 114758 105986 114810
rect 106038 114758 106050 114810
rect 106102 114758 106114 114810
rect 106166 114758 106178 114810
rect 106230 114758 108836 114810
rect 104052 114736 108836 114758
rect 1104 114266 7912 114288
rect 1104 114214 4874 114266
rect 4926 114214 4938 114266
rect 4990 114214 5002 114266
rect 5054 114214 5066 114266
rect 5118 114214 5130 114266
rect 5182 114214 7912 114266
rect 1104 114192 7912 114214
rect 104052 114266 108836 114288
rect 104052 114214 106658 114266
rect 106710 114214 106722 114266
rect 106774 114214 106786 114266
rect 106838 114214 106850 114266
rect 106902 114214 106914 114266
rect 106966 114214 108836 114266
rect 104052 114192 108836 114214
rect 1104 113722 7912 113744
rect 1104 113670 4214 113722
rect 4266 113670 4278 113722
rect 4330 113670 4342 113722
rect 4394 113670 4406 113722
rect 4458 113670 4470 113722
rect 4522 113670 7912 113722
rect 1104 113648 7912 113670
rect 104052 113722 108836 113744
rect 104052 113670 105922 113722
rect 105974 113670 105986 113722
rect 106038 113670 106050 113722
rect 106102 113670 106114 113722
rect 106166 113670 106178 113722
rect 106230 113670 108836 113722
rect 104052 113648 108836 113670
rect 104342 113568 104348 113620
rect 104400 113608 104406 113620
rect 105630 113608 105636 113620
rect 104400 113580 105636 113608
rect 104400 113568 104406 113580
rect 105630 113568 105636 113580
rect 105688 113608 105694 113620
rect 106001 113611 106059 113617
rect 106001 113608 106013 113611
rect 105688 113580 106013 113608
rect 105688 113568 105694 113580
rect 106001 113577 106013 113580
rect 106047 113577 106059 113611
rect 106001 113571 106059 113577
rect 104342 113432 104348 113484
rect 104400 113432 104406 113484
rect 104612 113407 104670 113413
rect 104612 113373 104624 113407
rect 104658 113373 104670 113407
rect 104612 113367 104670 113373
rect 104526 113296 104532 113348
rect 104584 113336 104590 113348
rect 104636 113336 104664 113367
rect 104584 113308 104664 113336
rect 104584 113296 104590 113308
rect 102870 113228 102876 113280
rect 102928 113268 102934 113280
rect 105725 113271 105783 113277
rect 105725 113268 105737 113271
rect 102928 113240 105737 113268
rect 102928 113228 102934 113240
rect 105725 113237 105737 113240
rect 105771 113268 105783 113271
rect 105817 113271 105875 113277
rect 105817 113268 105829 113271
rect 105771 113240 105829 113268
rect 105771 113237 105783 113240
rect 105725 113231 105783 113237
rect 105817 113237 105829 113240
rect 105863 113237 105875 113271
rect 105817 113231 105875 113237
rect 1104 113178 7912 113200
rect 1104 113126 4874 113178
rect 4926 113126 4938 113178
rect 4990 113126 5002 113178
rect 5054 113126 5066 113178
rect 5118 113126 5130 113178
rect 5182 113126 7912 113178
rect 1104 113104 7912 113126
rect 104052 113178 108836 113200
rect 104052 113126 106658 113178
rect 106710 113126 106722 113178
rect 106774 113126 106786 113178
rect 106838 113126 106850 113178
rect 106902 113126 106914 113178
rect 106966 113126 108836 113178
rect 104052 113104 108836 113126
rect 104437 113067 104495 113073
rect 104437 113033 104449 113067
rect 104483 113064 104495 113067
rect 104526 113064 104532 113076
rect 104483 113036 104532 113064
rect 104483 113033 104495 113036
rect 104437 113027 104495 113033
rect 104526 113024 104532 113036
rect 104584 113024 104590 113076
rect 1104 112634 7912 112656
rect 1104 112582 4214 112634
rect 4266 112582 4278 112634
rect 4330 112582 4342 112634
rect 4394 112582 4406 112634
rect 4458 112582 4470 112634
rect 4522 112582 7912 112634
rect 1104 112560 7912 112582
rect 104052 112634 108836 112656
rect 104052 112582 105922 112634
rect 105974 112582 105986 112634
rect 106038 112582 106050 112634
rect 106102 112582 106114 112634
rect 106166 112582 106178 112634
rect 106230 112582 108836 112634
rect 104052 112560 108836 112582
rect 1104 112090 7912 112112
rect 1104 112038 4874 112090
rect 4926 112038 4938 112090
rect 4990 112038 5002 112090
rect 5054 112038 5066 112090
rect 5118 112038 5130 112090
rect 5182 112038 7912 112090
rect 1104 112016 7912 112038
rect 104052 112090 108836 112112
rect 104052 112038 106658 112090
rect 106710 112038 106722 112090
rect 106774 112038 106786 112090
rect 106838 112038 106850 112090
rect 106902 112038 106914 112090
rect 106966 112038 108836 112090
rect 104052 112016 108836 112038
rect 1104 111546 7912 111568
rect 1104 111494 4214 111546
rect 4266 111494 4278 111546
rect 4330 111494 4342 111546
rect 4394 111494 4406 111546
rect 4458 111494 4470 111546
rect 4522 111494 7912 111546
rect 1104 111472 7912 111494
rect 104052 111546 108836 111568
rect 104052 111494 105922 111546
rect 105974 111494 105986 111546
rect 106038 111494 106050 111546
rect 106102 111494 106114 111546
rect 106166 111494 106178 111546
rect 106230 111494 108836 111546
rect 104052 111472 108836 111494
rect 1581 111367 1639 111373
rect 1581 111333 1593 111367
rect 1627 111364 1639 111367
rect 9490 111364 9496 111376
rect 1627 111336 9496 111364
rect 1627 111333 1639 111336
rect 1581 111327 1639 111333
rect 9490 111324 9496 111336
rect 9548 111324 9554 111376
rect 1302 111188 1308 111240
rect 1360 111228 1366 111240
rect 1397 111231 1455 111237
rect 1397 111228 1409 111231
rect 1360 111200 1409 111228
rect 1360 111188 1366 111200
rect 1397 111197 1409 111200
rect 1443 111228 1455 111231
rect 1673 111231 1731 111237
rect 1673 111228 1685 111231
rect 1443 111200 1685 111228
rect 1443 111197 1455 111200
rect 1397 111191 1455 111197
rect 1673 111197 1685 111200
rect 1719 111197 1731 111231
rect 1673 111191 1731 111197
rect 1104 111002 7912 111024
rect 1104 110950 4874 111002
rect 4926 110950 4938 111002
rect 4990 110950 5002 111002
rect 5054 110950 5066 111002
rect 5118 110950 5130 111002
rect 5182 110950 7912 111002
rect 1104 110928 7912 110950
rect 104052 111002 108836 111024
rect 104052 110950 106658 111002
rect 106710 110950 106722 111002
rect 106774 110950 106786 111002
rect 106838 110950 106850 111002
rect 106902 110950 106914 111002
rect 106966 110950 108836 111002
rect 104052 110928 108836 110950
rect 1104 110458 7912 110480
rect 1104 110406 4214 110458
rect 4266 110406 4278 110458
rect 4330 110406 4342 110458
rect 4394 110406 4406 110458
rect 4458 110406 4470 110458
rect 4522 110406 7912 110458
rect 1104 110384 7912 110406
rect 104052 110458 108836 110480
rect 104052 110406 105922 110458
rect 105974 110406 105986 110458
rect 106038 110406 106050 110458
rect 106102 110406 106114 110458
rect 106166 110406 106178 110458
rect 106230 110406 108836 110458
rect 104052 110384 108836 110406
rect 1104 109914 7912 109936
rect 1104 109862 4874 109914
rect 4926 109862 4938 109914
rect 4990 109862 5002 109914
rect 5054 109862 5066 109914
rect 5118 109862 5130 109914
rect 5182 109862 7912 109914
rect 1104 109840 7912 109862
rect 104052 109914 108836 109936
rect 104052 109862 106658 109914
rect 106710 109862 106722 109914
rect 106774 109862 106786 109914
rect 106838 109862 106850 109914
rect 106902 109862 106914 109914
rect 106966 109862 108836 109914
rect 104052 109840 108836 109862
rect 1302 109624 1308 109676
rect 1360 109664 1366 109676
rect 1397 109667 1455 109673
rect 1397 109664 1409 109667
rect 1360 109636 1409 109664
rect 1360 109624 1366 109636
rect 1397 109633 1409 109636
rect 1443 109664 1455 109667
rect 1673 109667 1731 109673
rect 1673 109664 1685 109667
rect 1443 109636 1685 109664
rect 1443 109633 1455 109636
rect 1397 109627 1455 109633
rect 1673 109633 1685 109636
rect 1719 109633 1731 109667
rect 1673 109627 1731 109633
rect 1581 109531 1639 109537
rect 1581 109497 1593 109531
rect 1627 109528 1639 109531
rect 9490 109528 9496 109540
rect 1627 109500 9496 109528
rect 1627 109497 1639 109500
rect 1581 109491 1639 109497
rect 9490 109488 9496 109500
rect 9548 109488 9554 109540
rect 1104 109370 7912 109392
rect 1104 109318 4214 109370
rect 4266 109318 4278 109370
rect 4330 109318 4342 109370
rect 4394 109318 4406 109370
rect 4458 109318 4470 109370
rect 4522 109318 7912 109370
rect 1104 109296 7912 109318
rect 104052 109370 108836 109392
rect 104052 109318 105922 109370
rect 105974 109318 105986 109370
rect 106038 109318 106050 109370
rect 106102 109318 106114 109370
rect 106166 109318 106178 109370
rect 106230 109318 108836 109370
rect 104052 109296 108836 109318
rect 1104 108826 7912 108848
rect 1104 108774 4874 108826
rect 4926 108774 4938 108826
rect 4990 108774 5002 108826
rect 5054 108774 5066 108826
rect 5118 108774 5130 108826
rect 5182 108774 7912 108826
rect 1104 108752 7912 108774
rect 104052 108826 108836 108848
rect 104052 108774 106658 108826
rect 106710 108774 106722 108826
rect 106774 108774 106786 108826
rect 106838 108774 106850 108826
rect 106902 108774 106914 108826
rect 106966 108774 108836 108826
rect 104052 108752 108836 108774
rect 1302 108536 1308 108588
rect 1360 108576 1366 108588
rect 1397 108579 1455 108585
rect 1397 108576 1409 108579
rect 1360 108548 1409 108576
rect 1360 108536 1366 108548
rect 1397 108545 1409 108548
rect 1443 108576 1455 108579
rect 1673 108579 1731 108585
rect 1673 108576 1685 108579
rect 1443 108548 1685 108576
rect 1443 108545 1455 108548
rect 1397 108539 1455 108545
rect 1673 108545 1685 108548
rect 1719 108545 1731 108579
rect 1673 108539 1731 108545
rect 1581 108443 1639 108449
rect 1581 108409 1593 108443
rect 1627 108440 1639 108443
rect 9490 108440 9496 108452
rect 1627 108412 9496 108440
rect 1627 108409 1639 108412
rect 1581 108403 1639 108409
rect 9490 108400 9496 108412
rect 9548 108400 9554 108452
rect 1104 108282 7912 108304
rect 1104 108230 4214 108282
rect 4266 108230 4278 108282
rect 4330 108230 4342 108282
rect 4394 108230 4406 108282
rect 4458 108230 4470 108282
rect 4522 108230 7912 108282
rect 1104 108208 7912 108230
rect 104052 108282 108836 108304
rect 104052 108230 105922 108282
rect 105974 108230 105986 108282
rect 106038 108230 106050 108282
rect 106102 108230 106114 108282
rect 106166 108230 106178 108282
rect 106230 108230 108836 108282
rect 104052 108208 108836 108230
rect 1104 107738 7912 107760
rect 1104 107686 4874 107738
rect 4926 107686 4938 107738
rect 4990 107686 5002 107738
rect 5054 107686 5066 107738
rect 5118 107686 5130 107738
rect 5182 107686 7912 107738
rect 1104 107664 7912 107686
rect 104052 107738 108836 107760
rect 104052 107686 106658 107738
rect 106710 107686 106722 107738
rect 106774 107686 106786 107738
rect 106838 107686 106850 107738
rect 106902 107686 106914 107738
rect 106966 107686 108836 107738
rect 104052 107664 108836 107686
rect 1104 107194 7912 107216
rect 1104 107142 4214 107194
rect 4266 107142 4278 107194
rect 4330 107142 4342 107194
rect 4394 107142 4406 107194
rect 4458 107142 4470 107194
rect 4522 107142 7912 107194
rect 1104 107120 7912 107142
rect 104052 107194 108836 107216
rect 104052 107142 105922 107194
rect 105974 107142 105986 107194
rect 106038 107142 106050 107194
rect 106102 107142 106114 107194
rect 106166 107142 106178 107194
rect 106230 107142 108836 107194
rect 104052 107120 108836 107142
rect 105630 107040 105636 107092
rect 105688 107080 105694 107092
rect 105814 107080 105820 107092
rect 105688 107052 105820 107080
rect 105688 107040 105694 107052
rect 105814 107040 105820 107052
rect 105872 107080 105878 107092
rect 106369 107083 106427 107089
rect 106369 107080 106381 107083
rect 105872 107052 106381 107080
rect 105872 107040 105878 107052
rect 106369 107049 106381 107052
rect 106415 107049 106427 107083
rect 106369 107043 106427 107049
rect 1581 107015 1639 107021
rect 1581 106981 1593 107015
rect 1627 107012 1639 107015
rect 9490 107012 9496 107024
rect 1627 106984 9496 107012
rect 1627 106981 1639 106984
rect 1581 106975 1639 106981
rect 9490 106972 9496 106984
rect 9548 106972 9554 107024
rect 1210 106836 1216 106888
rect 1268 106876 1274 106888
rect 1397 106879 1455 106885
rect 1397 106876 1409 106879
rect 1268 106848 1409 106876
rect 1268 106836 1274 106848
rect 1397 106845 1409 106848
rect 1443 106876 1455 106879
rect 1673 106879 1731 106885
rect 1673 106876 1685 106879
rect 1443 106848 1685 106876
rect 1443 106845 1455 106848
rect 1397 106839 1455 106845
rect 1673 106845 1685 106848
rect 1719 106845 1731 106879
rect 1673 106839 1731 106845
rect 104345 106811 104403 106817
rect 104345 106777 104357 106811
rect 104391 106808 104403 106811
rect 105078 106808 105084 106820
rect 104391 106780 105084 106808
rect 104391 106777 104403 106780
rect 104345 106771 104403 106777
rect 105078 106768 105084 106780
rect 105136 106808 105142 106820
rect 106277 106811 106335 106817
rect 106277 106808 106289 106811
rect 105136 106780 106289 106808
rect 105136 106768 105142 106780
rect 106277 106777 106289 106780
rect 106323 106777 106335 106811
rect 106277 106771 106335 106777
rect 1104 106650 7912 106672
rect 1104 106598 4874 106650
rect 4926 106598 4938 106650
rect 4990 106598 5002 106650
rect 5054 106598 5066 106650
rect 5118 106598 5130 106650
rect 5182 106598 7912 106650
rect 1104 106576 7912 106598
rect 104052 106650 108836 106672
rect 104052 106598 106658 106650
rect 106710 106598 106722 106650
rect 106774 106598 106786 106650
rect 106838 106598 106850 106650
rect 106902 106598 106914 106650
rect 106966 106598 108836 106650
rect 104052 106576 108836 106598
rect 1104 106106 7912 106128
rect 1104 106054 4214 106106
rect 4266 106054 4278 106106
rect 4330 106054 4342 106106
rect 4394 106054 4406 106106
rect 4458 106054 4470 106106
rect 4522 106054 7912 106106
rect 1104 106032 7912 106054
rect 104052 106106 108836 106128
rect 104052 106054 105922 106106
rect 105974 106054 105986 106106
rect 106038 106054 106050 106106
rect 106102 106054 106114 106106
rect 106166 106054 106178 106106
rect 106230 106054 108836 106106
rect 104052 106032 108836 106054
rect 1581 105927 1639 105933
rect 1581 105893 1593 105927
rect 1627 105924 1639 105927
rect 9490 105924 9496 105936
rect 1627 105896 9496 105924
rect 1627 105893 1639 105896
rect 1581 105887 1639 105893
rect 9490 105884 9496 105896
rect 9548 105884 9554 105936
rect 1302 105748 1308 105800
rect 1360 105788 1366 105800
rect 1397 105791 1455 105797
rect 1397 105788 1409 105791
rect 1360 105760 1409 105788
rect 1360 105748 1366 105760
rect 1397 105757 1409 105760
rect 1443 105788 1455 105791
rect 1673 105791 1731 105797
rect 1673 105788 1685 105791
rect 1443 105760 1685 105788
rect 1443 105757 1455 105760
rect 1397 105751 1455 105757
rect 1673 105757 1685 105760
rect 1719 105757 1731 105791
rect 1673 105751 1731 105757
rect 1104 105562 7912 105584
rect 1104 105510 4874 105562
rect 4926 105510 4938 105562
rect 4990 105510 5002 105562
rect 5054 105510 5066 105562
rect 5118 105510 5130 105562
rect 5182 105510 7912 105562
rect 1104 105488 7912 105510
rect 104052 105562 108836 105584
rect 104052 105510 106658 105562
rect 106710 105510 106722 105562
rect 106774 105510 106786 105562
rect 106838 105510 106850 105562
rect 106902 105510 106914 105562
rect 106966 105510 108836 105562
rect 104052 105488 108836 105510
rect 1104 105018 7912 105040
rect 1104 104966 4214 105018
rect 4266 104966 4278 105018
rect 4330 104966 4342 105018
rect 4394 104966 4406 105018
rect 4458 104966 4470 105018
rect 4522 104966 7912 105018
rect 1104 104944 7912 104966
rect 104052 105018 108836 105040
rect 104052 104966 105922 105018
rect 105974 104966 105986 105018
rect 106038 104966 106050 105018
rect 106102 104966 106114 105018
rect 106166 104966 106178 105018
rect 106230 104966 108836 105018
rect 104052 104944 108836 104966
rect 1104 104474 7912 104496
rect 1104 104422 4874 104474
rect 4926 104422 4938 104474
rect 4990 104422 5002 104474
rect 5054 104422 5066 104474
rect 5118 104422 5130 104474
rect 5182 104422 7912 104474
rect 1104 104400 7912 104422
rect 104052 104474 108836 104496
rect 104052 104422 106658 104474
rect 106710 104422 106722 104474
rect 106774 104422 106786 104474
rect 106838 104422 106850 104474
rect 106902 104422 106914 104474
rect 106966 104422 108836 104474
rect 104052 104400 108836 104422
rect 1302 104184 1308 104236
rect 1360 104224 1366 104236
rect 1397 104227 1455 104233
rect 1397 104224 1409 104227
rect 1360 104196 1409 104224
rect 1360 104184 1366 104196
rect 1397 104193 1409 104196
rect 1443 104224 1455 104227
rect 1673 104227 1731 104233
rect 1673 104224 1685 104227
rect 1443 104196 1685 104224
rect 1443 104193 1455 104196
rect 1397 104187 1455 104193
rect 1673 104193 1685 104196
rect 1719 104193 1731 104227
rect 1673 104187 1731 104193
rect 1581 104091 1639 104097
rect 1581 104057 1593 104091
rect 1627 104088 1639 104091
rect 9490 104088 9496 104100
rect 1627 104060 9496 104088
rect 1627 104057 1639 104060
rect 1581 104051 1639 104057
rect 9490 104048 9496 104060
rect 9548 104048 9554 104100
rect 1104 103930 7912 103952
rect 1104 103878 4214 103930
rect 4266 103878 4278 103930
rect 4330 103878 4342 103930
rect 4394 103878 4406 103930
rect 4458 103878 4470 103930
rect 4522 103878 7912 103930
rect 1104 103856 7912 103878
rect 104052 103930 108836 103952
rect 104052 103878 105922 103930
rect 105974 103878 105986 103930
rect 106038 103878 106050 103930
rect 106102 103878 106114 103930
rect 106166 103878 106178 103930
rect 106230 103878 108836 103930
rect 104052 103856 108836 103878
rect 1104 103386 7912 103408
rect 1104 103334 4874 103386
rect 4926 103334 4938 103386
rect 4990 103334 5002 103386
rect 5054 103334 5066 103386
rect 5118 103334 5130 103386
rect 5182 103334 7912 103386
rect 1104 103312 7912 103334
rect 104052 103386 108836 103408
rect 104052 103334 106658 103386
rect 106710 103334 106722 103386
rect 106774 103334 106786 103386
rect 106838 103334 106850 103386
rect 106902 103334 106914 103386
rect 106966 103334 108836 103386
rect 104052 103312 108836 103334
rect 1104 102842 7912 102864
rect 1104 102790 4214 102842
rect 4266 102790 4278 102842
rect 4330 102790 4342 102842
rect 4394 102790 4406 102842
rect 4458 102790 4470 102842
rect 4522 102790 7912 102842
rect 1104 102768 7912 102790
rect 104052 102842 108836 102864
rect 104052 102790 105922 102842
rect 105974 102790 105986 102842
rect 106038 102790 106050 102842
rect 106102 102790 106114 102842
rect 106166 102790 106178 102842
rect 106230 102790 108836 102842
rect 104052 102768 108836 102790
rect 1104 102298 7912 102320
rect 1104 102246 4874 102298
rect 4926 102246 4938 102298
rect 4990 102246 5002 102298
rect 5054 102246 5066 102298
rect 5118 102246 5130 102298
rect 5182 102246 7912 102298
rect 1104 102224 7912 102246
rect 104052 102298 108836 102320
rect 104052 102246 106658 102298
rect 106710 102246 106722 102298
rect 106774 102246 106786 102298
rect 106838 102246 106850 102298
rect 106902 102246 106914 102298
rect 106966 102246 108836 102298
rect 104052 102224 108836 102246
rect 7282 102144 7288 102196
rect 7340 102184 7346 102196
rect 9122 102184 9128 102196
rect 7340 102156 9128 102184
rect 7340 102144 7346 102156
rect 9122 102144 9128 102156
rect 9180 102144 9186 102196
rect 1104 101754 7912 101776
rect 1104 101702 4214 101754
rect 4266 101702 4278 101754
rect 4330 101702 4342 101754
rect 4394 101702 4406 101754
rect 4458 101702 4470 101754
rect 4522 101702 7912 101754
rect 1104 101680 7912 101702
rect 104052 101754 108836 101776
rect 104052 101702 105922 101754
rect 105974 101702 105986 101754
rect 106038 101702 106050 101754
rect 106102 101702 106114 101754
rect 106166 101702 106178 101754
rect 106230 101702 108836 101754
rect 104052 101680 108836 101702
rect 1104 101210 7912 101232
rect 1104 101158 4874 101210
rect 4926 101158 4938 101210
rect 4990 101158 5002 101210
rect 5054 101158 5066 101210
rect 5118 101158 5130 101210
rect 5182 101158 7912 101210
rect 1104 101136 7912 101158
rect 104052 101210 108836 101232
rect 104052 101158 106658 101210
rect 106710 101158 106722 101210
rect 106774 101158 106786 101210
rect 106838 101158 106850 101210
rect 106902 101158 106914 101210
rect 106966 101158 108836 101210
rect 104052 101136 108836 101158
rect 7374 101056 7380 101108
rect 7432 101096 7438 101108
rect 7561 101099 7619 101105
rect 7561 101096 7573 101099
rect 7432 101068 7573 101096
rect 7432 101056 7438 101068
rect 7561 101065 7573 101068
rect 7607 101096 7619 101099
rect 9030 101096 9036 101108
rect 7607 101068 9036 101096
rect 7607 101065 7619 101068
rect 7561 101059 7619 101065
rect 9030 101056 9036 101068
rect 9088 101056 9094 101108
rect 104618 101037 104624 101040
rect 104612 101028 104624 101037
rect 104579 101000 104624 101028
rect 104612 100991 104624 101000
rect 104618 100988 104624 100991
rect 104676 100988 104682 101040
rect 104345 100895 104403 100901
rect 104345 100861 104357 100895
rect 104391 100861 104403 100895
rect 104345 100855 104403 100861
rect 104360 100756 104388 100855
rect 105814 100852 105820 100904
rect 105872 100852 105878 100904
rect 105630 100784 105636 100836
rect 105688 100824 105694 100836
rect 105832 100824 105860 100852
rect 106001 100827 106059 100833
rect 106001 100824 106013 100827
rect 105688 100796 106013 100824
rect 105688 100784 105694 100796
rect 106001 100793 106013 100796
rect 106047 100793 106059 100827
rect 106001 100787 106059 100793
rect 105648 100756 105676 100784
rect 104360 100728 105676 100756
rect 105725 100759 105783 100765
rect 105725 100725 105737 100759
rect 105771 100756 105783 100759
rect 105814 100756 105820 100768
rect 105771 100728 105820 100756
rect 105771 100725 105783 100728
rect 105725 100719 105783 100725
rect 105814 100716 105820 100728
rect 105872 100716 105878 100768
rect 1104 100666 7912 100688
rect 1104 100614 4214 100666
rect 4266 100614 4278 100666
rect 4330 100614 4342 100666
rect 4394 100614 4406 100666
rect 4458 100614 4470 100666
rect 4522 100614 7912 100666
rect 1104 100592 7912 100614
rect 104052 100666 108836 100688
rect 104052 100614 105922 100666
rect 105974 100614 105986 100666
rect 106038 100614 106050 100666
rect 106102 100614 106114 100666
rect 106166 100614 106178 100666
rect 106230 100614 108836 100666
rect 104052 100592 108836 100614
rect 104437 100555 104495 100561
rect 104437 100521 104449 100555
rect 104483 100552 104495 100555
rect 104618 100552 104624 100564
rect 104483 100524 104624 100552
rect 104483 100521 104495 100524
rect 104437 100515 104495 100521
rect 104618 100512 104624 100524
rect 104676 100512 104682 100564
rect 6181 100351 6239 100357
rect 6181 100317 6193 100351
rect 6227 100348 6239 100351
rect 7466 100348 7472 100360
rect 6227 100320 7472 100348
rect 6227 100317 6239 100320
rect 6181 100311 6239 100317
rect 7466 100308 7472 100320
rect 7524 100308 7530 100360
rect 6448 100283 6506 100289
rect 6448 100249 6460 100283
rect 6494 100280 6506 100283
rect 7374 100280 7380 100292
rect 6494 100252 7380 100280
rect 6494 100249 6506 100252
rect 6448 100243 6506 100249
rect 7374 100240 7380 100252
rect 7432 100240 7438 100292
rect 7282 100172 7288 100224
rect 7340 100212 7346 100224
rect 7561 100215 7619 100221
rect 7561 100212 7573 100215
rect 7340 100184 7573 100212
rect 7340 100172 7346 100184
rect 7561 100181 7573 100184
rect 7607 100181 7619 100215
rect 7561 100175 7619 100181
rect 1104 100122 7912 100144
rect 1104 100070 4874 100122
rect 4926 100070 4938 100122
rect 4990 100070 5002 100122
rect 5054 100070 5066 100122
rect 5118 100070 5130 100122
rect 5182 100070 7912 100122
rect 1104 100048 7912 100070
rect 104052 100122 108836 100144
rect 104052 100070 106658 100122
rect 106710 100070 106722 100122
rect 106774 100070 106786 100122
rect 106838 100070 106850 100122
rect 106902 100070 106914 100122
rect 106966 100070 108836 100122
rect 104052 100048 108836 100070
rect 7466 99968 7472 100020
rect 7524 99968 7530 100020
rect 7282 99628 7288 99680
rect 7340 99628 7346 99680
rect 1104 99578 7912 99600
rect 1104 99526 4214 99578
rect 4266 99526 4278 99578
rect 4330 99526 4342 99578
rect 4394 99526 4406 99578
rect 4458 99526 4470 99578
rect 4522 99526 7912 99578
rect 1104 99504 7912 99526
rect 104052 99578 108836 99600
rect 104052 99526 105922 99578
rect 105974 99526 105986 99578
rect 106038 99526 106050 99578
rect 106102 99526 106114 99578
rect 106166 99526 106178 99578
rect 106230 99526 108836 99578
rect 104052 99504 108836 99526
rect 1104 99034 7912 99056
rect 1104 98982 4874 99034
rect 4926 98982 4938 99034
rect 4990 98982 5002 99034
rect 5054 98982 5066 99034
rect 5118 98982 5130 99034
rect 5182 98982 7912 99034
rect 1104 98960 7912 98982
rect 104052 99034 108836 99056
rect 104052 98982 106658 99034
rect 106710 98982 106722 99034
rect 106774 98982 106786 99034
rect 106838 98982 106850 99034
rect 106902 98982 106914 99034
rect 106966 98982 108836 99034
rect 104052 98960 108836 98982
rect 1104 98490 7912 98512
rect 1104 98438 4214 98490
rect 4266 98438 4278 98490
rect 4330 98438 4342 98490
rect 4394 98438 4406 98490
rect 4458 98438 4470 98490
rect 4522 98438 7912 98490
rect 1104 98416 7912 98438
rect 104052 98490 108836 98512
rect 104052 98438 105922 98490
rect 105974 98438 105986 98490
rect 106038 98438 106050 98490
rect 106102 98438 106114 98490
rect 106166 98438 106178 98490
rect 106230 98438 108836 98490
rect 104052 98416 108836 98438
rect 1104 97946 7912 97968
rect 1104 97894 4874 97946
rect 4926 97894 4938 97946
rect 4990 97894 5002 97946
rect 5054 97894 5066 97946
rect 5118 97894 5130 97946
rect 5182 97894 7912 97946
rect 1104 97872 7912 97894
rect 104052 97946 108836 97968
rect 104052 97894 106658 97946
rect 106710 97894 106722 97946
rect 106774 97894 106786 97946
rect 106838 97894 106850 97946
rect 106902 97894 106914 97946
rect 106966 97894 108836 97946
rect 104052 97872 108836 97894
rect 1104 97402 7912 97424
rect 1104 97350 4214 97402
rect 4266 97350 4278 97402
rect 4330 97350 4342 97402
rect 4394 97350 4406 97402
rect 4458 97350 4470 97402
rect 4522 97350 7912 97402
rect 1104 97328 7912 97350
rect 104052 97402 108836 97424
rect 104052 97350 105922 97402
rect 105974 97350 105986 97402
rect 106038 97350 106050 97402
rect 106102 97350 106114 97402
rect 106166 97350 106178 97402
rect 106230 97350 108836 97402
rect 104052 97328 108836 97350
rect 1104 96858 7912 96880
rect 1104 96806 4874 96858
rect 4926 96806 4938 96858
rect 4990 96806 5002 96858
rect 5054 96806 5066 96858
rect 5118 96806 5130 96858
rect 5182 96806 7912 96858
rect 1104 96784 7912 96806
rect 104052 96858 108836 96880
rect 104052 96806 106658 96858
rect 106710 96806 106722 96858
rect 106774 96806 106786 96858
rect 106838 96806 106850 96858
rect 106902 96806 106914 96858
rect 106966 96806 108836 96858
rect 104052 96784 108836 96806
rect 102778 96568 102784 96620
rect 102836 96608 102842 96620
rect 104601 96611 104659 96617
rect 104601 96608 104613 96611
rect 102836 96580 104613 96608
rect 102836 96568 102842 96580
rect 1104 96314 7912 96336
rect 1104 96262 4214 96314
rect 4266 96262 4278 96314
rect 4330 96262 4342 96314
rect 4394 96262 4406 96314
rect 4458 96262 4470 96314
rect 4522 96262 7912 96314
rect 1104 96240 7912 96262
rect 103992 96200 104020 96580
rect 104601 96577 104613 96580
rect 104647 96577 104659 96611
rect 104601 96571 104659 96577
rect 104342 96500 104348 96552
rect 104400 96500 104406 96552
rect 105630 96472 105636 96484
rect 105556 96444 105636 96472
rect 104342 96364 104348 96416
rect 104400 96404 104406 96416
rect 105556 96404 105584 96444
rect 105630 96432 105636 96444
rect 105688 96472 105694 96484
rect 106001 96475 106059 96481
rect 106001 96472 106013 96475
rect 105688 96444 106013 96472
rect 105688 96432 105694 96444
rect 106001 96441 106013 96444
rect 106047 96441 106059 96475
rect 106001 96435 106059 96441
rect 104400 96376 105584 96404
rect 104400 96364 104406 96376
rect 105722 96364 105728 96416
rect 105780 96404 105786 96416
rect 105817 96407 105875 96413
rect 105817 96404 105829 96407
rect 105780 96376 105829 96404
rect 105780 96364 105786 96376
rect 105817 96373 105829 96376
rect 105863 96373 105875 96407
rect 105817 96367 105875 96373
rect 104052 96314 108836 96336
rect 104052 96262 105922 96314
rect 105974 96262 105986 96314
rect 106038 96262 106050 96314
rect 106102 96262 106114 96314
rect 106166 96262 106178 96314
rect 106230 96262 108836 96314
rect 104052 96240 108836 96262
rect 104345 96203 104403 96209
rect 104345 96200 104357 96203
rect 103992 96172 104357 96200
rect 104345 96169 104357 96172
rect 104391 96169 104403 96203
rect 104345 96163 104403 96169
rect 102962 96092 102968 96144
rect 103020 96132 103026 96144
rect 105722 96132 105728 96144
rect 103020 96104 105728 96132
rect 103020 96092 103026 96104
rect 105722 96092 105728 96104
rect 105780 96092 105786 96144
rect 1104 95770 7912 95792
rect 1104 95718 4874 95770
rect 4926 95718 4938 95770
rect 4990 95718 5002 95770
rect 5054 95718 5066 95770
rect 5118 95718 5130 95770
rect 5182 95718 7912 95770
rect 1104 95696 7912 95718
rect 104052 95770 108836 95792
rect 104052 95718 106658 95770
rect 106710 95718 106722 95770
rect 106774 95718 106786 95770
rect 106838 95718 106850 95770
rect 106902 95718 106914 95770
rect 106966 95718 108836 95770
rect 104052 95696 108836 95718
rect 7466 95616 7472 95668
rect 7524 95616 7530 95668
rect 104345 95319 104403 95325
rect 104345 95316 104357 95319
rect 103486 95288 104357 95316
rect 1104 95226 7912 95248
rect 1104 95174 4214 95226
rect 4266 95174 4278 95226
rect 4330 95174 4342 95226
rect 4394 95174 4406 95226
rect 4458 95174 4470 95226
rect 4522 95174 7912 95226
rect 1104 95152 7912 95174
rect 102502 95140 102508 95192
rect 102560 95180 102566 95192
rect 103486 95180 103514 95288
rect 104345 95285 104357 95288
rect 104391 95285 104403 95319
rect 104345 95279 104403 95285
rect 102560 95152 103514 95180
rect 104052 95226 108836 95248
rect 104052 95174 105922 95226
rect 105974 95174 105986 95226
rect 106038 95174 106050 95226
rect 106102 95174 106114 95226
rect 106166 95174 106178 95226
rect 106230 95174 108836 95226
rect 104052 95152 108836 95174
rect 102560 95140 102566 95152
rect 7466 94936 7472 94988
rect 7524 94936 7530 94988
rect 5721 94843 5779 94849
rect 5721 94809 5733 94843
rect 5767 94840 5779 94843
rect 5810 94840 5816 94852
rect 5767 94812 5816 94840
rect 5767 94809 5779 94812
rect 5721 94803 5779 94809
rect 5810 94800 5816 94812
rect 5868 94800 5874 94852
rect 1104 94682 7912 94704
rect 1104 94630 4874 94682
rect 4926 94630 4938 94682
rect 4990 94630 5002 94682
rect 5054 94630 5066 94682
rect 5118 94630 5130 94682
rect 5182 94630 7912 94682
rect 1104 94608 7912 94630
rect 104052 94682 108836 94704
rect 104052 94630 106658 94682
rect 106710 94630 106722 94682
rect 106774 94630 106786 94682
rect 106838 94630 106850 94682
rect 106902 94630 106914 94682
rect 106966 94630 108836 94682
rect 104052 94608 108836 94630
rect 6549 94435 6607 94441
rect 6549 94401 6561 94435
rect 6595 94432 6607 94435
rect 6641 94435 6699 94441
rect 6641 94432 6653 94435
rect 6595 94404 6653 94432
rect 6595 94401 6607 94404
rect 6549 94395 6607 94401
rect 6641 94401 6653 94404
rect 6687 94432 6699 94435
rect 7466 94432 7472 94444
rect 6687 94404 7472 94432
rect 6687 94401 6699 94404
rect 6641 94395 6699 94401
rect 7466 94392 7472 94404
rect 7524 94392 7530 94444
rect 1104 94138 7912 94160
rect 1104 94086 4214 94138
rect 4266 94086 4278 94138
rect 4330 94086 4342 94138
rect 4394 94086 4406 94138
rect 4458 94086 4470 94138
rect 4522 94086 7912 94138
rect 1104 94064 7912 94086
rect 104052 94138 108836 94160
rect 104052 94086 105922 94138
rect 105974 94086 105986 94138
rect 106038 94086 106050 94138
rect 106102 94086 106114 94138
rect 106166 94086 106178 94138
rect 106230 94086 108836 94138
rect 104052 94064 108836 94086
rect 6181 93823 6239 93829
rect 6181 93789 6193 93823
rect 6227 93820 6239 93823
rect 7466 93820 7472 93832
rect 6227 93792 7472 93820
rect 6227 93789 6239 93792
rect 6181 93783 6239 93789
rect 7466 93780 7472 93792
rect 7524 93780 7530 93832
rect 6448 93755 6506 93761
rect 6448 93721 6460 93755
rect 6494 93752 6506 93755
rect 8938 93752 8944 93764
rect 6494 93724 8944 93752
rect 6494 93721 6506 93724
rect 6448 93715 6506 93721
rect 7098 93644 7104 93696
rect 7156 93684 7162 93696
rect 7561 93687 7619 93693
rect 7561 93684 7573 93687
rect 7156 93656 7573 93684
rect 7156 93644 7162 93656
rect 7561 93653 7573 93656
rect 7607 93653 7619 93687
rect 7561 93647 7619 93653
rect 1104 93594 7912 93616
rect 1104 93542 4874 93594
rect 4926 93542 4938 93594
rect 4990 93542 5002 93594
rect 5054 93542 5066 93594
rect 5118 93542 5130 93594
rect 5182 93542 7912 93594
rect 1104 93520 7912 93542
rect 7377 93483 7435 93489
rect 7377 93449 7389 93483
rect 7423 93480 7435 93483
rect 7944 93480 7972 93724
rect 8938 93712 8944 93724
rect 8996 93712 9002 93764
rect 102410 93644 102416 93696
rect 102468 93684 102474 93696
rect 104345 93687 104403 93693
rect 104345 93684 104357 93687
rect 102468 93656 104357 93684
rect 102468 93644 102474 93656
rect 104345 93653 104357 93656
rect 104391 93653 104403 93687
rect 104345 93647 104403 93653
rect 104052 93594 108836 93616
rect 104052 93542 106658 93594
rect 106710 93542 106722 93594
rect 106774 93542 106786 93594
rect 106838 93542 106850 93594
rect 106902 93542 106914 93594
rect 106966 93542 108836 93594
rect 104052 93520 108836 93542
rect 7423 93452 7972 93480
rect 7423 93449 7435 93452
rect 7377 93443 7435 93449
rect 7098 93100 7104 93152
rect 7156 93100 7162 93152
rect 7466 93100 7472 93152
rect 7524 93100 7530 93152
rect 1104 93050 7912 93072
rect 1104 92998 4214 93050
rect 4266 92998 4278 93050
rect 4330 92998 4342 93050
rect 4394 92998 4406 93050
rect 4458 92998 4470 93050
rect 4522 92998 7912 93050
rect 1104 92976 7912 92998
rect 104052 93050 108836 93072
rect 104052 92998 105922 93050
rect 105974 92998 105986 93050
rect 106038 92998 106050 93050
rect 106102 92998 106114 93050
rect 106166 92998 106178 93050
rect 106230 92998 108836 93050
rect 104052 92976 108836 92998
rect 103882 92556 103888 92608
rect 103940 92596 103946 92608
rect 104345 92599 104403 92605
rect 104345 92596 104357 92599
rect 103940 92568 104357 92596
rect 103940 92556 103946 92568
rect 104345 92565 104357 92568
rect 104391 92565 104403 92599
rect 104345 92559 104403 92565
rect 1104 92506 7912 92528
rect 1104 92454 4874 92506
rect 4926 92454 4938 92506
rect 4990 92454 5002 92506
rect 5054 92454 5066 92506
rect 5118 92454 5130 92506
rect 5182 92454 7912 92506
rect 1104 92432 7912 92454
rect 104052 92506 108836 92528
rect 104052 92454 106658 92506
rect 106710 92454 106722 92506
rect 106774 92454 106786 92506
rect 106838 92454 106850 92506
rect 106902 92454 106914 92506
rect 106966 92454 108836 92506
rect 104052 92432 108836 92454
rect 1104 91962 7912 91984
rect 1104 91910 4214 91962
rect 4266 91910 4278 91962
rect 4330 91910 4342 91962
rect 4394 91910 4406 91962
rect 4458 91910 4470 91962
rect 4522 91910 7912 91962
rect 1104 91888 7912 91910
rect 104052 91962 108836 91984
rect 104052 91910 105922 91962
rect 105974 91910 105986 91962
rect 106038 91910 106050 91962
rect 106102 91910 106114 91962
rect 106166 91910 106178 91962
rect 106230 91910 108836 91962
rect 104052 91888 108836 91910
rect 104345 91579 104403 91585
rect 104345 91576 104357 91579
rect 103992 91548 104357 91576
rect 1104 91418 7912 91440
rect 1104 91366 4874 91418
rect 4926 91366 4938 91418
rect 4990 91366 5002 91418
rect 5054 91366 5066 91418
rect 5118 91366 5130 91418
rect 5182 91366 7912 91418
rect 1104 91344 7912 91366
rect 102778 91060 102784 91112
rect 102836 91100 102842 91112
rect 103992 91100 104020 91548
rect 104345 91545 104357 91548
rect 104391 91545 104403 91579
rect 104345 91539 104403 91545
rect 105078 91536 105084 91588
rect 105136 91576 105142 91588
rect 105357 91579 105415 91585
rect 105357 91576 105369 91579
rect 105136 91548 105369 91576
rect 105136 91536 105142 91548
rect 105357 91545 105369 91548
rect 105403 91545 105415 91579
rect 105357 91539 105415 91545
rect 104052 91418 108836 91440
rect 104052 91366 106658 91418
rect 106710 91366 106722 91418
rect 106774 91366 106786 91418
rect 106838 91366 106850 91418
rect 106902 91366 106914 91418
rect 106966 91366 108836 91418
rect 104052 91344 108836 91366
rect 104345 91103 104403 91109
rect 104345 91100 104357 91103
rect 102836 91072 104357 91100
rect 102836 91060 102842 91072
rect 104345 91069 104357 91072
rect 104391 91069 104403 91103
rect 104345 91063 104403 91069
rect 1104 90874 7912 90896
rect 1104 90822 4214 90874
rect 4266 90822 4278 90874
rect 4330 90822 4342 90874
rect 4394 90822 4406 90874
rect 4458 90822 4470 90874
rect 4522 90822 7912 90874
rect 1104 90800 7912 90822
rect 104052 90874 108836 90896
rect 104052 90822 105922 90874
rect 105974 90822 105986 90874
rect 106038 90822 106050 90874
rect 106102 90822 106114 90874
rect 106166 90822 106178 90874
rect 106230 90822 108836 90874
rect 104052 90800 108836 90822
rect 1104 90330 7912 90352
rect 1104 90278 4874 90330
rect 4926 90278 4938 90330
rect 4990 90278 5002 90330
rect 5054 90278 5066 90330
rect 5118 90278 5130 90330
rect 5182 90278 7912 90330
rect 1104 90256 7912 90278
rect 104052 90330 108836 90352
rect 104052 90278 106658 90330
rect 106710 90278 106722 90330
rect 106774 90278 106786 90330
rect 106838 90278 106850 90330
rect 106902 90278 106914 90330
rect 106966 90278 108836 90330
rect 104052 90256 108836 90278
rect 1104 89786 7912 89808
rect 1104 89734 4214 89786
rect 4266 89734 4278 89786
rect 4330 89734 4342 89786
rect 4394 89734 4406 89786
rect 4458 89734 4470 89786
rect 4522 89734 7912 89786
rect 1104 89712 7912 89734
rect 104052 89786 108836 89808
rect 104052 89734 105922 89786
rect 105974 89734 105986 89786
rect 106038 89734 106050 89786
rect 106102 89734 106114 89786
rect 106166 89734 106178 89786
rect 106230 89734 108836 89786
rect 104052 89712 108836 89734
rect 1104 89242 7912 89264
rect 1104 89190 4874 89242
rect 4926 89190 4938 89242
rect 4990 89190 5002 89242
rect 5054 89190 5066 89242
rect 5118 89190 5130 89242
rect 5182 89190 7912 89242
rect 1104 89168 7912 89190
rect 104052 89242 108836 89264
rect 104052 89190 106658 89242
rect 106710 89190 106722 89242
rect 106774 89190 106786 89242
rect 106838 89190 106850 89242
rect 106902 89190 106914 89242
rect 106966 89190 108836 89242
rect 104052 89168 108836 89190
rect 1302 88952 1308 89004
rect 1360 88992 1366 89004
rect 1489 88995 1547 89001
rect 1489 88992 1501 88995
rect 1360 88964 1501 88992
rect 1360 88952 1366 88964
rect 1489 88961 1501 88964
rect 1535 88992 1547 88995
rect 1949 88995 2007 89001
rect 1949 88992 1961 88995
rect 1535 88964 1961 88992
rect 1535 88961 1547 88964
rect 1489 88955 1547 88961
rect 1949 88961 1961 88964
rect 1995 88961 2007 88995
rect 1949 88955 2007 88961
rect 1673 88859 1731 88865
rect 1673 88825 1685 88859
rect 1719 88856 1731 88859
rect 1857 88859 1915 88865
rect 1857 88856 1869 88859
rect 1719 88828 1869 88856
rect 1719 88825 1731 88828
rect 1673 88819 1731 88825
rect 1857 88825 1869 88828
rect 1903 88856 1915 88859
rect 7558 88856 7564 88868
rect 1903 88828 7564 88856
rect 1903 88825 1915 88828
rect 1857 88819 1915 88825
rect 7558 88816 7564 88828
rect 7616 88816 7622 88868
rect 1104 88698 7912 88720
rect 1104 88646 4214 88698
rect 4266 88646 4278 88698
rect 4330 88646 4342 88698
rect 4394 88646 4406 88698
rect 4458 88646 4470 88698
rect 4522 88646 7912 88698
rect 1104 88624 7912 88646
rect 104052 88698 108836 88720
rect 104052 88646 105922 88698
rect 105974 88646 105986 88698
rect 106038 88646 106050 88698
rect 106102 88646 106114 88698
rect 106166 88646 106178 88698
rect 106230 88646 108836 88698
rect 104052 88624 108836 88646
rect 1104 88154 7912 88176
rect 1104 88102 4874 88154
rect 4926 88102 4938 88154
rect 4990 88102 5002 88154
rect 5054 88102 5066 88154
rect 5118 88102 5130 88154
rect 5182 88102 7912 88154
rect 1104 88080 7912 88102
rect 104052 88154 108836 88176
rect 104052 88102 106658 88154
rect 106710 88102 106722 88154
rect 106774 88102 106786 88154
rect 106838 88102 106850 88154
rect 106902 88102 106914 88154
rect 106966 88102 108836 88154
rect 104052 88080 108836 88102
rect 1210 87864 1216 87916
rect 1268 87904 1274 87916
rect 1489 87907 1547 87913
rect 1489 87904 1501 87907
rect 1268 87876 1501 87904
rect 1268 87864 1274 87876
rect 1489 87873 1501 87876
rect 1535 87904 1547 87907
rect 1949 87907 2007 87913
rect 1949 87904 1961 87907
rect 1535 87876 1961 87904
rect 1535 87873 1547 87876
rect 1489 87867 1547 87873
rect 1949 87873 1961 87876
rect 1995 87873 2007 87907
rect 1949 87867 2007 87873
rect 1673 87771 1731 87777
rect 1673 87737 1685 87771
rect 1719 87768 1731 87771
rect 1857 87771 1915 87777
rect 1857 87768 1869 87771
rect 1719 87740 1869 87768
rect 1719 87737 1731 87740
rect 1673 87731 1731 87737
rect 1857 87737 1869 87740
rect 1903 87768 1915 87771
rect 8938 87768 8944 87780
rect 1903 87740 8944 87768
rect 1903 87737 1915 87740
rect 1857 87731 1915 87737
rect 8938 87728 8944 87740
rect 8996 87728 9002 87780
rect 1104 87610 7912 87632
rect 1104 87558 4214 87610
rect 4266 87558 4278 87610
rect 4330 87558 4342 87610
rect 4394 87558 4406 87610
rect 4458 87558 4470 87610
rect 4522 87558 7912 87610
rect 1104 87536 7912 87558
rect 104052 87610 108836 87632
rect 104052 87558 105922 87610
rect 105974 87558 105986 87610
rect 106038 87558 106050 87610
rect 106102 87558 106114 87610
rect 106166 87558 106178 87610
rect 106230 87558 108836 87610
rect 104052 87536 108836 87558
rect 1210 87184 1216 87236
rect 1268 87224 1274 87236
rect 1489 87227 1547 87233
rect 1489 87224 1501 87227
rect 1268 87196 1501 87224
rect 1268 87184 1274 87196
rect 1489 87193 1501 87196
rect 1535 87224 1547 87227
rect 1949 87227 2007 87233
rect 1949 87224 1961 87227
rect 1535 87196 1961 87224
rect 1535 87193 1547 87196
rect 1489 87187 1547 87193
rect 1949 87193 1961 87196
rect 1995 87193 2007 87227
rect 1949 87187 2007 87193
rect 1581 87159 1639 87165
rect 1581 87125 1593 87159
rect 1627 87156 1639 87159
rect 1854 87156 1860 87168
rect 1627 87128 1860 87156
rect 1627 87125 1639 87128
rect 1581 87119 1639 87125
rect 1854 87116 1860 87128
rect 1912 87116 1918 87168
rect 1104 87066 7912 87088
rect 1104 87014 4874 87066
rect 4926 87014 4938 87066
rect 4990 87014 5002 87066
rect 5054 87014 5066 87066
rect 5118 87014 5130 87066
rect 5182 87014 7912 87066
rect 1104 86992 7912 87014
rect 104052 87066 108836 87088
rect 104052 87014 106658 87066
rect 106710 87014 106722 87066
rect 106774 87014 106786 87066
rect 106838 87014 106850 87066
rect 106902 87014 106914 87066
rect 106966 87014 108836 87066
rect 104052 86992 108836 87014
rect 1302 86776 1308 86828
rect 1360 86816 1366 86828
rect 1489 86819 1547 86825
rect 1489 86816 1501 86819
rect 1360 86788 1501 86816
rect 1360 86776 1366 86788
rect 1489 86785 1501 86788
rect 1535 86816 1547 86819
rect 1949 86819 2007 86825
rect 1949 86816 1961 86819
rect 1535 86788 1961 86816
rect 1535 86785 1547 86788
rect 1489 86779 1547 86785
rect 1949 86785 1961 86788
rect 1995 86785 2007 86819
rect 1949 86779 2007 86785
rect 1673 86683 1731 86689
rect 1673 86649 1685 86683
rect 1719 86680 1731 86683
rect 1857 86683 1915 86689
rect 1857 86680 1869 86683
rect 1719 86652 1869 86680
rect 1719 86649 1731 86652
rect 1673 86643 1731 86649
rect 1857 86649 1869 86652
rect 1903 86680 1915 86683
rect 8386 86680 8392 86692
rect 1903 86652 8392 86680
rect 1903 86649 1915 86652
rect 1857 86643 1915 86649
rect 8386 86640 8392 86652
rect 8444 86640 8450 86692
rect 1104 86522 7912 86544
rect 1104 86470 4214 86522
rect 4266 86470 4278 86522
rect 4330 86470 4342 86522
rect 4394 86470 4406 86522
rect 4458 86470 4470 86522
rect 4522 86470 7912 86522
rect 1104 86448 7912 86470
rect 104052 86522 108836 86544
rect 104052 86470 105922 86522
rect 105974 86470 105986 86522
rect 106038 86470 106050 86522
rect 106102 86470 106114 86522
rect 106166 86470 106178 86522
rect 106230 86470 108836 86522
rect 104052 86448 108836 86470
rect 1302 86164 1308 86216
rect 1360 86204 1366 86216
rect 1397 86207 1455 86213
rect 1397 86204 1409 86207
rect 1360 86176 1409 86204
rect 1360 86164 1366 86176
rect 1397 86173 1409 86176
rect 1443 86204 1455 86207
rect 1673 86207 1731 86213
rect 1673 86204 1685 86207
rect 1443 86176 1685 86204
rect 1443 86173 1455 86176
rect 1397 86167 1455 86173
rect 1673 86173 1685 86176
rect 1719 86173 1731 86207
rect 1673 86167 1731 86173
rect 1581 86071 1639 86077
rect 1581 86037 1593 86071
rect 1627 86068 1639 86071
rect 5534 86068 5540 86080
rect 1627 86040 5540 86068
rect 1627 86037 1639 86040
rect 1581 86031 1639 86037
rect 5534 86028 5540 86040
rect 5592 86028 5598 86080
rect 1104 85978 7912 86000
rect 1104 85926 4874 85978
rect 4926 85926 4938 85978
rect 4990 85926 5002 85978
rect 5054 85926 5066 85978
rect 5118 85926 5130 85978
rect 5182 85926 7912 85978
rect 1104 85904 7912 85926
rect 104052 85978 108836 86000
rect 104052 85926 106658 85978
rect 106710 85926 106722 85978
rect 106774 85926 106786 85978
rect 106838 85926 106850 85978
rect 106902 85926 106914 85978
rect 106966 85926 108836 85978
rect 104052 85904 108836 85926
rect 1854 85552 1860 85604
rect 1912 85592 1918 85604
rect 8570 85592 8576 85604
rect 1912 85564 8576 85592
rect 1912 85552 1918 85564
rect 8570 85552 8576 85564
rect 8628 85552 8634 85604
rect 1104 85434 7912 85456
rect 1104 85382 4214 85434
rect 4266 85382 4278 85434
rect 4330 85382 4342 85434
rect 4394 85382 4406 85434
rect 4458 85382 4470 85434
rect 4522 85382 7912 85434
rect 1104 85360 7912 85382
rect 104052 85434 108836 85456
rect 104052 85382 105922 85434
rect 105974 85382 105986 85434
rect 106038 85382 106050 85434
rect 106102 85382 106114 85434
rect 106166 85382 106178 85434
rect 106230 85382 108836 85434
rect 104052 85360 108836 85382
rect 1210 85008 1216 85060
rect 1268 85048 1274 85060
rect 1489 85051 1547 85057
rect 1489 85048 1501 85051
rect 1268 85020 1501 85048
rect 1268 85008 1274 85020
rect 1489 85017 1501 85020
rect 1535 85048 1547 85051
rect 1949 85051 2007 85057
rect 1949 85048 1961 85051
rect 1535 85020 1961 85048
rect 1535 85017 1547 85020
rect 1489 85011 1547 85017
rect 1949 85017 1961 85020
rect 1995 85017 2007 85051
rect 1949 85011 2007 85017
rect 1581 84983 1639 84989
rect 1581 84949 1593 84983
rect 1627 84980 1639 84983
rect 1857 84983 1915 84989
rect 1857 84980 1869 84983
rect 1627 84952 1869 84980
rect 1627 84949 1639 84952
rect 1581 84943 1639 84949
rect 1857 84949 1869 84952
rect 1903 84980 1915 84983
rect 2038 84980 2044 84992
rect 1903 84952 2044 84980
rect 1903 84949 1915 84952
rect 1857 84943 1915 84949
rect 2038 84940 2044 84952
rect 2096 84940 2102 84992
rect 1104 84890 7912 84912
rect 1104 84838 4874 84890
rect 4926 84838 4938 84890
rect 4990 84838 5002 84890
rect 5054 84838 5066 84890
rect 5118 84838 5130 84890
rect 5182 84838 7912 84890
rect 1104 84816 7912 84838
rect 104052 84890 108836 84912
rect 104052 84838 106658 84890
rect 106710 84838 106722 84890
rect 106774 84838 106786 84890
rect 106838 84838 106850 84890
rect 106902 84838 106914 84890
rect 106966 84838 108836 84890
rect 104052 84816 108836 84838
rect 1302 84600 1308 84652
rect 1360 84640 1366 84652
rect 1489 84643 1547 84649
rect 1489 84640 1501 84643
rect 1360 84612 1501 84640
rect 1360 84600 1366 84612
rect 1489 84609 1501 84612
rect 1535 84640 1547 84643
rect 1949 84643 2007 84649
rect 1949 84640 1961 84643
rect 1535 84612 1961 84640
rect 1535 84609 1547 84612
rect 1489 84603 1547 84609
rect 1949 84609 1961 84612
rect 1995 84609 2007 84643
rect 1949 84603 2007 84609
rect 1673 84507 1731 84513
rect 1673 84473 1685 84507
rect 1719 84504 1731 84507
rect 1765 84507 1823 84513
rect 1765 84504 1777 84507
rect 1719 84476 1777 84504
rect 1719 84473 1731 84476
rect 1673 84467 1731 84473
rect 1765 84473 1777 84476
rect 1811 84504 1823 84507
rect 1854 84504 1860 84516
rect 1811 84476 1860 84504
rect 1811 84473 1823 84476
rect 1765 84467 1823 84473
rect 1854 84464 1860 84476
rect 1912 84464 1918 84516
rect 1104 84346 7912 84368
rect 1104 84294 4214 84346
rect 4266 84294 4278 84346
rect 4330 84294 4342 84346
rect 4394 84294 4406 84346
rect 4458 84294 4470 84346
rect 4522 84294 7912 84346
rect 1104 84272 7912 84294
rect 104052 84346 108836 84368
rect 104052 84294 105922 84346
rect 105974 84294 105986 84346
rect 106038 84294 106050 84346
rect 106102 84294 106114 84346
rect 106166 84294 106178 84346
rect 106230 84294 108836 84346
rect 104052 84272 108836 84294
rect 1854 84124 1860 84176
rect 1912 84164 1918 84176
rect 9306 84164 9312 84176
rect 1912 84136 9312 84164
rect 1912 84124 1918 84136
rect 9306 84124 9312 84136
rect 9364 84124 9370 84176
rect 1302 83988 1308 84040
rect 1360 84028 1366 84040
rect 1397 84031 1455 84037
rect 1397 84028 1409 84031
rect 1360 84000 1409 84028
rect 1360 83988 1366 84000
rect 1397 83997 1409 84000
rect 1443 84028 1455 84031
rect 1949 84031 2007 84037
rect 1949 84028 1961 84031
rect 1443 84000 1961 84028
rect 1443 83997 1455 84000
rect 1397 83991 1455 83997
rect 1949 83997 1961 84000
rect 1995 83997 2007 84031
rect 1949 83991 2007 83997
rect 1581 83895 1639 83901
rect 1581 83861 1593 83895
rect 1627 83892 1639 83895
rect 1857 83895 1915 83901
rect 1857 83892 1869 83895
rect 1627 83864 1869 83892
rect 1627 83861 1639 83864
rect 1581 83855 1639 83861
rect 1857 83861 1869 83864
rect 1903 83892 1915 83895
rect 2498 83892 2504 83904
rect 1903 83864 2504 83892
rect 1903 83861 1915 83864
rect 1857 83855 1915 83861
rect 2498 83852 2504 83864
rect 2556 83852 2562 83904
rect 1104 83802 7912 83824
rect 1104 83750 4874 83802
rect 4926 83750 4938 83802
rect 4990 83750 5002 83802
rect 5054 83750 5066 83802
rect 5118 83750 5130 83802
rect 5182 83750 7912 83802
rect 1104 83728 7912 83750
rect 104052 83802 108836 83824
rect 104052 83750 106658 83802
rect 106710 83750 106722 83802
rect 106774 83750 106786 83802
rect 106838 83750 106850 83802
rect 106902 83750 106914 83802
rect 106966 83750 108836 83802
rect 104052 83728 108836 83750
rect 1302 83512 1308 83564
rect 1360 83552 1366 83564
rect 1489 83555 1547 83561
rect 1489 83552 1501 83555
rect 1360 83524 1501 83552
rect 1360 83512 1366 83524
rect 1489 83521 1501 83524
rect 1535 83552 1547 83555
rect 1949 83555 2007 83561
rect 1949 83552 1961 83555
rect 1535 83524 1961 83552
rect 1535 83521 1547 83524
rect 1489 83515 1547 83521
rect 1949 83521 1961 83524
rect 1995 83521 2007 83555
rect 1949 83515 2007 83521
rect 2038 83444 2044 83496
rect 2096 83484 2102 83496
rect 9214 83484 9220 83496
rect 2096 83456 9220 83484
rect 2096 83444 2102 83456
rect 9214 83444 9220 83456
rect 9272 83444 9278 83496
rect 1581 83351 1639 83357
rect 1581 83317 1593 83351
rect 1627 83348 1639 83351
rect 1857 83351 1915 83357
rect 1857 83348 1869 83351
rect 1627 83320 1869 83348
rect 1627 83317 1639 83320
rect 1581 83311 1639 83317
rect 1857 83317 1869 83320
rect 1903 83348 1915 83351
rect 2038 83348 2044 83360
rect 1903 83320 2044 83348
rect 1903 83317 1915 83320
rect 1857 83311 1915 83317
rect 2038 83308 2044 83320
rect 2096 83308 2102 83360
rect 1104 83258 7912 83280
rect 1104 83206 4214 83258
rect 4266 83206 4278 83258
rect 4330 83206 4342 83258
rect 4394 83206 4406 83258
rect 4458 83206 4470 83258
rect 4522 83206 7912 83258
rect 1104 83184 7912 83206
rect 104052 83258 108836 83280
rect 104052 83206 105922 83258
rect 105974 83206 105986 83258
rect 106038 83206 106050 83258
rect 106102 83206 106114 83258
rect 106166 83206 106178 83258
rect 106230 83206 108836 83258
rect 104052 83184 108836 83206
rect 1104 82714 7912 82736
rect 1104 82662 4874 82714
rect 4926 82662 4938 82714
rect 4990 82662 5002 82714
rect 5054 82662 5066 82714
rect 5118 82662 5130 82714
rect 5182 82662 7912 82714
rect 1104 82640 7912 82662
rect 104052 82714 108836 82736
rect 104052 82662 106658 82714
rect 106710 82662 106722 82714
rect 106774 82662 106786 82714
rect 106838 82662 106850 82714
rect 106902 82662 106914 82714
rect 106966 82662 108836 82714
rect 104052 82640 108836 82662
rect 1210 82424 1216 82476
rect 1268 82464 1274 82476
rect 1489 82467 1547 82473
rect 1489 82464 1501 82467
rect 1268 82436 1501 82464
rect 1268 82424 1274 82436
rect 1489 82433 1501 82436
rect 1535 82464 1547 82467
rect 1949 82467 2007 82473
rect 1949 82464 1961 82467
rect 1535 82436 1961 82464
rect 1535 82433 1547 82436
rect 1489 82427 1547 82433
rect 1949 82433 1961 82436
rect 1995 82433 2007 82467
rect 1949 82427 2007 82433
rect 4985 82467 5043 82473
rect 4985 82433 4997 82467
rect 5031 82464 5043 82467
rect 5031 82436 5212 82464
rect 5031 82433 5043 82436
rect 4985 82427 5043 82433
rect 5184 82405 5212 82436
rect 4249 82399 4307 82405
rect 4249 82365 4261 82399
rect 4295 82365 4307 82399
rect 4249 82359 4307 82365
rect 5169 82399 5227 82405
rect 5169 82365 5181 82399
rect 5215 82396 5227 82399
rect 5258 82396 5264 82408
rect 5215 82368 5264 82396
rect 5215 82365 5227 82368
rect 5169 82359 5227 82365
rect 1581 82263 1639 82269
rect 1581 82229 1593 82263
rect 1627 82260 1639 82263
rect 1857 82263 1915 82269
rect 1857 82260 1869 82263
rect 1627 82232 1869 82260
rect 1627 82229 1639 82232
rect 1581 82223 1639 82229
rect 1857 82229 1869 82232
rect 1903 82260 1915 82263
rect 2682 82260 2688 82272
rect 1903 82232 2688 82260
rect 1903 82229 1915 82232
rect 1857 82223 1915 82229
rect 2682 82220 2688 82232
rect 2740 82220 2746 82272
rect 4264 82260 4292 82359
rect 5258 82356 5264 82368
rect 5316 82356 5322 82408
rect 5353 82263 5411 82269
rect 5353 82260 5365 82263
rect 4264 82232 5365 82260
rect 5353 82229 5365 82232
rect 5399 82260 5411 82263
rect 5810 82260 5816 82272
rect 5399 82232 5816 82260
rect 5399 82229 5411 82232
rect 5353 82223 5411 82229
rect 5810 82220 5816 82232
rect 5868 82260 5874 82272
rect 6178 82260 6184 82272
rect 5868 82232 6184 82260
rect 5868 82220 5874 82232
rect 6178 82220 6184 82232
rect 6236 82220 6242 82272
rect 1104 82170 7912 82192
rect 1104 82118 4214 82170
rect 4266 82118 4278 82170
rect 4330 82118 4342 82170
rect 4394 82118 4406 82170
rect 4458 82118 4470 82170
rect 4522 82118 7912 82170
rect 1104 82096 7912 82118
rect 104052 82170 108836 82192
rect 104052 82118 105922 82170
rect 105974 82118 105986 82170
rect 106038 82118 106050 82170
rect 106102 82118 106114 82170
rect 106166 82118 106178 82170
rect 106230 82118 108836 82170
rect 104052 82096 108836 82118
rect 1210 81744 1216 81796
rect 1268 81784 1274 81796
rect 1489 81787 1547 81793
rect 1489 81784 1501 81787
rect 1268 81756 1501 81784
rect 1268 81744 1274 81756
rect 1489 81753 1501 81756
rect 1535 81784 1547 81787
rect 1949 81787 2007 81793
rect 1949 81784 1961 81787
rect 1535 81756 1961 81784
rect 1535 81753 1547 81756
rect 1489 81747 1547 81753
rect 1949 81753 1961 81756
rect 1995 81753 2007 81787
rect 1949 81747 2007 81753
rect 1581 81719 1639 81725
rect 1581 81685 1593 81719
rect 1627 81716 1639 81719
rect 1854 81716 1860 81728
rect 1627 81688 1860 81716
rect 1627 81685 1639 81688
rect 1581 81679 1639 81685
rect 1854 81676 1860 81688
rect 1912 81676 1918 81728
rect 1104 81626 7912 81648
rect 1104 81574 4874 81626
rect 4926 81574 4938 81626
rect 4990 81574 5002 81626
rect 5054 81574 5066 81626
rect 5118 81574 5130 81626
rect 5182 81574 7912 81626
rect 1104 81552 7912 81574
rect 104052 81626 108836 81648
rect 104052 81574 106658 81626
rect 106710 81574 106722 81626
rect 106774 81574 106786 81626
rect 106838 81574 106850 81626
rect 106902 81574 106914 81626
rect 106966 81574 108836 81626
rect 104052 81552 108836 81574
rect 1302 81336 1308 81388
rect 1360 81376 1366 81388
rect 1489 81379 1547 81385
rect 1489 81376 1501 81379
rect 1360 81348 1501 81376
rect 1360 81336 1366 81348
rect 1489 81345 1501 81348
rect 1535 81376 1547 81379
rect 1949 81379 2007 81385
rect 1949 81376 1961 81379
rect 1535 81348 1961 81376
rect 1535 81345 1547 81348
rect 1489 81339 1547 81345
rect 1949 81345 1961 81348
rect 1995 81345 2007 81379
rect 1949 81339 2007 81345
rect 2038 81268 2044 81320
rect 2096 81308 2102 81320
rect 9766 81308 9772 81320
rect 2096 81280 9772 81308
rect 2096 81268 2102 81280
rect 9766 81268 9772 81280
rect 9824 81268 9830 81320
rect 1673 81243 1731 81249
rect 1673 81209 1685 81243
rect 1719 81240 1731 81243
rect 1857 81243 1915 81249
rect 1857 81240 1869 81243
rect 1719 81212 1869 81240
rect 1719 81209 1731 81212
rect 1673 81203 1731 81209
rect 1857 81209 1869 81212
rect 1903 81240 1915 81243
rect 9582 81240 9588 81252
rect 1903 81212 9588 81240
rect 1903 81209 1915 81212
rect 1857 81203 1915 81209
rect 9582 81200 9588 81212
rect 9640 81200 9646 81252
rect 1104 81082 7912 81104
rect 1104 81030 4214 81082
rect 4266 81030 4278 81082
rect 4330 81030 4342 81082
rect 4394 81030 4406 81082
rect 4458 81030 4470 81082
rect 4522 81030 7912 81082
rect 1104 81008 7912 81030
rect 104052 81082 108836 81104
rect 104052 81030 105922 81082
rect 105974 81030 105986 81082
rect 106038 81030 106050 81082
rect 106102 81030 106114 81082
rect 106166 81030 106178 81082
rect 106230 81030 108836 81082
rect 104052 81008 108836 81030
rect 1854 80792 1860 80844
rect 1912 80832 1918 80844
rect 9674 80832 9680 80844
rect 1912 80804 9680 80832
rect 1912 80792 1918 80804
rect 9674 80792 9680 80804
rect 9732 80792 9738 80844
rect 1302 80724 1308 80776
rect 1360 80764 1366 80776
rect 1397 80767 1455 80773
rect 1397 80764 1409 80767
rect 1360 80736 1409 80764
rect 1360 80724 1366 80736
rect 1397 80733 1409 80736
rect 1443 80733 1455 80767
rect 1397 80727 1455 80733
rect 1673 80767 1731 80773
rect 1673 80733 1685 80767
rect 1719 80764 1731 80767
rect 1719 80736 2452 80764
rect 1719 80733 1731 80736
rect 1673 80727 1731 80733
rect 2424 80637 2452 80736
rect 2682 80724 2688 80776
rect 2740 80764 2746 80776
rect 9858 80764 9864 80776
rect 2740 80736 9864 80764
rect 2740 80724 2746 80736
rect 9858 80724 9864 80736
rect 9916 80724 9922 80776
rect 107746 80724 107752 80776
rect 107804 80764 107810 80776
rect 108209 80767 108267 80773
rect 108209 80764 108221 80767
rect 107804 80736 108221 80764
rect 107804 80724 107810 80736
rect 108209 80733 108221 80736
rect 108255 80733 108267 80767
rect 108209 80727 108267 80733
rect 108482 80724 108488 80776
rect 108540 80724 108546 80776
rect 2498 80656 2504 80708
rect 2556 80696 2562 80708
rect 9950 80696 9956 80708
rect 2556 80668 9956 80696
rect 2556 80656 2562 80668
rect 9950 80656 9956 80668
rect 10008 80656 10014 80708
rect 2409 80631 2467 80637
rect 2409 80597 2421 80631
rect 2455 80628 2467 80631
rect 5534 80628 5540 80640
rect 2455 80600 5540 80628
rect 2455 80597 2467 80600
rect 2409 80591 2467 80597
rect 5534 80588 5540 80600
rect 5592 80588 5598 80640
rect 1104 80538 7912 80560
rect 1104 80486 4874 80538
rect 4926 80486 4938 80538
rect 4990 80486 5002 80538
rect 5054 80486 5066 80538
rect 5118 80486 5130 80538
rect 5182 80486 7912 80538
rect 1104 80464 7912 80486
rect 104052 80538 108836 80560
rect 104052 80486 106658 80538
rect 106710 80486 106722 80538
rect 106774 80486 106786 80538
rect 106838 80486 106850 80538
rect 106902 80486 106914 80538
rect 106966 80486 108836 80538
rect 104052 80464 108836 80486
rect 1302 80316 1308 80368
rect 1360 80356 1366 80368
rect 1397 80359 1455 80365
rect 1397 80356 1409 80359
rect 1360 80328 1409 80356
rect 1360 80316 1366 80328
rect 1397 80325 1409 80328
rect 1443 80325 1455 80359
rect 1397 80319 1455 80325
rect 108482 80316 108488 80368
rect 108540 80316 108546 80368
rect 101950 80044 101956 80096
rect 102008 80084 102014 80096
rect 105814 80084 105820 80096
rect 102008 80056 105820 80084
rect 102008 80044 102014 80056
rect 105814 80044 105820 80056
rect 105872 80044 105878 80096
rect 1104 79994 7912 80016
rect 1104 79942 4214 79994
rect 4266 79942 4278 79994
rect 4330 79942 4342 79994
rect 4394 79942 4406 79994
rect 4458 79942 4470 79994
rect 4522 79942 7912 79994
rect 9950 79976 9956 80028
rect 10008 80016 10014 80028
rect 43254 80016 43260 80028
rect 10008 79988 43260 80016
rect 10008 79976 10014 79988
rect 43254 79976 43260 79988
rect 43312 79976 43318 80028
rect 104052 79994 108836 80016
rect 1104 79920 7912 79942
rect 9766 79908 9772 79960
rect 9824 79948 9830 79960
rect 40954 79948 40960 79960
rect 9824 79920 40960 79948
rect 9824 79908 9830 79920
rect 40954 79908 40960 79920
rect 41012 79908 41018 79960
rect 104052 79942 105922 79994
rect 105974 79942 105986 79994
rect 106038 79942 106050 79994
rect 106102 79942 106114 79994
rect 106166 79942 106178 79994
rect 106230 79942 108836 79994
rect 104052 79920 108836 79942
rect 9858 79840 9864 79892
rect 9916 79880 9922 79892
rect 39758 79880 39764 79892
rect 9916 79852 39764 79880
rect 9916 79840 9922 79852
rect 39758 79840 39764 79852
rect 39816 79840 39822 79892
rect 7558 79772 7564 79824
rect 7616 79812 7622 79824
rect 36262 79812 36268 79824
rect 7616 79784 36268 79812
rect 7616 79772 7622 79784
rect 36262 79772 36268 79784
rect 36320 79772 36326 79824
rect 9674 79704 9680 79756
rect 9732 79744 9738 79756
rect 38654 79744 38660 79756
rect 9732 79716 38660 79744
rect 9732 79704 9738 79716
rect 38654 79704 38660 79716
rect 38712 79704 38718 79756
rect 8938 79636 8944 79688
rect 8996 79676 9002 79688
rect 33962 79676 33968 79688
rect 8996 79648 33968 79676
rect 8996 79636 9002 79648
rect 33962 79636 33968 79648
rect 34020 79636 34026 79688
rect 97994 79636 98000 79688
rect 98052 79676 98058 79688
rect 108209 79679 108267 79685
rect 108209 79676 108221 79679
rect 98052 79648 108221 79676
rect 98052 79636 98058 79648
rect 108209 79645 108221 79648
rect 108255 79645 108267 79679
rect 108209 79639 108267 79645
rect 1210 79568 1216 79620
rect 1268 79608 1274 79620
rect 1489 79611 1547 79617
rect 1489 79608 1501 79611
rect 1268 79580 1501 79608
rect 1268 79568 1274 79580
rect 1489 79577 1501 79580
rect 1535 79577 1547 79611
rect 1489 79571 1547 79577
rect 1673 79611 1731 79617
rect 1673 79577 1685 79611
rect 1719 79608 1731 79611
rect 1857 79611 1915 79617
rect 1857 79608 1869 79611
rect 1719 79580 1869 79608
rect 1719 79577 1731 79580
rect 1673 79571 1731 79577
rect 1857 79577 1869 79580
rect 1903 79608 1915 79611
rect 1903 79580 6914 79608
rect 1903 79577 1915 79580
rect 1857 79571 1915 79577
rect 1504 79540 1532 79571
rect 1949 79543 2007 79549
rect 1949 79540 1961 79543
rect 1504 79512 1961 79540
rect 1949 79509 1961 79512
rect 1995 79509 2007 79543
rect 6886 79540 6914 79580
rect 8570 79568 8576 79620
rect 8628 79608 8634 79620
rect 31662 79608 31668 79620
rect 8628 79580 31668 79608
rect 8628 79568 8634 79580
rect 31662 79568 31668 79580
rect 31720 79568 31726 79620
rect 37458 79540 37464 79552
rect 6886 79512 37464 79540
rect 1949 79503 2007 79509
rect 37458 79500 37464 79512
rect 37516 79500 37522 79552
rect 108390 79500 108396 79552
rect 108448 79500 108454 79552
rect 1104 79450 7912 79472
rect 1104 79398 4874 79450
rect 4926 79398 4938 79450
rect 4990 79398 5002 79450
rect 5054 79398 5066 79450
rect 5118 79398 5130 79450
rect 5182 79398 7912 79450
rect 92106 79432 92112 79484
rect 92164 79472 92170 79484
rect 102870 79472 102876 79484
rect 92164 79444 102876 79472
rect 92164 79432 92170 79444
rect 102870 79432 102876 79444
rect 102928 79432 102934 79484
rect 104052 79450 108836 79472
rect 1104 79376 7912 79398
rect 90266 79364 90272 79416
rect 90324 79404 90330 79416
rect 102962 79404 102968 79416
rect 90324 79376 102968 79404
rect 90324 79364 90330 79376
rect 102962 79364 102968 79376
rect 103020 79364 103026 79416
rect 104052 79398 106658 79450
rect 106710 79398 106722 79450
rect 106774 79398 106786 79450
rect 106838 79398 106850 79450
rect 106902 79398 106914 79450
rect 106966 79398 108836 79450
rect 104052 79376 108836 79398
rect 73798 79296 73804 79348
rect 73856 79336 73862 79348
rect 102778 79336 102784 79348
rect 73856 79308 102784 79336
rect 73856 79296 73862 79308
rect 102778 79296 102784 79308
rect 102836 79296 102842 79348
rect 1302 79160 1308 79212
rect 1360 79200 1366 79212
rect 1489 79203 1547 79209
rect 1489 79200 1501 79203
rect 1360 79172 1501 79200
rect 1360 79160 1366 79172
rect 1489 79169 1501 79172
rect 1535 79200 1547 79203
rect 1949 79203 2007 79209
rect 1949 79200 1961 79203
rect 1535 79172 1961 79200
rect 1535 79169 1547 79172
rect 1489 79163 1547 79169
rect 1949 79169 1961 79172
rect 1995 79169 2007 79203
rect 1949 79163 2007 79169
rect 96798 79160 96804 79212
rect 96856 79200 96862 79212
rect 108209 79203 108267 79209
rect 108209 79200 108221 79203
rect 96856 79172 108221 79200
rect 96856 79160 96862 79172
rect 108209 79169 108221 79172
rect 108255 79169 108267 79203
rect 108209 79163 108267 79169
rect 1673 79067 1731 79073
rect 1673 79033 1685 79067
rect 1719 79064 1731 79067
rect 1857 79067 1915 79073
rect 1857 79064 1869 79067
rect 1719 79036 1869 79064
rect 1719 79033 1731 79036
rect 1673 79027 1731 79033
rect 1857 79033 1869 79036
rect 1903 79064 1915 79067
rect 1903 79036 6914 79064
rect 1903 79033 1915 79036
rect 1857 79027 1915 79033
rect 6886 78996 6914 79036
rect 42150 78996 42156 79008
rect 6886 78968 42156 78996
rect 42150 78956 42156 78968
rect 42208 78956 42214 79008
rect 108390 78956 108396 79008
rect 108448 78956 108454 79008
rect 1104 78906 7912 78928
rect 1104 78854 4214 78906
rect 4266 78854 4278 78906
rect 4330 78854 4342 78906
rect 4394 78854 4406 78906
rect 4458 78854 4470 78906
rect 4522 78854 7912 78906
rect 1104 78832 7912 78854
rect 104052 78906 108836 78928
rect 104052 78854 105922 78906
rect 105974 78854 105986 78906
rect 106038 78854 106050 78906
rect 106102 78854 106114 78906
rect 106166 78854 106178 78906
rect 106230 78854 108836 78906
rect 104052 78832 108836 78854
rect 7282 78616 7288 78668
rect 7340 78656 7346 78668
rect 13998 78656 14004 78668
rect 7340 78628 14004 78656
rect 7340 78616 7346 78628
rect 13998 78616 14004 78628
rect 14056 78616 14062 78668
rect 95878 78616 95884 78668
rect 95936 78656 95942 78668
rect 102042 78656 102048 78668
rect 95936 78628 102048 78656
rect 95936 78616 95942 78628
rect 102042 78616 102048 78628
rect 102100 78616 102106 78668
rect 107654 78548 107660 78600
rect 107712 78588 107718 78600
rect 108209 78591 108267 78597
rect 108209 78588 108221 78591
rect 107712 78560 108221 78588
rect 107712 78548 107718 78560
rect 108209 78557 108221 78560
rect 108255 78557 108267 78591
rect 108209 78551 108267 78557
rect 1302 78480 1308 78532
rect 1360 78520 1366 78532
rect 1489 78523 1547 78529
rect 1489 78520 1501 78523
rect 1360 78492 1501 78520
rect 1360 78480 1366 78492
rect 1489 78489 1501 78492
rect 1535 78489 1547 78523
rect 1489 78483 1547 78489
rect 1673 78523 1731 78529
rect 1673 78489 1685 78523
rect 1719 78520 1731 78523
rect 1857 78523 1915 78529
rect 1857 78520 1869 78523
rect 1719 78492 1869 78520
rect 1719 78489 1731 78492
rect 1673 78483 1731 78489
rect 1857 78489 1869 78492
rect 1903 78520 1915 78523
rect 1903 78492 6914 78520
rect 1903 78489 1915 78492
rect 1857 78483 1915 78489
rect 1504 78452 1532 78483
rect 1949 78455 2007 78461
rect 1949 78452 1961 78455
rect 1504 78424 1961 78452
rect 1949 78421 1961 78424
rect 1995 78421 2007 78455
rect 6886 78452 6914 78492
rect 29546 78452 29552 78464
rect 6886 78424 29552 78452
rect 1949 78415 2007 78421
rect 29546 78412 29552 78424
rect 29604 78412 29610 78464
rect 108390 78412 108396 78464
rect 108448 78412 108454 78464
rect 1104 78362 7912 78384
rect 1104 78310 4874 78362
rect 4926 78310 4938 78362
rect 4990 78310 5002 78362
rect 5054 78310 5066 78362
rect 5118 78310 5130 78362
rect 5182 78310 7912 78362
rect 1104 78288 7912 78310
rect 104052 78362 108836 78384
rect 104052 78310 106658 78362
rect 106710 78310 106722 78362
rect 106774 78310 106786 78362
rect 106838 78310 106850 78362
rect 106902 78310 106914 78362
rect 106966 78310 108836 78362
rect 104052 78288 108836 78310
rect 91922 78140 91928 78192
rect 91980 78180 91986 78192
rect 102318 78180 102324 78192
rect 91980 78152 102324 78180
rect 91980 78140 91986 78152
rect 102318 78140 102324 78152
rect 102376 78140 102382 78192
rect 1302 78072 1308 78124
rect 1360 78112 1366 78124
rect 1489 78115 1547 78121
rect 1489 78112 1501 78115
rect 1360 78084 1501 78112
rect 1360 78072 1366 78084
rect 1489 78081 1501 78084
rect 1535 78112 1547 78115
rect 1949 78115 2007 78121
rect 1949 78112 1961 78115
rect 1535 78084 1961 78112
rect 1535 78081 1547 78084
rect 1489 78075 1547 78081
rect 1949 78081 1961 78084
rect 1995 78081 2007 78115
rect 1949 78075 2007 78081
rect 2038 78072 2044 78124
rect 2096 78112 2102 78124
rect 35342 78112 35348 78124
rect 2096 78084 35348 78112
rect 2096 78072 2102 78084
rect 35342 78072 35348 78084
rect 35400 78072 35406 78124
rect 108206 78072 108212 78124
rect 108264 78072 108270 78124
rect 16206 78004 16212 78056
rect 16264 78044 16270 78056
rect 25406 78044 25412 78056
rect 16264 78016 25412 78044
rect 16264 78004 16270 78016
rect 25406 78004 25412 78016
rect 25464 78004 25470 78056
rect 92382 78004 92388 78056
rect 92440 78044 92446 78056
rect 102410 78044 102416 78056
rect 92440 78016 102416 78044
rect 92440 78004 92446 78016
rect 102410 78004 102416 78016
rect 102468 78004 102474 78056
rect 1673 77979 1731 77985
rect 1673 77945 1685 77979
rect 1719 77976 1731 77979
rect 1857 77979 1915 77985
rect 1857 77976 1869 77979
rect 1719 77948 1869 77976
rect 1719 77945 1731 77948
rect 1673 77939 1731 77945
rect 1857 77945 1869 77948
rect 1903 77976 1915 77979
rect 1903 77948 6914 77976
rect 1903 77945 1915 77948
rect 1857 77939 1915 77945
rect 6886 77908 6914 77948
rect 7098 77936 7104 77988
rect 7156 77976 7162 77988
rect 17126 77976 17132 77988
rect 7156 77948 17132 77976
rect 7156 77936 7162 77948
rect 17126 77936 17132 77948
rect 17184 77936 17190 77988
rect 89898 77936 89904 77988
rect 89956 77976 89962 77988
rect 102134 77976 102140 77988
rect 89956 77948 102140 77976
rect 89956 77936 89962 77948
rect 102134 77936 102140 77948
rect 102192 77936 102198 77988
rect 26050 77908 26056 77920
rect 6886 77880 26056 77908
rect 26050 77868 26056 77880
rect 26108 77868 26114 77920
rect 87230 77868 87236 77920
rect 87288 77908 87294 77920
rect 101950 77908 101956 77920
rect 87288 77880 101956 77908
rect 87288 77868 87294 77880
rect 101950 77868 101956 77880
rect 102008 77868 102014 77920
rect 108390 77868 108396 77920
rect 108448 77868 108454 77920
rect 1104 77818 108836 77840
rect 1104 77766 4214 77818
rect 4266 77766 4278 77818
rect 4330 77766 4342 77818
rect 4394 77766 4406 77818
rect 4458 77766 4470 77818
rect 4522 77766 34934 77818
rect 34986 77766 34998 77818
rect 35050 77766 35062 77818
rect 35114 77766 35126 77818
rect 35178 77766 35190 77818
rect 35242 77766 65654 77818
rect 65706 77766 65718 77818
rect 65770 77766 65782 77818
rect 65834 77766 65846 77818
rect 65898 77766 65910 77818
rect 65962 77766 96374 77818
rect 96426 77766 96438 77818
rect 96490 77766 96502 77818
rect 96554 77766 96566 77818
rect 96618 77766 96630 77818
rect 96682 77766 105922 77818
rect 105974 77766 105986 77818
rect 106038 77766 106050 77818
rect 106102 77766 106114 77818
rect 106166 77766 106178 77818
rect 106230 77766 108836 77818
rect 1104 77744 108836 77766
rect 8018 77664 8024 77716
rect 8076 77704 8082 77716
rect 8076 77676 15240 77704
rect 8076 77664 8082 77676
rect 11054 77596 11060 77648
rect 11112 77636 11118 77648
rect 14737 77639 14795 77645
rect 14737 77636 14749 77639
rect 11112 77608 14749 77636
rect 11112 77596 11118 77608
rect 14737 77605 14749 77608
rect 14783 77605 14795 77639
rect 14737 77599 14795 77605
rect 15212 77568 15240 77676
rect 16114 77664 16120 77716
rect 16172 77704 16178 77716
rect 16669 77707 16727 77713
rect 16669 77704 16681 77707
rect 16172 77676 16681 77704
rect 16172 77664 16178 77676
rect 16669 77673 16681 77676
rect 16715 77673 16727 77707
rect 16669 77667 16727 77673
rect 26050 77664 26056 77716
rect 26108 77664 26114 77716
rect 26970 77664 26976 77716
rect 27028 77664 27034 77716
rect 28166 77664 28172 77716
rect 28224 77664 28230 77716
rect 29546 77664 29552 77716
rect 29604 77664 29610 77716
rect 30466 77664 30472 77716
rect 30524 77664 30530 77716
rect 31754 77664 31760 77716
rect 31812 77664 31818 77716
rect 32858 77664 32864 77716
rect 32916 77664 32922 77716
rect 33962 77664 33968 77716
rect 34020 77664 34026 77716
rect 35253 77707 35311 77713
rect 35253 77673 35265 77707
rect 35299 77704 35311 77707
rect 35342 77704 35348 77716
rect 35299 77676 35348 77704
rect 35299 77673 35311 77676
rect 35253 77667 35311 77673
rect 35342 77664 35348 77676
rect 35400 77664 35406 77716
rect 36262 77664 36268 77716
rect 36320 77704 36326 77716
rect 36357 77707 36415 77713
rect 36357 77704 36369 77707
rect 36320 77676 36369 77704
rect 36320 77664 36326 77676
rect 36357 77673 36369 77676
rect 36403 77673 36415 77707
rect 36357 77667 36415 77673
rect 37458 77664 37464 77716
rect 37516 77664 37522 77716
rect 38654 77664 38660 77716
rect 38712 77664 38718 77716
rect 39758 77664 39764 77716
rect 39816 77704 39822 77716
rect 39853 77707 39911 77713
rect 39853 77704 39865 77707
rect 39816 77676 39865 77704
rect 39816 77664 39822 77676
rect 39853 77673 39865 77676
rect 39899 77673 39911 77707
rect 39853 77667 39911 77673
rect 40954 77664 40960 77716
rect 41012 77704 41018 77716
rect 41049 77707 41107 77713
rect 41049 77704 41061 77707
rect 41012 77676 41061 77704
rect 41012 77664 41018 77676
rect 41049 77673 41061 77676
rect 41095 77673 41107 77707
rect 41049 77667 41107 77673
rect 42150 77664 42156 77716
rect 42208 77664 42214 77716
rect 43254 77664 43260 77716
rect 43312 77704 43318 77716
rect 43349 77707 43407 77713
rect 43349 77704 43361 77707
rect 43312 77676 43361 77704
rect 43312 77664 43318 77676
rect 43349 77673 43361 77676
rect 43395 77673 43407 77707
rect 43349 77667 43407 77673
rect 91186 77664 91192 77716
rect 91244 77704 91250 77716
rect 94866 77704 94872 77716
rect 91244 77676 94872 77704
rect 91244 77664 91250 77676
rect 94866 77664 94872 77676
rect 94924 77664 94930 77716
rect 94961 77707 95019 77713
rect 94961 77673 94973 77707
rect 95007 77704 95019 77707
rect 97902 77704 97908 77716
rect 95007 77676 97908 77704
rect 95007 77673 95019 77676
rect 94961 77667 95019 77673
rect 97902 77664 97908 77676
rect 97960 77664 97966 77716
rect 99098 77664 99104 77716
rect 99156 77704 99162 77716
rect 104342 77704 104348 77716
rect 99156 77676 104348 77704
rect 99156 77664 99162 77676
rect 104342 77664 104348 77676
rect 104400 77664 104406 77716
rect 25777 77639 25835 77645
rect 25777 77605 25789 77639
rect 25823 77636 25835 77639
rect 27522 77636 27528 77648
rect 25823 77608 27528 77636
rect 25823 77605 25835 77608
rect 25777 77599 25835 77605
rect 27522 77596 27528 77608
rect 27580 77596 27586 77648
rect 87230 77636 87236 77648
rect 86604 77608 87236 77636
rect 83737 77571 83795 77577
rect 83737 77568 83749 77571
rect 15212 77540 24532 77568
rect 16485 77503 16543 77509
rect 16485 77469 16497 77503
rect 16531 77500 16543 77503
rect 19886 77500 19892 77512
rect 16531 77472 19892 77500
rect 16531 77469 16543 77472
rect 16485 77463 16543 77469
rect 19886 77460 19892 77472
rect 19944 77500 19950 77512
rect 24121 77503 24179 77509
rect 24121 77500 24133 77503
rect 19944 77472 24133 77500
rect 19944 77460 19950 77472
rect 24121 77469 24133 77472
rect 24167 77500 24179 77503
rect 24397 77503 24455 77509
rect 24397 77500 24409 77503
rect 24167 77472 24409 77500
rect 24167 77469 24179 77472
rect 24121 77463 24179 77469
rect 24397 77469 24409 77472
rect 24443 77469 24455 77503
rect 24504 77500 24532 77540
rect 83384 77540 83749 77568
rect 24653 77503 24711 77509
rect 24653 77500 24665 77503
rect 24504 77472 24665 77500
rect 24397 77463 24455 77469
rect 24653 77469 24665 77472
rect 24699 77500 24711 77503
rect 25869 77503 25927 77509
rect 25869 77500 25881 77503
rect 24699 77472 25881 77500
rect 24699 77469 24711 77472
rect 24653 77463 24711 77469
rect 25869 77469 25881 77472
rect 25915 77469 25927 77503
rect 25869 77463 25927 77469
rect 54481 77503 54539 77509
rect 54481 77469 54493 77503
rect 54527 77500 54539 77503
rect 55030 77500 55036 77512
rect 54527 77472 55036 77500
rect 54527 77469 54539 77472
rect 54481 77463 54539 77469
rect 55030 77460 55036 77472
rect 55088 77460 55094 77512
rect 15778 77404 16160 77432
rect 14642 77324 14648 77376
rect 14700 77324 14706 77376
rect 16132 77364 16160 77404
rect 16206 77392 16212 77444
rect 16264 77392 16270 77444
rect 55122 77432 55128 77444
rect 55083 77404 55128 77432
rect 55122 77392 55128 77404
rect 55180 77432 55186 77444
rect 55309 77435 55367 77441
rect 55309 77432 55321 77435
rect 55180 77404 55321 77432
rect 55180 77392 55186 77404
rect 55309 77401 55321 77404
rect 55355 77401 55367 77435
rect 55309 77395 55367 77401
rect 20714 77364 20720 77376
rect 16132 77336 20720 77364
rect 20714 77324 20720 77336
rect 20772 77324 20778 77376
rect 23474 77324 23480 77376
rect 23532 77324 23538 77376
rect 55030 77324 55036 77376
rect 55088 77364 55094 77376
rect 56597 77367 56655 77373
rect 56597 77364 56609 77367
rect 55088 77336 56609 77364
rect 55088 77324 55094 77336
rect 56597 77333 56609 77336
rect 56643 77364 56655 77367
rect 57149 77367 57207 77373
rect 57149 77364 57161 77367
rect 56643 77336 57161 77364
rect 56643 77333 56655 77336
rect 56597 77327 56655 77333
rect 57149 77333 57161 77336
rect 57195 77364 57207 77367
rect 59262 77364 59268 77376
rect 57195 77336 59268 77364
rect 57195 77333 57207 77336
rect 57149 77327 57207 77333
rect 59262 77324 59268 77336
rect 59320 77324 59326 77376
rect 82814 77324 82820 77376
rect 82872 77364 82878 77376
rect 83384 77373 83412 77540
rect 83737 77537 83749 77540
rect 83783 77568 83795 77571
rect 85945 77571 86003 77577
rect 85945 77568 85957 77571
rect 83783 77540 85957 77568
rect 83783 77537 83795 77540
rect 83737 77531 83795 77537
rect 85945 77537 85957 77540
rect 85991 77568 86003 77571
rect 86402 77568 86408 77580
rect 85991 77540 86408 77568
rect 85991 77537 86003 77540
rect 85945 77531 86003 77537
rect 86402 77528 86408 77540
rect 86460 77528 86466 77580
rect 86604 77577 86632 77608
rect 87230 77596 87236 77608
rect 87288 77596 87294 77648
rect 89441 77639 89499 77645
rect 89441 77605 89453 77639
rect 89487 77636 89499 77639
rect 89622 77636 89628 77648
rect 89487 77608 89628 77636
rect 89487 77605 89499 77608
rect 89441 77599 89499 77605
rect 89622 77596 89628 77608
rect 89680 77636 89686 77648
rect 89714 77636 89720 77648
rect 89680 77608 89720 77636
rect 89680 77596 89686 77608
rect 89714 77596 89720 77608
rect 89772 77596 89778 77648
rect 89806 77596 89812 77648
rect 89864 77636 89870 77648
rect 90453 77639 90511 77645
rect 89864 77608 90036 77636
rect 89864 77596 89870 77608
rect 86589 77571 86647 77577
rect 86589 77537 86601 77571
rect 86635 77537 86647 77571
rect 89898 77568 89904 77580
rect 86589 77531 86647 77537
rect 86696 77540 89904 77568
rect 83921 77503 83979 77509
rect 83921 77469 83933 77503
rect 83967 77500 83979 77503
rect 84565 77503 84623 77509
rect 84565 77500 84577 77503
rect 83967 77472 84577 77500
rect 83967 77469 83979 77472
rect 83921 77463 83979 77469
rect 84565 77469 84577 77472
rect 84611 77500 84623 77503
rect 86696 77500 86724 77540
rect 89898 77528 89904 77540
rect 89956 77528 89962 77580
rect 90008 77509 90036 77608
rect 90453 77605 90465 77639
rect 90499 77636 90511 77639
rect 90542 77636 90548 77648
rect 90499 77608 90548 77636
rect 90499 77605 90511 77608
rect 90453 77599 90511 77605
rect 90542 77596 90548 77608
rect 90600 77636 90606 77648
rect 91097 77639 91155 77645
rect 90600 77608 90680 77636
rect 90600 77596 90606 77608
rect 90652 77577 90680 77608
rect 91097 77605 91109 77639
rect 91143 77636 91155 77639
rect 91922 77636 91928 77648
rect 91143 77608 91928 77636
rect 91143 77605 91155 77608
rect 91097 77599 91155 77605
rect 91922 77596 91928 77608
rect 91980 77596 91986 77648
rect 94133 77639 94191 77645
rect 94133 77605 94145 77639
rect 94179 77636 94191 77639
rect 96522 77636 96528 77648
rect 94179 77608 96528 77636
rect 94179 77605 94191 77608
rect 94133 77599 94191 77605
rect 96522 77596 96528 77608
rect 96580 77596 96586 77648
rect 98917 77639 98975 77645
rect 98917 77605 98929 77639
rect 98963 77636 98975 77639
rect 108206 77636 108212 77648
rect 98963 77608 108212 77636
rect 98963 77605 98975 77608
rect 98917 77599 98975 77605
rect 108206 77596 108212 77608
rect 108264 77596 108270 77648
rect 90637 77571 90695 77577
rect 90637 77537 90649 77571
rect 90683 77537 90695 77571
rect 94593 77571 94651 77577
rect 94593 77568 94605 77571
rect 90637 77531 90695 77537
rect 93780 77540 94605 77568
rect 89993 77503 90051 77509
rect 84611 77472 86724 77500
rect 87064 77472 89944 77500
rect 84611 77469 84623 77472
rect 84565 77463 84623 77469
rect 83369 77367 83427 77373
rect 83369 77364 83381 77367
rect 82872 77336 83381 77364
rect 82872 77324 82878 77336
rect 83369 77333 83381 77336
rect 83415 77333 83427 77367
rect 83369 77327 83427 77333
rect 84010 77324 84016 77376
rect 84068 77324 84074 77376
rect 84381 77367 84439 77373
rect 84381 77333 84393 77367
rect 84427 77364 84439 77367
rect 85850 77364 85856 77376
rect 84427 77336 85856 77364
rect 84427 77333 84439 77336
rect 84381 77327 84439 77333
rect 85850 77324 85856 77336
rect 85908 77324 85914 77376
rect 86681 77367 86739 77373
rect 86681 77333 86693 77367
rect 86727 77364 86739 77367
rect 86770 77364 86776 77376
rect 86727 77336 86776 77364
rect 86727 77333 86739 77336
rect 86681 77327 86739 77333
rect 86770 77324 86776 77336
rect 86828 77324 86834 77376
rect 87064 77373 87092 77472
rect 89533 77435 89591 77441
rect 89533 77401 89545 77435
rect 89579 77401 89591 77435
rect 89533 77395 89591 77401
rect 87049 77367 87107 77373
rect 87049 77333 87061 77367
rect 87095 77333 87107 77367
rect 89548 77364 89576 77395
rect 89622 77392 89628 77444
rect 89680 77432 89686 77444
rect 89717 77435 89775 77441
rect 89717 77432 89729 77435
rect 89680 77404 89729 77432
rect 89680 77392 89686 77404
rect 89717 77401 89729 77404
rect 89763 77401 89775 77435
rect 89916 77432 89944 77472
rect 89993 77469 90005 77503
rect 90039 77469 90051 77503
rect 92474 77500 92480 77512
rect 89993 77463 90051 77469
rect 90100 77472 92480 77500
rect 90100 77432 90128 77472
rect 92474 77460 92480 77472
rect 92532 77460 92538 77512
rect 93780 77509 93808 77540
rect 94593 77537 94605 77540
rect 94639 77568 94651 77571
rect 105078 77568 105084 77580
rect 94639 77540 105084 77568
rect 94639 77537 94651 77540
rect 94593 77531 94651 77537
rect 105078 77528 105084 77540
rect 105136 77528 105142 77580
rect 93765 77503 93823 77509
rect 93765 77469 93777 77503
rect 93811 77469 93823 77503
rect 93765 77463 93823 77469
rect 93946 77460 93952 77512
rect 94004 77500 94010 77512
rect 94041 77503 94099 77509
rect 94041 77500 94053 77503
rect 94004 77472 94053 77500
rect 94004 77460 94010 77472
rect 94041 77469 94053 77472
rect 94087 77469 94099 77503
rect 94041 77463 94099 77469
rect 94866 77460 94872 77512
rect 94924 77500 94930 77512
rect 95145 77503 95203 77509
rect 95145 77500 95157 77503
rect 94924 77472 95157 77500
rect 94924 77460 94930 77472
rect 95145 77469 95157 77472
rect 95191 77469 95203 77503
rect 95145 77463 95203 77469
rect 96890 77460 96896 77512
rect 96948 77500 96954 77512
rect 97169 77503 97227 77509
rect 97169 77500 97181 77503
rect 96948 77472 97181 77500
rect 96948 77460 96954 77472
rect 97169 77469 97181 77472
rect 97215 77469 97227 77503
rect 97169 77463 97227 77469
rect 89916 77404 90128 77432
rect 89717 77395 89775 77401
rect 91462 77392 91468 77444
rect 91520 77432 91526 77444
rect 92014 77432 92020 77444
rect 91520 77404 92020 77432
rect 91520 77392 91526 77404
rect 92014 77392 92020 77404
rect 92072 77392 92078 77444
rect 94685 77435 94743 77441
rect 94685 77432 94697 77435
rect 92584 77404 94697 77432
rect 92584 77376 92612 77404
rect 94685 77401 94697 77404
rect 94731 77401 94743 77435
rect 94685 77395 94743 77401
rect 95234 77392 95240 77444
rect 95292 77432 95298 77444
rect 97445 77435 97503 77441
rect 97445 77432 97457 77435
rect 95292 77404 97457 77432
rect 95292 77392 95298 77404
rect 97445 77401 97457 77404
rect 97491 77401 97503 77435
rect 97445 77395 97503 77401
rect 97902 77392 97908 77444
rect 97960 77392 97966 77444
rect 89806 77364 89812 77376
rect 89548 77336 89812 77364
rect 87049 77327 87107 77333
rect 89806 77324 89812 77336
rect 89864 77324 89870 77376
rect 89901 77367 89959 77373
rect 89901 77333 89913 77367
rect 89947 77364 89959 77367
rect 90082 77364 90088 77376
rect 89947 77336 90088 77364
rect 89947 77333 89959 77336
rect 89901 77327 89959 77333
rect 90082 77324 90088 77336
rect 90140 77324 90146 77376
rect 91554 77324 91560 77376
rect 91612 77324 91618 77376
rect 91833 77367 91891 77373
rect 91833 77333 91845 77367
rect 91879 77364 91891 77367
rect 92198 77364 92204 77376
rect 91879 77336 92204 77364
rect 91879 77333 91891 77336
rect 91833 77327 91891 77333
rect 92198 77324 92204 77336
rect 92256 77324 92262 77376
rect 92477 77367 92535 77373
rect 92477 77333 92489 77367
rect 92523 77364 92535 77367
rect 92566 77364 92572 77376
rect 92523 77336 92572 77364
rect 92523 77333 92535 77336
rect 92477 77327 92535 77333
rect 92566 77324 92572 77336
rect 92624 77324 92630 77376
rect 93946 77324 93952 77376
rect 94004 77364 94010 77376
rect 94317 77367 94375 77373
rect 94317 77364 94329 77367
rect 94004 77336 94329 77364
rect 94004 77324 94010 77336
rect 94317 77333 94329 77336
rect 94363 77333 94375 77367
rect 94317 77327 94375 77333
rect 97626 77324 97632 77376
rect 97684 77364 97690 77376
rect 99098 77364 99104 77376
rect 97684 77336 99104 77364
rect 97684 77324 97690 77336
rect 99098 77324 99104 77336
rect 99156 77324 99162 77376
rect 1104 77274 108836 77296
rect 1104 77222 4874 77274
rect 4926 77222 4938 77274
rect 4990 77222 5002 77274
rect 5054 77222 5066 77274
rect 5118 77222 5130 77274
rect 5182 77222 35594 77274
rect 35646 77222 35658 77274
rect 35710 77222 35722 77274
rect 35774 77222 35786 77274
rect 35838 77222 35850 77274
rect 35902 77222 66314 77274
rect 66366 77222 66378 77274
rect 66430 77222 66442 77274
rect 66494 77222 66506 77274
rect 66558 77222 66570 77274
rect 66622 77222 97034 77274
rect 97086 77222 97098 77274
rect 97150 77222 97162 77274
rect 97214 77222 97226 77274
rect 97278 77222 97290 77274
rect 97342 77222 106658 77274
rect 106710 77222 106722 77274
rect 106774 77222 106786 77274
rect 106838 77222 106850 77274
rect 106902 77222 106914 77274
rect 106966 77222 108836 77274
rect 1104 77200 108836 77222
rect 1581 77163 1639 77169
rect 1581 77129 1593 77163
rect 1627 77160 1639 77163
rect 1857 77163 1915 77169
rect 1857 77160 1869 77163
rect 1627 77132 1869 77160
rect 1627 77129 1639 77132
rect 1581 77123 1639 77129
rect 1857 77129 1869 77132
rect 1903 77160 1915 77163
rect 2038 77160 2044 77172
rect 1903 77132 2044 77160
rect 1903 77129 1915 77132
rect 1857 77123 1915 77129
rect 2038 77120 2044 77132
rect 2096 77120 2102 77172
rect 8110 77120 8116 77172
rect 8168 77160 8174 77172
rect 46934 77160 46940 77172
rect 8168 77132 46940 77160
rect 8168 77120 8174 77132
rect 46934 77120 46940 77132
rect 46992 77120 46998 77172
rect 86402 77120 86408 77172
rect 86460 77160 86466 77172
rect 88521 77163 88579 77169
rect 88521 77160 88533 77163
rect 86460 77132 88533 77160
rect 86460 77120 86466 77132
rect 20714 77052 20720 77104
rect 20772 77092 20778 77104
rect 22373 77095 22431 77101
rect 22373 77092 22385 77095
rect 20772 77064 22385 77092
rect 20772 77052 20778 77064
rect 22373 77061 22385 77064
rect 22419 77061 22431 77095
rect 22373 77055 22431 77061
rect 24670 77052 24676 77104
rect 24728 77052 24734 77104
rect 25222 77052 25228 77104
rect 25280 77092 25286 77104
rect 25869 77095 25927 77101
rect 25869 77092 25881 77095
rect 25280 77064 25881 77092
rect 25280 77052 25286 77064
rect 25869 77061 25881 77064
rect 25915 77061 25927 77095
rect 25869 77055 25927 77061
rect 1210 76984 1216 77036
rect 1268 77024 1274 77036
rect 1489 77027 1547 77033
rect 1489 77024 1501 77027
rect 1268 76996 1501 77024
rect 1268 76984 1274 76996
rect 1489 76993 1501 76996
rect 1535 77024 1547 77027
rect 1949 77027 2007 77033
rect 1949 77024 1961 77027
rect 1535 76996 1961 77024
rect 1535 76993 1547 76996
rect 1489 76987 1547 76993
rect 1949 76993 1961 76996
rect 1995 76993 2007 77027
rect 1949 76987 2007 76993
rect 22462 76984 22468 77036
rect 22520 76984 22526 77036
rect 25777 77027 25835 77033
rect 23860 76996 25360 77024
rect 8202 76916 8208 76968
rect 8260 76956 8266 76968
rect 23860 76956 23888 76996
rect 8260 76928 23888 76956
rect 8260 76916 8266 76928
rect 9122 76848 9128 76900
rect 9180 76888 9186 76900
rect 25222 76888 25228 76900
rect 9180 76860 25228 76888
rect 9180 76848 9186 76860
rect 25222 76848 25228 76860
rect 25280 76848 25286 76900
rect 25332 76888 25360 76996
rect 25777 76993 25789 77027
rect 25823 77024 25835 77027
rect 32950 77024 32956 77036
rect 25823 76996 32956 77024
rect 25823 76993 25835 76996
rect 25777 76987 25835 76993
rect 32950 76984 32956 76996
rect 33008 76984 33014 77036
rect 26053 76959 26111 76965
rect 26053 76925 26065 76959
rect 26099 76956 26111 76959
rect 26326 76956 26332 76968
rect 26099 76928 26332 76956
rect 26099 76925 26111 76928
rect 26053 76919 26111 76925
rect 26326 76916 26332 76928
rect 26384 76916 26390 76968
rect 88352 76956 88380 77132
rect 88521 77129 88533 77132
rect 88567 77129 88579 77163
rect 88521 77123 88579 77129
rect 89533 77163 89591 77169
rect 89533 77129 89545 77163
rect 89579 77129 89591 77163
rect 89533 77123 89591 77129
rect 89073 77095 89131 77101
rect 89073 77061 89085 77095
rect 89119 77092 89131 77095
rect 89548 77092 89576 77123
rect 89714 77120 89720 77172
rect 89772 77160 89778 77172
rect 90177 77163 90235 77169
rect 90177 77160 90189 77163
rect 89772 77132 90189 77160
rect 89772 77120 89778 77132
rect 90177 77129 90189 77132
rect 90223 77160 90235 77163
rect 90358 77160 90364 77172
rect 90223 77132 90364 77160
rect 90223 77129 90235 77132
rect 90177 77123 90235 77129
rect 90358 77120 90364 77132
rect 90416 77120 90422 77172
rect 91741 77163 91799 77169
rect 91741 77129 91753 77163
rect 91787 77160 91799 77163
rect 95234 77160 95240 77172
rect 91787 77132 95240 77160
rect 91787 77129 91799 77132
rect 91741 77123 91799 77129
rect 95234 77120 95240 77132
rect 95292 77120 95298 77172
rect 96890 77160 96896 77172
rect 95804 77132 96896 77160
rect 89119 77064 89392 77092
rect 89548 77064 92888 77092
rect 89119 77061 89131 77064
rect 89073 77055 89131 77061
rect 88426 76984 88432 77036
rect 88484 77024 88490 77036
rect 89165 77027 89223 77033
rect 89165 77024 89177 77027
rect 88484 76996 89177 77024
rect 88484 76984 88490 76996
rect 89165 76993 89177 76996
rect 89211 76993 89223 77027
rect 89364 77024 89392 77064
rect 89717 77027 89775 77033
rect 89717 77024 89729 77027
rect 89364 76996 89729 77024
rect 89165 76987 89223 76993
rect 89717 76993 89729 76996
rect 89763 77024 89775 77027
rect 90266 77024 90272 77036
rect 89763 76996 90272 77024
rect 89763 76993 89775 76996
rect 89717 76987 89775 76993
rect 90266 76984 90272 76996
rect 90324 76984 90330 77036
rect 90358 76984 90364 77036
rect 90416 76984 90422 77036
rect 90542 76984 90548 77036
rect 90600 76984 90606 77036
rect 91373 77027 91431 77033
rect 91373 77024 91385 77027
rect 90652 76996 91385 77024
rect 88889 76959 88947 76965
rect 88889 76956 88901 76959
rect 88352 76928 88901 76956
rect 88889 76925 88901 76928
rect 88935 76925 88947 76959
rect 88889 76919 88947 76925
rect 41322 76888 41328 76900
rect 25332 76860 41328 76888
rect 41322 76848 41328 76860
rect 41380 76848 41386 76900
rect 88904 76888 88932 76919
rect 89254 76916 89260 76968
rect 89312 76956 89318 76968
rect 90652 76956 90680 76996
rect 91373 76993 91385 76996
rect 91419 76993 91431 77027
rect 91373 76987 91431 76993
rect 91922 76984 91928 77036
rect 91980 76984 91986 77036
rect 92106 76984 92112 77036
rect 92164 76984 92170 77036
rect 92661 77027 92719 77033
rect 92661 76993 92673 77027
rect 92707 76993 92719 77027
rect 92661 76987 92719 76993
rect 89312 76928 90680 76956
rect 91097 76959 91155 76965
rect 89312 76916 89318 76928
rect 91097 76925 91109 76959
rect 91143 76925 91155 76959
rect 91097 76919 91155 76925
rect 91281 76959 91339 76965
rect 91281 76925 91293 76959
rect 91327 76956 91339 76959
rect 92124 76956 92152 76984
rect 91327 76928 92152 76956
rect 91327 76925 91339 76928
rect 91281 76919 91339 76925
rect 90821 76891 90879 76897
rect 90821 76888 90833 76891
rect 88904 76860 90833 76888
rect 90821 76857 90833 76860
rect 90867 76888 90879 76891
rect 91112 76888 91140 76919
rect 90867 76860 91140 76888
rect 90867 76857 90879 76860
rect 90821 76851 90879 76857
rect 22370 76780 22376 76832
rect 22428 76820 22434 76832
rect 22557 76823 22615 76829
rect 22557 76820 22569 76823
rect 22428 76792 22569 76820
rect 22428 76780 22434 76792
rect 22557 76789 22569 76792
rect 22603 76789 22615 76823
rect 22557 76783 22615 76789
rect 25406 76780 25412 76832
rect 25464 76780 25470 76832
rect 26326 76780 26332 76832
rect 26384 76780 26390 76832
rect 55030 76780 55036 76832
rect 55088 76780 55094 76832
rect 90450 76780 90456 76832
rect 90508 76780 90514 76832
rect 92566 76780 92572 76832
rect 92624 76820 92630 76832
rect 92676 76820 92704 76987
rect 92860 76956 92888 77064
rect 93946 76984 93952 77036
rect 94004 77024 94010 77036
rect 95804 77033 95832 77132
rect 96890 77120 96896 77132
rect 96948 77160 96954 77172
rect 97626 77160 97632 77172
rect 96948 77132 97632 77160
rect 96948 77120 96954 77132
rect 97626 77120 97632 77132
rect 97684 77120 97690 77172
rect 96522 77052 96528 77104
rect 96580 77052 96586 77104
rect 98730 77052 98736 77104
rect 98788 77092 98794 77104
rect 99469 77095 99527 77101
rect 99469 77092 99481 77095
rect 98788 77064 99481 77092
rect 98788 77052 98794 77064
rect 99469 77061 99481 77064
rect 99515 77061 99527 77095
rect 99469 77055 99527 77061
rect 94225 77027 94283 77033
rect 94225 77024 94237 77027
rect 94004 76996 94237 77024
rect 94004 76984 94010 76996
rect 94225 76993 94237 76996
rect 94271 76993 94283 77027
rect 94225 76987 94283 76993
rect 95789 77027 95847 77033
rect 95789 76993 95801 77027
rect 95835 76993 95847 77027
rect 95789 76987 95847 76993
rect 99098 76984 99104 77036
rect 99156 76984 99162 77036
rect 99282 76984 99288 77036
rect 99340 76984 99346 77036
rect 99561 77027 99619 77033
rect 99561 76993 99573 77027
rect 99607 76993 99619 77027
rect 99561 76987 99619 76993
rect 96065 76959 96123 76965
rect 96065 76956 96077 76959
rect 92860 76928 96077 76956
rect 96065 76925 96077 76928
rect 96111 76925 96123 76959
rect 96065 76919 96123 76925
rect 99190 76916 99196 76968
rect 99248 76956 99254 76968
rect 99576 76956 99604 76987
rect 100110 76984 100116 77036
rect 100168 77024 100174 77036
rect 100481 77027 100539 77033
rect 100481 77024 100493 77027
rect 100168 76996 100493 77024
rect 100168 76984 100174 76996
rect 100481 76993 100493 76996
rect 100527 76993 100539 77027
rect 100481 76987 100539 76993
rect 100665 77027 100723 77033
rect 100665 76993 100677 77027
rect 100711 77024 100723 77027
rect 100754 77024 100760 77036
rect 100711 76996 100760 77024
rect 100711 76993 100723 76996
rect 100665 76987 100723 76993
rect 100754 76984 100760 76996
rect 100812 76984 100818 77036
rect 108209 77027 108267 77033
rect 108209 76993 108221 77027
rect 108255 76993 108267 77027
rect 108209 76987 108267 76993
rect 99248 76928 99604 76956
rect 99248 76916 99254 76928
rect 100570 76916 100576 76968
rect 100628 76956 100634 76968
rect 108224 76956 108252 76987
rect 100628 76928 108252 76956
rect 100628 76916 100634 76928
rect 97537 76891 97595 76897
rect 97537 76857 97549 76891
rect 97583 76888 97595 76891
rect 107654 76888 107660 76900
rect 97583 76860 107660 76888
rect 97583 76857 97595 76860
rect 97537 76851 97595 76857
rect 107654 76848 107660 76860
rect 107712 76848 107718 76900
rect 108390 76848 108396 76900
rect 108448 76848 108454 76900
rect 93121 76823 93179 76829
rect 93121 76820 93133 76823
rect 92624 76792 93133 76820
rect 92624 76780 92630 76792
rect 93121 76789 93133 76792
rect 93167 76789 93179 76823
rect 93121 76783 93179 76789
rect 94038 76780 94044 76832
rect 94096 76780 94102 76832
rect 98454 76780 98460 76832
rect 98512 76820 98518 76832
rect 99193 76823 99251 76829
rect 99193 76820 99205 76823
rect 98512 76792 99205 76820
rect 98512 76780 98518 76792
rect 99193 76789 99205 76792
rect 99239 76789 99251 76823
rect 99193 76783 99251 76789
rect 100481 76823 100539 76829
rect 100481 76789 100493 76823
rect 100527 76820 100539 76823
rect 101030 76820 101036 76832
rect 100527 76792 101036 76820
rect 100527 76789 100539 76792
rect 100481 76783 100539 76789
rect 101030 76780 101036 76792
rect 101088 76780 101094 76832
rect 1104 76730 108836 76752
rect 1104 76678 4214 76730
rect 4266 76678 4278 76730
rect 4330 76678 4342 76730
rect 4394 76678 4406 76730
rect 4458 76678 4470 76730
rect 4522 76678 34934 76730
rect 34986 76678 34998 76730
rect 35050 76678 35062 76730
rect 35114 76678 35126 76730
rect 35178 76678 35190 76730
rect 35242 76678 65654 76730
rect 65706 76678 65718 76730
rect 65770 76678 65782 76730
rect 65834 76678 65846 76730
rect 65898 76678 65910 76730
rect 65962 76678 96374 76730
rect 96426 76678 96438 76730
rect 96490 76678 96502 76730
rect 96554 76678 96566 76730
rect 96618 76678 96630 76730
rect 96682 76678 108836 76730
rect 1104 76656 108836 76678
rect 9398 76576 9404 76628
rect 9456 76616 9462 76628
rect 9456 76588 31754 76616
rect 9456 76576 9462 76588
rect 19334 76508 19340 76560
rect 19392 76548 19398 76560
rect 23201 76551 23259 76557
rect 23201 76548 23213 76551
rect 19392 76520 23213 76548
rect 19392 76508 19398 76520
rect 23201 76517 23213 76520
rect 23247 76517 23259 76551
rect 23201 76511 23259 76517
rect 13998 76440 14004 76492
rect 14056 76480 14062 76492
rect 23017 76483 23075 76489
rect 23017 76480 23029 76483
rect 14056 76452 23029 76480
rect 14056 76440 14062 76452
rect 23017 76449 23029 76452
rect 23063 76480 23075 76483
rect 23661 76483 23719 76489
rect 23661 76480 23673 76483
rect 23063 76452 23673 76480
rect 23063 76449 23075 76452
rect 23017 76443 23075 76449
rect 23661 76449 23673 76452
rect 23707 76449 23719 76483
rect 23661 76443 23719 76449
rect 23845 76483 23903 76489
rect 23845 76449 23857 76483
rect 23891 76480 23903 76483
rect 24121 76483 24179 76489
rect 24121 76480 24133 76483
rect 23891 76452 24133 76480
rect 23891 76449 23903 76452
rect 23845 76443 23903 76449
rect 24121 76449 24133 76452
rect 24167 76480 24179 76483
rect 26326 76480 26332 76492
rect 24167 76452 26332 76480
rect 24167 76449 24179 76452
rect 24121 76443 24179 76449
rect 26326 76440 26332 76452
rect 26384 76480 26390 76492
rect 27341 76483 27399 76489
rect 27341 76480 27353 76483
rect 26384 76452 27353 76480
rect 26384 76440 26390 76452
rect 27341 76449 27353 76452
rect 27387 76449 27399 76483
rect 27341 76443 27399 76449
rect 1673 76415 1731 76421
rect 1673 76381 1685 76415
rect 1719 76412 1731 76415
rect 14550 76412 14556 76424
rect 1719 76384 14556 76412
rect 1719 76381 1731 76384
rect 1673 76375 1731 76381
rect 14550 76372 14556 76384
rect 14608 76372 14614 76424
rect 17126 76372 17132 76424
rect 17184 76412 17190 76424
rect 26513 76415 26571 76421
rect 26513 76412 26525 76415
rect 17184 76384 26525 76412
rect 17184 76372 17190 76384
rect 26513 76381 26525 76384
rect 26559 76412 26571 76415
rect 27157 76415 27215 76421
rect 27157 76412 27169 76415
rect 26559 76384 27169 76412
rect 26559 76381 26571 76384
rect 26513 76375 26571 76381
rect 27157 76381 27169 76384
rect 27203 76381 27215 76415
rect 27356 76412 27384 76443
rect 27522 76440 27528 76492
rect 27580 76480 27586 76492
rect 28997 76483 29055 76489
rect 28997 76480 29009 76483
rect 27580 76452 29009 76480
rect 27580 76440 27586 76452
rect 28997 76449 29009 76452
rect 29043 76449 29055 76483
rect 28997 76443 29055 76449
rect 29089 76483 29147 76489
rect 29089 76449 29101 76483
rect 29135 76449 29147 76483
rect 29089 76443 29147 76449
rect 27617 76415 27675 76421
rect 27617 76412 27629 76415
rect 27356 76384 27629 76412
rect 27157 76375 27215 76381
rect 27617 76381 27629 76384
rect 27663 76412 27675 76415
rect 29104 76412 29132 76443
rect 27663 76384 29132 76412
rect 31726 76412 31754 76588
rect 41322 76576 41328 76628
rect 41380 76576 41386 76628
rect 46934 76576 46940 76628
rect 46992 76576 46998 76628
rect 58618 76576 58624 76628
rect 58676 76616 58682 76628
rect 59262 76616 59268 76628
rect 58676 76588 59268 76616
rect 58676 76576 58682 76588
rect 59262 76576 59268 76588
rect 59320 76616 59326 76628
rect 60461 76619 60519 76625
rect 60461 76616 60473 76619
rect 59320 76588 60473 76616
rect 59320 76576 59326 76588
rect 60461 76585 60473 76588
rect 60507 76585 60519 76619
rect 60461 76579 60519 76585
rect 66993 76619 67051 76625
rect 66993 76585 67005 76619
rect 67039 76616 67051 76619
rect 68922 76616 68928 76628
rect 67039 76588 68928 76616
rect 67039 76585 67051 76588
rect 66993 76579 67051 76585
rect 60476 76480 60504 76579
rect 68922 76576 68928 76588
rect 68980 76576 68986 76628
rect 92474 76576 92480 76628
rect 92532 76616 92538 76628
rect 94501 76619 94559 76625
rect 92532 76588 94084 76616
rect 92532 76576 92538 76588
rect 94056 76548 94084 76588
rect 94501 76585 94513 76619
rect 94547 76616 94559 76619
rect 97994 76616 98000 76628
rect 94547 76588 98000 76616
rect 94547 76585 94559 76588
rect 94501 76579 94559 76585
rect 97994 76576 98000 76588
rect 98052 76576 98058 76628
rect 99098 76576 99104 76628
rect 99156 76616 99162 76628
rect 99156 76588 99880 76616
rect 99156 76576 99162 76588
rect 95418 76548 95424 76560
rect 94056 76520 95424 76548
rect 95418 76508 95424 76520
rect 95476 76508 95482 76560
rect 99282 76508 99288 76560
rect 99340 76548 99346 76560
rect 99340 76520 99696 76548
rect 99340 76508 99346 76520
rect 60737 76483 60795 76489
rect 60737 76480 60749 76483
rect 60476 76452 60749 76480
rect 60737 76449 60749 76452
rect 60783 76449 60795 76483
rect 60737 76443 60795 76449
rect 82538 76440 82544 76492
rect 82596 76480 82602 76492
rect 82722 76480 82728 76492
rect 82596 76452 82728 76480
rect 82596 76440 82602 76452
rect 82722 76440 82728 76452
rect 82780 76480 82786 76492
rect 82817 76483 82875 76489
rect 82817 76480 82829 76483
rect 82780 76452 82829 76480
rect 82780 76440 82786 76452
rect 82817 76449 82829 76452
rect 82863 76449 82875 76483
rect 82817 76443 82875 76449
rect 85850 76440 85856 76492
rect 85908 76480 85914 76492
rect 93029 76483 93087 76489
rect 93029 76480 93041 76483
rect 85908 76452 93041 76480
rect 85908 76440 85914 76452
rect 93029 76449 93041 76452
rect 93075 76449 93087 76483
rect 93029 76443 93087 76449
rect 98089 76483 98147 76489
rect 98089 76449 98101 76483
rect 98135 76480 98147 76483
rect 98270 76480 98276 76492
rect 98135 76452 98276 76480
rect 98135 76449 98147 76452
rect 98089 76443 98147 76449
rect 98270 76440 98276 76452
rect 98328 76480 98334 76492
rect 98328 76452 99420 76480
rect 98328 76440 98334 76452
rect 41233 76415 41291 76421
rect 31726 76384 41092 76412
rect 27663 76381 27675 76384
rect 27617 76375 27675 76381
rect 842 76236 848 76288
rect 900 76276 906 76288
rect 1489 76279 1547 76285
rect 1489 76276 1501 76279
rect 900 76248 1501 76276
rect 900 76236 906 76248
rect 1489 76245 1501 76248
rect 1535 76245 1547 76279
rect 1489 76239 1547 76245
rect 23566 76236 23572 76288
rect 23624 76236 23630 76288
rect 24854 76236 24860 76288
rect 24912 76276 24918 76288
rect 26697 76279 26755 76285
rect 26697 76276 26709 76279
rect 24912 76248 26709 76276
rect 24912 76236 24918 76248
rect 26697 76245 26709 76248
rect 26743 76245 26755 76279
rect 26697 76239 26755 76245
rect 27065 76279 27123 76285
rect 27065 76245 27077 76279
rect 27111 76276 27123 76279
rect 28442 76276 28448 76288
rect 27111 76248 28448 76276
rect 27111 76245 27123 76248
rect 27065 76239 27123 76245
rect 28442 76236 28448 76248
rect 28500 76236 28506 76288
rect 28534 76236 28540 76288
rect 28592 76236 28598 76288
rect 28828 76276 28856 76384
rect 28905 76347 28963 76353
rect 28905 76313 28917 76347
rect 28951 76344 28963 76347
rect 30282 76344 30288 76356
rect 28951 76316 30288 76344
rect 28951 76313 28963 76316
rect 28905 76307 28963 76313
rect 30282 76304 30288 76316
rect 30340 76304 30346 76356
rect 40966 76347 41024 76353
rect 40966 76313 40978 76347
rect 41012 76313 41024 76347
rect 41064 76344 41092 76384
rect 41233 76381 41245 76415
rect 41279 76412 41291 76415
rect 41601 76415 41659 76421
rect 41601 76412 41613 76415
rect 41279 76384 41613 76412
rect 41279 76381 41291 76384
rect 41233 76375 41291 76381
rect 41601 76381 41613 76384
rect 41647 76412 41659 76415
rect 44269 76415 44327 76421
rect 44269 76412 44281 76415
rect 41647 76384 44281 76412
rect 41647 76381 41659 76384
rect 41601 76375 41659 76381
rect 44269 76381 44281 76384
rect 44315 76412 44327 76415
rect 44637 76415 44695 76421
rect 44637 76412 44649 76415
rect 44315 76384 44649 76412
rect 44315 76381 44327 76384
rect 44269 76375 44327 76381
rect 44637 76381 44649 76384
rect 44683 76412 44695 76415
rect 46845 76415 46903 76421
rect 46845 76412 46857 76415
rect 44683 76384 46857 76412
rect 44683 76381 44695 76384
rect 44637 76375 44695 76381
rect 46845 76381 46857 76384
rect 46891 76412 46903 76415
rect 47121 76415 47179 76421
rect 47121 76412 47133 76415
rect 46891 76384 47133 76412
rect 46891 76381 46903 76384
rect 46845 76375 46903 76381
rect 47121 76381 47133 76384
rect 47167 76412 47179 76415
rect 55030 76412 55036 76424
rect 47167 76384 55036 76412
rect 47167 76381 47179 76384
rect 47121 76375 47179 76381
rect 55030 76372 55036 76384
rect 55088 76372 55094 76424
rect 62853 76415 62911 76421
rect 62853 76381 62865 76415
rect 62899 76412 62911 76415
rect 64325 76415 64383 76421
rect 64325 76412 64337 76415
rect 62899 76384 64337 76412
rect 62899 76381 62911 76384
rect 62853 76375 62911 76381
rect 64325 76381 64337 76384
rect 64371 76412 64383 76415
rect 65613 76415 65671 76421
rect 65613 76412 65625 76415
rect 64371 76384 65625 76412
rect 64371 76381 64383 76384
rect 64325 76375 64383 76381
rect 65613 76381 65625 76384
rect 65659 76412 65671 76415
rect 67177 76415 67235 76421
rect 67177 76412 67189 76415
rect 65659 76384 67189 76412
rect 65659 76381 65671 76384
rect 65613 76375 65671 76381
rect 67177 76381 67189 76384
rect 67223 76412 67235 76415
rect 67637 76415 67695 76421
rect 67637 76412 67649 76415
rect 67223 76384 67649 76412
rect 67223 76381 67235 76384
rect 67177 76375 67235 76381
rect 67637 76381 67649 76384
rect 67683 76412 67695 76415
rect 85117 76415 85175 76421
rect 67683 76384 69152 76412
rect 67683 76381 67695 76384
rect 67637 76375 67695 76381
rect 69124 76356 69152 76384
rect 85117 76381 85129 76415
rect 85163 76412 85175 76415
rect 85209 76415 85267 76421
rect 85209 76412 85221 76415
rect 85163 76384 85221 76412
rect 85163 76381 85175 76384
rect 85117 76375 85175 76381
rect 85209 76381 85221 76384
rect 85255 76412 85267 76415
rect 86862 76412 86868 76424
rect 85255 76384 86868 76412
rect 85255 76381 85267 76384
rect 85209 76375 85267 76381
rect 86862 76372 86868 76384
rect 86920 76372 86926 76424
rect 92753 76415 92811 76421
rect 92753 76412 92765 76415
rect 92584 76384 92765 76412
rect 44002 76347 44060 76353
rect 44002 76344 44014 76347
rect 41064 76316 44014 76344
rect 40966 76307 41024 76313
rect 44002 76313 44014 76316
rect 44048 76344 44060 76347
rect 44361 76347 44419 76353
rect 44361 76344 44373 76347
rect 44048 76316 44373 76344
rect 44048 76313 44060 76316
rect 44002 76307 44060 76313
rect 44361 76313 44373 76316
rect 44407 76313 44419 76347
rect 44361 76307 44419 76313
rect 46600 76347 46658 76353
rect 46600 76313 46612 76347
rect 46646 76344 46658 76347
rect 46934 76344 46940 76356
rect 46646 76316 46940 76344
rect 46646 76313 46658 76316
rect 46600 76307 46658 76313
rect 29641 76279 29699 76285
rect 29641 76276 29653 76279
rect 28828 76248 29653 76276
rect 29641 76245 29653 76248
rect 29687 76276 29699 76279
rect 33042 76276 33048 76288
rect 29687 76248 33048 76276
rect 29687 76245 29699 76248
rect 29641 76239 29699 76245
rect 33042 76236 33048 76248
rect 33100 76236 33106 76288
rect 39850 76236 39856 76288
rect 39908 76236 39914 76288
rect 40972 76276 41000 76307
rect 46934 76304 46940 76316
rect 46992 76304 46998 76356
rect 61010 76353 61016 76356
rect 60277 76347 60335 76353
rect 60277 76313 60289 76347
rect 60323 76344 60335 76347
rect 61004 76344 61016 76353
rect 60323 76316 61016 76344
rect 60323 76313 60335 76316
rect 60277 76307 60335 76313
rect 61004 76307 61016 76316
rect 61010 76304 61016 76307
rect 61068 76304 61074 76356
rect 63126 76353 63132 76356
rect 62761 76347 62819 76353
rect 62761 76313 62773 76347
rect 62807 76344 62819 76347
rect 63120 76344 63132 76353
rect 62807 76316 63132 76344
rect 62807 76313 62819 76316
rect 62761 76307 62819 76313
rect 63120 76307 63132 76316
rect 63126 76304 63132 76307
rect 63184 76304 63190 76356
rect 65429 76347 65487 76353
rect 65429 76313 65441 76347
rect 65475 76344 65487 76347
rect 65880 76347 65938 76353
rect 65880 76344 65892 76347
rect 65475 76316 65892 76344
rect 65475 76313 65487 76316
rect 65429 76307 65487 76313
rect 65880 76313 65892 76316
rect 65926 76344 65938 76347
rect 65978 76344 65984 76356
rect 65926 76316 65984 76344
rect 65926 76313 65938 76316
rect 65880 76307 65938 76313
rect 65978 76304 65984 76316
rect 66036 76304 66042 76356
rect 67910 76353 67916 76356
rect 67545 76347 67603 76353
rect 67545 76313 67557 76347
rect 67591 76344 67603 76347
rect 67904 76344 67916 76353
rect 67591 76316 67916 76344
rect 67591 76313 67603 76316
rect 67545 76307 67603 76313
rect 67904 76307 67916 76316
rect 67910 76304 67916 76307
rect 67968 76304 67974 76356
rect 69106 76304 69112 76356
rect 69164 76304 69170 76356
rect 83001 76347 83059 76353
rect 83001 76313 83013 76347
rect 83047 76344 83059 76347
rect 83047 76316 83780 76344
rect 83047 76313 83059 76316
rect 83001 76307 83059 76313
rect 41322 76276 41328 76288
rect 40972 76248 41328 76276
rect 41322 76236 41328 76248
rect 41380 76236 41386 76288
rect 42886 76236 42892 76288
rect 42944 76236 42950 76288
rect 45462 76236 45468 76288
rect 45520 76236 45526 76288
rect 62114 76236 62120 76288
rect 62172 76236 62178 76288
rect 64230 76236 64236 76288
rect 64288 76236 64294 76288
rect 69017 76279 69075 76285
rect 69017 76245 69029 76279
rect 69063 76276 69075 76279
rect 74534 76276 74540 76288
rect 69063 76248 74540 76276
rect 69063 76245 69075 76248
rect 69017 76239 69075 76245
rect 74534 76236 74540 76248
rect 74592 76236 74598 76288
rect 82538 76236 82544 76288
rect 82596 76236 82602 76288
rect 83090 76236 83096 76288
rect 83148 76236 83154 76288
rect 83458 76236 83464 76288
rect 83516 76236 83522 76288
rect 83642 76236 83648 76288
rect 83700 76236 83706 76288
rect 83752 76285 83780 76316
rect 84838 76304 84844 76356
rect 84896 76353 84902 76356
rect 84896 76344 84908 76353
rect 84896 76316 84941 76344
rect 84896 76307 84908 76316
rect 84896 76304 84902 76307
rect 92584 76288 92612 76384
rect 92753 76381 92765 76384
rect 92799 76381 92811 76415
rect 92753 76375 92811 76381
rect 98454 76372 98460 76424
rect 98512 76372 98518 76424
rect 98638 76372 98644 76424
rect 98696 76372 98702 76424
rect 99006 76372 99012 76424
rect 99064 76372 99070 76424
rect 93486 76304 93492 76356
rect 93544 76304 93550 76356
rect 97718 76304 97724 76356
rect 97776 76344 97782 76356
rect 97813 76347 97871 76353
rect 97813 76344 97825 76347
rect 97776 76316 97825 76344
rect 97776 76304 97782 76316
rect 97813 76313 97825 76316
rect 97859 76313 97871 76347
rect 97813 76307 97871 76313
rect 98178 76304 98184 76356
rect 98236 76344 98242 76356
rect 99190 76344 99196 76356
rect 98236 76316 99196 76344
rect 98236 76304 98242 76316
rect 99190 76304 99196 76316
rect 99248 76344 99254 76356
rect 99392 76353 99420 76452
rect 99668 76421 99696 76520
rect 99852 76421 99880 76588
rect 100573 76483 100631 76489
rect 100573 76449 100585 76483
rect 100619 76480 100631 76483
rect 100938 76480 100944 76492
rect 100619 76452 100944 76480
rect 100619 76449 100631 76452
rect 100573 76443 100631 76449
rect 100938 76440 100944 76452
rect 100996 76440 101002 76492
rect 101030 76440 101036 76492
rect 101088 76440 101094 76492
rect 99653 76415 99711 76421
rect 99653 76381 99665 76415
rect 99699 76381 99711 76415
rect 99653 76375 99711 76381
rect 99837 76415 99895 76421
rect 99837 76381 99849 76415
rect 99883 76412 99895 76415
rect 100386 76412 100392 76424
rect 99883 76384 100392 76412
rect 99883 76381 99895 76384
rect 99837 76375 99895 76381
rect 100386 76372 100392 76384
rect 100444 76372 100450 76424
rect 101122 76372 101128 76424
rect 101180 76372 101186 76424
rect 108209 76415 108267 76421
rect 108209 76412 108221 76415
rect 108040 76384 108221 76412
rect 99285 76347 99343 76353
rect 99285 76344 99297 76347
rect 99248 76316 99297 76344
rect 99248 76304 99254 76316
rect 99285 76313 99297 76316
rect 99331 76313 99343 76347
rect 99285 76307 99343 76313
rect 99377 76347 99435 76353
rect 99377 76313 99389 76347
rect 99423 76344 99435 76347
rect 99558 76344 99564 76356
rect 99423 76316 99564 76344
rect 99423 76313 99435 76316
rect 99377 76307 99435 76313
rect 83737 76279 83795 76285
rect 83737 76245 83749 76279
rect 83783 76245 83795 76279
rect 83737 76239 83795 76245
rect 92566 76236 92572 76288
rect 92624 76236 92630 76288
rect 99300 76276 99328 76307
rect 99558 76304 99564 76316
rect 99616 76304 99622 76356
rect 100297 76347 100355 76353
rect 100297 76313 100309 76347
rect 100343 76344 100355 76347
rect 100343 76316 100800 76344
rect 100343 76313 100355 76316
rect 100297 76307 100355 76313
rect 99929 76279 99987 76285
rect 99929 76276 99941 76279
rect 99300 76248 99941 76276
rect 99929 76245 99941 76248
rect 99975 76245 99987 76279
rect 99929 76239 99987 76245
rect 100018 76236 100024 76288
rect 100076 76276 100082 76288
rect 100772 76285 100800 76316
rect 100389 76279 100447 76285
rect 100389 76276 100401 76279
rect 100076 76248 100401 76276
rect 100076 76236 100082 76248
rect 100389 76245 100401 76248
rect 100435 76245 100447 76279
rect 100389 76239 100447 76245
rect 100757 76279 100815 76285
rect 100757 76245 100769 76279
rect 100803 76245 100815 76279
rect 100757 76239 100815 76245
rect 107930 76236 107936 76288
rect 107988 76276 107994 76288
rect 108040 76285 108068 76384
rect 108209 76381 108221 76384
rect 108255 76381 108267 76415
rect 108209 76375 108267 76381
rect 108025 76279 108083 76285
rect 108025 76276 108037 76279
rect 107988 76248 108037 76276
rect 107988 76236 107994 76248
rect 108025 76245 108037 76248
rect 108071 76245 108083 76279
rect 108025 76239 108083 76245
rect 108390 76236 108396 76288
rect 108448 76236 108454 76288
rect 1104 76186 108836 76208
rect 1104 76134 4874 76186
rect 4926 76134 4938 76186
rect 4990 76134 5002 76186
rect 5054 76134 5066 76186
rect 5118 76134 5130 76186
rect 5182 76134 35594 76186
rect 35646 76134 35658 76186
rect 35710 76134 35722 76186
rect 35774 76134 35786 76186
rect 35838 76134 35850 76186
rect 35902 76134 66314 76186
rect 66366 76134 66378 76186
rect 66430 76134 66442 76186
rect 66494 76134 66506 76186
rect 66558 76134 66570 76186
rect 66622 76134 97034 76186
rect 97086 76134 97098 76186
rect 97150 76134 97162 76186
rect 97214 76134 97226 76186
rect 97278 76134 97290 76186
rect 97342 76134 108836 76186
rect 1104 76112 108836 76134
rect 14642 76032 14648 76084
rect 14700 76072 14706 76084
rect 14700 76044 16528 76072
rect 14700 76032 14706 76044
rect 16298 76004 16304 76016
rect 15778 75976 16304 76004
rect 16298 75964 16304 75976
rect 16356 75964 16362 76016
rect 1673 75939 1731 75945
rect 1673 75905 1685 75939
rect 1719 75936 1731 75939
rect 11054 75936 11060 75948
rect 1719 75908 11060 75936
rect 1719 75905 1731 75908
rect 1673 75899 1731 75905
rect 11054 75896 11060 75908
rect 11112 75896 11118 75948
rect 14550 75896 14556 75948
rect 14608 75936 14614 75948
rect 16500 75945 16528 76044
rect 16574 76032 16580 76084
rect 16632 76072 16638 76084
rect 22278 76072 22284 76084
rect 16632 76044 22284 76072
rect 16632 76032 16638 76044
rect 22278 76032 22284 76044
rect 22336 76032 22342 76084
rect 23566 76032 23572 76084
rect 23624 76072 23630 76084
rect 30558 76072 30564 76084
rect 23624 76044 30564 76072
rect 23624 76032 23630 76044
rect 30558 76032 30564 76044
rect 30616 76032 30622 76084
rect 62114 76032 62120 76084
rect 62172 76072 62178 76084
rect 68462 76072 68468 76084
rect 62172 76044 68468 76072
rect 62172 76032 62178 76044
rect 68462 76032 68468 76044
rect 68520 76032 68526 76084
rect 83642 76032 83648 76084
rect 83700 76072 83706 76084
rect 83737 76075 83795 76081
rect 83737 76072 83749 76075
rect 83700 76044 83749 76072
rect 83700 76032 83706 76044
rect 83737 76041 83749 76044
rect 83783 76072 83795 76075
rect 84838 76072 84844 76084
rect 83783 76044 84844 76072
rect 83783 76041 83795 76044
rect 83737 76035 83795 76041
rect 84838 76032 84844 76044
rect 84896 76032 84902 76084
rect 90069 76075 90127 76081
rect 90069 76041 90081 76075
rect 90115 76072 90127 76075
rect 90450 76072 90456 76084
rect 90115 76044 90456 76072
rect 90115 76041 90127 76044
rect 90069 76035 90127 76041
rect 90450 76032 90456 76044
rect 90508 76032 90514 76084
rect 90821 76075 90879 76081
rect 90821 76041 90833 76075
rect 90867 76072 90879 76075
rect 93486 76072 93492 76084
rect 90867 76044 93492 76072
rect 90867 76041 90879 76044
rect 90821 76035 90879 76041
rect 93486 76032 93492 76044
rect 93544 76032 93550 76084
rect 96893 76075 96951 76081
rect 96893 76041 96905 76075
rect 96939 76072 96951 76075
rect 100570 76072 100576 76084
rect 96939 76044 100576 76072
rect 96939 76041 96951 76044
rect 96893 76035 96951 76041
rect 100570 76032 100576 76044
rect 100628 76032 100634 76084
rect 100754 76032 100760 76084
rect 100812 76032 100818 76084
rect 108390 76032 108396 76084
rect 108448 76032 108454 76084
rect 64230 75964 64236 76016
rect 64288 76004 64294 76016
rect 70118 76004 70124 76016
rect 64288 75976 70124 76004
rect 64288 75964 64294 75976
rect 70118 75964 70124 75976
rect 70176 75964 70182 76016
rect 90266 75964 90272 76016
rect 90324 75964 90330 76016
rect 93394 76004 93400 76016
rect 90652 75976 93400 76004
rect 16485 75939 16543 75945
rect 14608 75908 14688 75936
rect 14608 75896 14614 75908
rect 14660 75868 14688 75908
rect 16485 75905 16497 75939
rect 16531 75936 16543 75939
rect 16531 75908 16896 75936
rect 16531 75905 16543 75908
rect 16485 75899 16543 75905
rect 14737 75871 14795 75877
rect 14737 75868 14749 75871
rect 14660 75840 14749 75868
rect 14737 75837 14749 75840
rect 14783 75837 14795 75871
rect 14737 75831 14795 75837
rect 16209 75871 16267 75877
rect 16209 75837 16221 75871
rect 16255 75868 16267 75871
rect 16868 75868 16896 75908
rect 83458 75896 83464 75948
rect 83516 75936 83522 75948
rect 90652 75936 90680 75976
rect 93394 75964 93400 75976
rect 93452 75964 93458 76016
rect 94038 75964 94044 76016
rect 94096 76004 94102 76016
rect 94096 75976 95910 76004
rect 94096 75964 94102 75976
rect 98454 75964 98460 76016
rect 98512 76004 98518 76016
rect 99469 76007 99527 76013
rect 99469 76004 99481 76007
rect 98512 75976 99481 76004
rect 98512 75964 98518 75976
rect 83516 75908 90680 75936
rect 90729 75939 90787 75945
rect 83516 75896 83522 75908
rect 90729 75905 90741 75939
rect 90775 75936 90787 75939
rect 91097 75939 91155 75945
rect 91097 75936 91109 75939
rect 90775 75908 91109 75936
rect 90775 75905 90787 75908
rect 90729 75899 90787 75905
rect 91097 75905 91109 75908
rect 91143 75936 91155 75939
rect 91186 75936 91192 75948
rect 91143 75908 91192 75936
rect 91143 75905 91155 75908
rect 91097 75899 91155 75905
rect 91186 75896 91192 75908
rect 91244 75896 91250 75948
rect 96890 75896 96896 75948
rect 96948 75936 96954 75948
rect 97718 75936 97724 75948
rect 96948 75908 97724 75936
rect 96948 75896 96954 75908
rect 97718 75896 97724 75908
rect 97776 75936 97782 75948
rect 98273 75939 98331 75945
rect 98273 75936 98285 75939
rect 97776 75908 98285 75936
rect 97776 75896 97782 75908
rect 98273 75905 98285 75908
rect 98319 75905 98331 75939
rect 98273 75899 98331 75905
rect 18046 75868 18052 75880
rect 16255 75840 16804 75868
rect 16868 75840 18052 75868
rect 16255 75837 16267 75840
rect 16209 75831 16267 75837
rect 16776 75800 16804 75840
rect 18046 75828 18052 75840
rect 18104 75828 18110 75880
rect 95145 75871 95203 75877
rect 95145 75837 95157 75871
rect 95191 75837 95203 75871
rect 95145 75831 95203 75837
rect 19334 75800 19340 75812
rect 16776 75772 19340 75800
rect 19334 75760 19340 75772
rect 19392 75760 19398 75812
rect 88153 75803 88211 75809
rect 88153 75769 88165 75803
rect 88199 75800 88211 75803
rect 88242 75800 88248 75812
rect 88199 75772 88248 75800
rect 88199 75769 88211 75772
rect 88153 75763 88211 75769
rect 88242 75760 88248 75772
rect 88300 75800 88306 75812
rect 88889 75803 88947 75809
rect 88889 75800 88901 75803
rect 88300 75772 88901 75800
rect 88300 75760 88306 75772
rect 88889 75769 88901 75772
rect 88935 75800 88947 75803
rect 89714 75800 89720 75812
rect 88935 75772 89720 75800
rect 88935 75769 88947 75772
rect 88889 75763 88947 75769
rect 89714 75760 89720 75772
rect 89772 75760 89778 75812
rect 1486 75692 1492 75744
rect 1544 75692 1550 75744
rect 87969 75735 88027 75741
rect 87969 75701 87981 75735
rect 88015 75732 88027 75735
rect 88058 75732 88064 75744
rect 88015 75704 88064 75732
rect 88015 75701 88027 75704
rect 87969 75695 88027 75701
rect 88058 75692 88064 75704
rect 88116 75692 88122 75744
rect 89898 75692 89904 75744
rect 89956 75692 89962 75744
rect 90082 75692 90088 75744
rect 90140 75692 90146 75744
rect 92566 75692 92572 75744
rect 92624 75732 92630 75744
rect 94961 75735 95019 75741
rect 94961 75732 94973 75735
rect 92624 75704 94973 75732
rect 92624 75692 92630 75704
rect 94961 75701 94973 75704
rect 95007 75732 95019 75735
rect 95160 75732 95188 75831
rect 95418 75828 95424 75880
rect 95476 75828 95482 75880
rect 97813 75871 97871 75877
rect 97813 75837 97825 75871
rect 97859 75837 97871 75871
rect 97813 75831 97871 75837
rect 97905 75871 97963 75877
rect 97905 75837 97917 75871
rect 97951 75868 97963 75871
rect 97994 75868 98000 75880
rect 97951 75840 98000 75868
rect 97951 75837 97963 75840
rect 97905 75831 97963 75837
rect 97828 75800 97856 75831
rect 97994 75828 98000 75840
rect 98052 75828 98058 75880
rect 98288 75868 98316 75899
rect 98546 75896 98552 75948
rect 98604 75896 98610 75948
rect 98638 75896 98644 75948
rect 98696 75896 98702 75948
rect 98730 75896 98736 75948
rect 98788 75896 98794 75948
rect 98932 75945 98960 75976
rect 99469 75973 99481 75976
rect 99515 75973 99527 76007
rect 99469 75967 99527 75973
rect 98917 75939 98975 75945
rect 98917 75905 98929 75939
rect 98963 75905 98975 75939
rect 98917 75899 98975 75905
rect 99006 75896 99012 75948
rect 99064 75936 99070 75948
rect 99253 75939 99311 75945
rect 99253 75936 99265 75939
rect 99064 75908 99265 75936
rect 99064 75896 99070 75908
rect 99253 75905 99265 75908
rect 99299 75905 99311 75939
rect 99253 75899 99311 75905
rect 99377 75939 99435 75945
rect 99377 75905 99389 75939
rect 99423 75905 99435 75939
rect 99377 75899 99435 75905
rect 98454 75868 98460 75880
rect 98288 75840 98460 75868
rect 98454 75828 98460 75840
rect 98512 75828 98518 75880
rect 98564 75868 98592 75896
rect 99024 75868 99052 75896
rect 98564 75840 99052 75868
rect 98178 75800 98184 75812
rect 97828 75772 98184 75800
rect 98178 75760 98184 75772
rect 98236 75760 98242 75812
rect 98638 75760 98644 75812
rect 98696 75800 98702 75812
rect 99392 75800 99420 75899
rect 99558 75896 99564 75948
rect 99616 75936 99622 75948
rect 99653 75939 99711 75945
rect 99653 75936 99665 75939
rect 99616 75908 99665 75936
rect 99616 75896 99622 75908
rect 99653 75905 99665 75908
rect 99699 75905 99711 75939
rect 99653 75899 99711 75905
rect 99745 75939 99803 75945
rect 99745 75905 99757 75939
rect 99791 75905 99803 75939
rect 99745 75899 99803 75905
rect 99760 75868 99788 75899
rect 100018 75896 100024 75948
rect 100076 75936 100082 75948
rect 100573 75939 100631 75945
rect 100573 75936 100585 75939
rect 100076 75908 100585 75936
rect 100076 75896 100082 75908
rect 100573 75905 100585 75908
rect 100619 75905 100631 75939
rect 108209 75939 108267 75945
rect 108209 75936 108221 75939
rect 100573 75899 100631 75905
rect 108040 75908 108221 75936
rect 100202 75868 100208 75880
rect 99760 75840 100208 75868
rect 100202 75828 100208 75840
rect 100260 75828 100266 75880
rect 100386 75828 100392 75880
rect 100444 75828 100450 75880
rect 101674 75828 101680 75880
rect 101732 75868 101738 75880
rect 104066 75868 104072 75880
rect 101732 75840 104072 75868
rect 101732 75828 101738 75840
rect 104066 75828 104072 75840
rect 104124 75828 104130 75880
rect 98696 75772 99420 75800
rect 98696 75760 98702 75772
rect 100294 75760 100300 75812
rect 100352 75800 100358 75812
rect 108040 75809 108068 75908
rect 108209 75905 108221 75908
rect 108255 75905 108267 75939
rect 108209 75899 108267 75905
rect 108025 75803 108083 75809
rect 108025 75800 108037 75803
rect 100352 75772 108037 75800
rect 100352 75760 100358 75772
rect 108025 75769 108037 75772
rect 108071 75769 108083 75803
rect 108025 75763 108083 75769
rect 95007 75704 95188 75732
rect 95007 75701 95019 75704
rect 94961 75695 95019 75701
rect 97534 75692 97540 75744
rect 97592 75732 97598 75744
rect 97629 75735 97687 75741
rect 97629 75732 97641 75735
rect 97592 75704 97641 75732
rect 97592 75692 97598 75704
rect 97629 75701 97641 75704
rect 97675 75701 97687 75735
rect 97629 75695 97687 75701
rect 98362 75692 98368 75744
rect 98420 75692 98426 75744
rect 99098 75692 99104 75744
rect 99156 75692 99162 75744
rect 99190 75692 99196 75744
rect 99248 75732 99254 75744
rect 107930 75732 107936 75744
rect 99248 75704 107936 75732
rect 99248 75692 99254 75704
rect 107930 75692 107936 75704
rect 107988 75692 107994 75744
rect 1104 75642 108836 75664
rect 1104 75590 4214 75642
rect 4266 75590 4278 75642
rect 4330 75590 4342 75642
rect 4394 75590 4406 75642
rect 4458 75590 4470 75642
rect 4522 75590 34934 75642
rect 34986 75590 34998 75642
rect 35050 75590 35062 75642
rect 35114 75590 35126 75642
rect 35178 75590 35190 75642
rect 35242 75590 65654 75642
rect 65706 75590 65718 75642
rect 65770 75590 65782 75642
rect 65834 75590 65846 75642
rect 65898 75590 65910 75642
rect 65962 75590 96374 75642
rect 96426 75590 96438 75642
rect 96490 75590 96502 75642
rect 96554 75590 96566 75642
rect 96618 75590 96630 75642
rect 96682 75590 108836 75642
rect 1104 75568 108836 75590
rect 22278 75488 22284 75540
rect 22336 75488 22342 75540
rect 90266 75528 90272 75540
rect 87708 75500 90272 75528
rect 87708 75469 87736 75500
rect 90266 75488 90272 75500
rect 90324 75528 90330 75540
rect 91002 75528 91008 75540
rect 90324 75500 91008 75528
rect 90324 75488 90330 75500
rect 91002 75488 91008 75500
rect 91060 75488 91066 75540
rect 94869 75531 94927 75537
rect 94869 75497 94881 75531
rect 94915 75528 94927 75531
rect 96798 75528 96804 75540
rect 94915 75500 96804 75528
rect 94915 75497 94927 75500
rect 94869 75491 94927 75497
rect 96798 75488 96804 75500
rect 96856 75488 96862 75540
rect 97994 75488 98000 75540
rect 98052 75528 98058 75540
rect 98052 75500 98592 75528
rect 98052 75488 98058 75500
rect 87693 75463 87751 75469
rect 87693 75429 87705 75463
rect 87739 75429 87751 75463
rect 87693 75423 87751 75429
rect 88242 75420 88248 75472
rect 88300 75460 88306 75472
rect 88337 75463 88395 75469
rect 88337 75460 88349 75463
rect 88300 75432 88349 75460
rect 88300 75420 88306 75432
rect 88337 75429 88349 75432
rect 88383 75429 88395 75463
rect 88337 75423 88395 75429
rect 97718 75420 97724 75472
rect 97776 75460 97782 75472
rect 98089 75463 98147 75469
rect 98089 75460 98101 75463
rect 97776 75432 98101 75460
rect 97776 75420 97782 75432
rect 98089 75429 98101 75432
rect 98135 75429 98147 75463
rect 98564 75460 98592 75500
rect 98638 75488 98644 75540
rect 98696 75528 98702 75540
rect 99009 75531 99067 75537
rect 99009 75528 99021 75531
rect 98696 75500 99021 75528
rect 98696 75488 98702 75500
rect 99009 75497 99021 75500
rect 99055 75497 99067 75531
rect 99009 75491 99067 75497
rect 99190 75488 99196 75540
rect 99248 75528 99254 75540
rect 101674 75528 101680 75540
rect 99248 75500 101680 75528
rect 99248 75488 99254 75500
rect 101674 75488 101680 75500
rect 101732 75488 101738 75540
rect 102873 75531 102931 75537
rect 102873 75497 102885 75531
rect 102919 75528 102931 75531
rect 103241 75531 103299 75537
rect 103241 75528 103253 75531
rect 102919 75500 103253 75528
rect 102919 75497 102931 75500
rect 102873 75491 102931 75497
rect 103241 75497 103253 75500
rect 103287 75528 103299 75531
rect 103287 75500 103836 75528
rect 103287 75497 103299 75500
rect 103241 75491 103299 75497
rect 99282 75460 99288 75472
rect 98564 75432 99288 75460
rect 98089 75423 98147 75429
rect 99282 75420 99288 75432
rect 99340 75460 99346 75472
rect 100757 75463 100815 75469
rect 100757 75460 100769 75463
rect 99340 75432 100769 75460
rect 99340 75420 99346 75432
rect 100757 75429 100769 75432
rect 100803 75429 100815 75463
rect 100757 75423 100815 75429
rect 103514 75420 103520 75472
rect 103572 75420 103578 75472
rect 87969 75395 88027 75401
rect 87969 75361 87981 75395
rect 88015 75392 88027 75395
rect 88260 75392 88288 75420
rect 88015 75364 88288 75392
rect 88720 75364 90956 75392
rect 88015 75361 88027 75364
rect 87969 75355 88027 75361
rect 1673 75327 1731 75333
rect 1673 75293 1685 75327
rect 1719 75324 1731 75327
rect 18138 75324 18144 75336
rect 1719 75296 18144 75324
rect 1719 75293 1731 75296
rect 1673 75287 1731 75293
rect 18138 75284 18144 75296
rect 18196 75284 18202 75336
rect 22370 75284 22376 75336
rect 22428 75284 22434 75336
rect 25593 75327 25651 75333
rect 25593 75293 25605 75327
rect 25639 75293 25651 75327
rect 25593 75287 25651 75293
rect 19150 75216 19156 75268
rect 19208 75256 19214 75268
rect 25501 75259 25559 75265
rect 25501 75256 25513 75259
rect 19208 75228 25513 75256
rect 19208 75216 19214 75228
rect 25501 75225 25513 75228
rect 25547 75225 25559 75259
rect 25501 75219 25559 75225
rect 842 75148 848 75200
rect 900 75188 906 75200
rect 1489 75191 1547 75197
rect 1489 75188 1501 75191
rect 900 75160 1501 75188
rect 900 75148 906 75160
rect 1489 75157 1501 75160
rect 1535 75157 1547 75191
rect 1489 75151 1547 75157
rect 22370 75148 22376 75200
rect 22428 75188 22434 75200
rect 22557 75191 22615 75197
rect 22557 75188 22569 75191
rect 22428 75160 22569 75188
rect 22428 75148 22434 75160
rect 22557 75157 22569 75160
rect 22603 75188 22615 75191
rect 24762 75188 24768 75200
rect 22603 75160 24768 75188
rect 22603 75157 22615 75160
rect 22557 75151 22615 75157
rect 24762 75148 24768 75160
rect 24820 75188 24826 75200
rect 25608 75188 25636 75287
rect 86862 75284 86868 75336
rect 86920 75324 86926 75336
rect 88720 75333 88748 75364
rect 88705 75327 88763 75333
rect 88705 75324 88717 75327
rect 86920 75296 88717 75324
rect 86920 75284 86926 75296
rect 88705 75293 88717 75296
rect 88751 75293 88763 75327
rect 88705 75287 88763 75293
rect 88150 75216 88156 75268
rect 88208 75216 88214 75268
rect 88981 75259 89039 75265
rect 88981 75225 88993 75259
rect 89027 75225 89039 75259
rect 88981 75219 89039 75225
rect 25685 75191 25743 75197
rect 25685 75188 25697 75191
rect 24820 75160 25697 75188
rect 24820 75148 24826 75160
rect 25685 75157 25697 75160
rect 25731 75157 25743 75191
rect 25685 75151 25743 75157
rect 87509 75191 87567 75197
rect 87509 75157 87521 75191
rect 87555 75188 87567 75191
rect 87782 75188 87788 75200
rect 87555 75160 87788 75188
rect 87555 75157 87567 75160
rect 87509 75151 87567 75157
rect 87782 75148 87788 75160
rect 87840 75148 87846 75200
rect 88996 75188 89024 75219
rect 89622 75216 89628 75268
rect 89680 75216 89686 75268
rect 90726 75216 90732 75268
rect 90784 75216 90790 75268
rect 89898 75188 89904 75200
rect 88996 75160 89904 75188
rect 89898 75148 89904 75160
rect 89956 75148 89962 75200
rect 90928 75197 90956 75364
rect 93394 75352 93400 75404
rect 93452 75352 93458 75404
rect 96890 75352 96896 75404
rect 96948 75392 96954 75404
rect 97169 75395 97227 75401
rect 97169 75392 97181 75395
rect 96948 75364 97181 75392
rect 96948 75352 96954 75364
rect 97169 75361 97181 75364
rect 97215 75361 97227 75395
rect 97169 75355 97227 75361
rect 97920 75364 99144 75392
rect 93121 75327 93179 75333
rect 93121 75324 93133 75327
rect 92952 75296 93133 75324
rect 91462 75216 91468 75268
rect 91520 75256 91526 75268
rect 92382 75256 92388 75268
rect 91520 75228 92388 75256
rect 91520 75216 91526 75228
rect 92382 75216 92388 75228
rect 92440 75216 92446 75268
rect 90913 75191 90971 75197
rect 90913 75157 90925 75191
rect 90959 75188 90971 75191
rect 91370 75188 91376 75200
rect 90959 75160 91376 75188
rect 90959 75157 90971 75160
rect 90913 75151 90971 75157
rect 91370 75148 91376 75160
rect 91428 75188 91434 75200
rect 92566 75188 92572 75200
rect 91428 75160 92572 75188
rect 91428 75148 91434 75160
rect 92566 75148 92572 75160
rect 92624 75188 92630 75200
rect 92952 75197 92980 75296
rect 93121 75293 93133 75296
rect 93167 75293 93179 75327
rect 93121 75287 93179 75293
rect 97920 75268 97948 75364
rect 98270 75284 98276 75336
rect 98328 75284 98334 75336
rect 98362 75284 98368 75336
rect 98420 75284 98426 75336
rect 99116 75333 99144 75364
rect 100938 75352 100944 75404
rect 100996 75392 101002 75404
rect 101309 75395 101367 75401
rect 101309 75392 101321 75395
rect 100996 75364 101321 75392
rect 100996 75352 101002 75364
rect 101309 75361 101321 75364
rect 101355 75392 101367 75395
rect 101398 75392 101404 75404
rect 101355 75364 101404 75392
rect 101355 75361 101367 75364
rect 101309 75355 101367 75361
rect 101398 75352 101404 75364
rect 101456 75352 101462 75404
rect 101950 75352 101956 75404
rect 102008 75352 102014 75404
rect 103146 75392 103152 75404
rect 102796 75364 103152 75392
rect 98917 75327 98975 75333
rect 98917 75293 98929 75327
rect 98963 75293 98975 75327
rect 98917 75287 98975 75293
rect 99101 75327 99159 75333
rect 99101 75293 99113 75327
rect 99147 75324 99159 75327
rect 99374 75324 99380 75336
rect 99147 75296 99380 75324
rect 99147 75293 99159 75296
rect 99101 75287 99159 75293
rect 93026 75216 93032 75268
rect 93084 75256 93090 75268
rect 97902 75256 97908 75268
rect 93084 75228 93886 75256
rect 97368 75228 97908 75256
rect 93084 75216 93090 75228
rect 92937 75191 92995 75197
rect 92937 75188 92949 75191
rect 92624 75160 92949 75188
rect 92624 75148 92630 75160
rect 92937 75157 92949 75160
rect 92983 75157 92995 75191
rect 92937 75151 92995 75157
rect 96798 75148 96804 75200
rect 96856 75188 96862 75200
rect 97368 75197 97396 75228
rect 97902 75216 97908 75228
rect 97960 75216 97966 75268
rect 98089 75259 98147 75265
rect 98089 75225 98101 75259
rect 98135 75256 98147 75259
rect 98730 75256 98736 75268
rect 98135 75228 98736 75256
rect 98135 75225 98147 75228
rect 98089 75219 98147 75225
rect 98730 75216 98736 75228
rect 98788 75216 98794 75268
rect 98932 75256 98960 75287
rect 99374 75284 99380 75296
rect 99432 75284 99438 75336
rect 100018 75284 100024 75336
rect 100076 75324 100082 75336
rect 102796 75333 102824 75364
rect 103146 75352 103152 75364
rect 103204 75352 103210 75404
rect 103330 75352 103336 75404
rect 103388 75392 103394 75404
rect 103388 75364 103744 75392
rect 103388 75352 103394 75364
rect 100297 75327 100355 75333
rect 100297 75324 100309 75327
rect 100076 75296 100309 75324
rect 100076 75284 100082 75296
rect 100297 75293 100309 75296
rect 100343 75293 100355 75327
rect 100297 75287 100355 75293
rect 100481 75327 100539 75333
rect 100481 75293 100493 75327
rect 100527 75293 100539 75327
rect 102045 75327 102103 75333
rect 102045 75324 102057 75327
rect 100481 75287 100539 75293
rect 101968 75296 102057 75324
rect 99466 75256 99472 75268
rect 98932 75228 99472 75256
rect 99466 75216 99472 75228
rect 99524 75216 99530 75268
rect 99926 75216 99932 75268
rect 99984 75256 99990 75268
rect 100386 75256 100392 75268
rect 99984 75228 100392 75256
rect 99984 75216 99990 75228
rect 100386 75216 100392 75228
rect 100444 75256 100450 75268
rect 100496 75256 100524 75287
rect 101968 75268 101996 75296
rect 102045 75293 102057 75296
rect 102091 75293 102103 75327
rect 102045 75287 102103 75293
rect 102781 75327 102839 75333
rect 102781 75293 102793 75327
rect 102827 75293 102839 75327
rect 102781 75287 102839 75293
rect 102962 75284 102968 75336
rect 103020 75284 103026 75336
rect 100444 75228 100524 75256
rect 101125 75259 101183 75265
rect 100444 75216 100450 75228
rect 101125 75225 101137 75259
rect 101171 75256 101183 75259
rect 101171 75228 101720 75256
rect 101171 75225 101183 75228
rect 101125 75219 101183 75225
rect 97353 75191 97411 75197
rect 97353 75188 97365 75191
rect 96856 75160 97365 75188
rect 96856 75148 96862 75160
rect 97353 75157 97365 75160
rect 97399 75157 97411 75191
rect 97353 75151 97411 75157
rect 97442 75148 97448 75200
rect 97500 75148 97506 75200
rect 97813 75191 97871 75197
rect 97813 75157 97825 75191
rect 97859 75188 97871 75191
rect 97994 75188 98000 75200
rect 97859 75160 98000 75188
rect 97859 75157 97871 75160
rect 97813 75151 97871 75157
rect 97994 75148 98000 75160
rect 98052 75148 98058 75200
rect 98178 75148 98184 75200
rect 98236 75188 98242 75200
rect 100294 75188 100300 75200
rect 98236 75160 100300 75188
rect 98236 75148 98242 75160
rect 100294 75148 100300 75160
rect 100352 75148 100358 75200
rect 100478 75148 100484 75200
rect 100536 75148 100542 75200
rect 101214 75148 101220 75200
rect 101272 75148 101278 75200
rect 101692 75197 101720 75228
rect 101950 75216 101956 75268
rect 102008 75216 102014 75268
rect 102870 75216 102876 75268
rect 102928 75256 102934 75268
rect 103209 75259 103267 75265
rect 103209 75256 103221 75259
rect 102928 75228 103221 75256
rect 102928 75216 102934 75228
rect 103209 75225 103221 75228
rect 103255 75256 103267 75259
rect 103255 75225 103284 75256
rect 103209 75219 103284 75225
rect 101677 75191 101735 75197
rect 101677 75157 101689 75191
rect 101723 75157 101735 75191
rect 101677 75151 101735 75157
rect 103054 75148 103060 75200
rect 103112 75148 103118 75200
rect 103256 75188 103284 75219
rect 103330 75216 103336 75268
rect 103388 75256 103394 75268
rect 103716 75265 103744 75364
rect 103808 75333 103836 75500
rect 104158 75488 104164 75540
rect 104216 75528 104222 75540
rect 104621 75531 104679 75537
rect 104621 75528 104633 75531
rect 104216 75500 104633 75528
rect 104216 75488 104222 75500
rect 104621 75497 104633 75500
rect 104667 75497 104679 75531
rect 104621 75491 104679 75497
rect 104802 75488 104808 75540
rect 104860 75528 104866 75540
rect 108025 75531 108083 75537
rect 108025 75528 108037 75531
rect 104860 75500 108037 75528
rect 104860 75488 104866 75500
rect 108025 75497 108037 75500
rect 108071 75497 108083 75531
rect 108025 75491 108083 75497
rect 103974 75420 103980 75472
rect 104032 75460 104038 75472
rect 104989 75463 105047 75469
rect 104989 75460 105001 75463
rect 104032 75432 105001 75460
rect 104032 75420 104038 75432
rect 104989 75429 105001 75432
rect 105035 75429 105047 75463
rect 104989 75423 105047 75429
rect 103992 75364 104848 75392
rect 103992 75333 104020 75364
rect 103793 75327 103851 75333
rect 103793 75293 103805 75327
rect 103839 75293 103851 75327
rect 103793 75287 103851 75293
rect 103885 75327 103943 75333
rect 103885 75293 103897 75327
rect 103931 75293 103943 75327
rect 103885 75287 103943 75293
rect 103977 75327 104035 75333
rect 103977 75293 103989 75327
rect 104023 75293 104035 75327
rect 103977 75287 104035 75293
rect 103425 75259 103483 75265
rect 103425 75256 103437 75259
rect 103388 75228 103437 75256
rect 103388 75216 103394 75228
rect 103425 75225 103437 75228
rect 103471 75225 103483 75259
rect 103425 75219 103483 75225
rect 103517 75259 103575 75265
rect 103517 75225 103529 75259
rect 103563 75225 103575 75259
rect 103517 75219 103575 75225
rect 103701 75259 103759 75265
rect 103701 75225 103713 75259
rect 103747 75225 103759 75259
rect 103900 75256 103928 75287
rect 104158 75284 104164 75336
rect 104216 75284 104222 75336
rect 104820 75324 104848 75364
rect 105096 75364 105400 75392
rect 105096 75333 105124 75364
rect 105372 75333 105400 75364
rect 105081 75327 105139 75333
rect 105081 75324 105093 75327
rect 104820 75296 105093 75324
rect 104066 75256 104072 75268
rect 103900 75228 104072 75256
rect 103701 75219 103759 75225
rect 103532 75188 103560 75219
rect 104066 75216 104072 75228
rect 104124 75256 104130 75268
rect 104820 75265 104848 75296
rect 105081 75293 105093 75296
rect 105127 75293 105139 75327
rect 105081 75287 105139 75293
rect 105173 75327 105231 75333
rect 105173 75293 105185 75327
rect 105219 75293 105231 75327
rect 105173 75287 105231 75293
rect 105357 75327 105415 75333
rect 105357 75293 105369 75327
rect 105403 75324 105415 75327
rect 107746 75324 107752 75336
rect 105403 75296 107752 75324
rect 105403 75293 105415 75296
rect 105357 75287 105415 75293
rect 104805 75259 104863 75265
rect 104124 75228 104572 75256
rect 104124 75216 104130 75228
rect 103256 75160 103560 75188
rect 104342 75148 104348 75200
rect 104400 75148 104406 75200
rect 104434 75148 104440 75200
rect 104492 75148 104498 75200
rect 104544 75188 104572 75228
rect 104805 75225 104817 75259
rect 104851 75225 104863 75259
rect 105188 75256 105216 75287
rect 107746 75284 107752 75296
rect 107804 75284 107810 75336
rect 108040 75324 108068 75491
rect 108209 75327 108267 75333
rect 108209 75324 108221 75327
rect 108040 75296 108221 75324
rect 108209 75293 108221 75296
rect 108255 75293 108267 75327
rect 108209 75287 108267 75293
rect 104805 75219 104863 75225
rect 104912 75228 105216 75256
rect 104605 75191 104663 75197
rect 104605 75188 104617 75191
rect 104544 75160 104617 75188
rect 104605 75157 104617 75160
rect 104651 75188 104663 75191
rect 104912 75188 104940 75228
rect 104651 75160 104940 75188
rect 104651 75157 104663 75160
rect 104605 75151 104663 75157
rect 105262 75148 105268 75200
rect 105320 75148 105326 75200
rect 108390 75148 108396 75200
rect 108448 75148 108454 75200
rect 1104 75098 108836 75120
rect 1104 75046 4874 75098
rect 4926 75046 4938 75098
rect 4990 75046 5002 75098
rect 5054 75046 5066 75098
rect 5118 75046 5130 75098
rect 5182 75046 35594 75098
rect 35646 75046 35658 75098
rect 35710 75046 35722 75098
rect 35774 75046 35786 75098
rect 35838 75046 35850 75098
rect 35902 75046 66314 75098
rect 66366 75046 66378 75098
rect 66430 75046 66442 75098
rect 66494 75046 66506 75098
rect 66558 75046 66570 75098
rect 66622 75046 97034 75098
rect 97086 75046 97098 75098
rect 97150 75046 97162 75098
rect 97214 75046 97226 75098
rect 97278 75046 97290 75098
rect 97342 75046 108836 75098
rect 1104 75024 108836 75046
rect 18046 74944 18052 74996
rect 18104 74984 18110 74996
rect 18966 74984 18972 74996
rect 18104 74956 18972 74984
rect 18104 74944 18110 74956
rect 18966 74944 18972 74956
rect 19024 74984 19030 74996
rect 19886 74984 19892 74996
rect 19024 74956 19892 74984
rect 19024 74944 19030 74956
rect 19886 74944 19892 74956
rect 19944 74944 19950 74996
rect 86862 74944 86868 74996
rect 86920 74984 86926 74996
rect 86920 74956 88012 74984
rect 86920 74944 86926 74956
rect 19150 74876 19156 74928
rect 19208 74876 19214 74928
rect 85666 74876 85672 74928
rect 85724 74916 85730 74928
rect 85724 74888 86618 74916
rect 85724 74876 85730 74888
rect 87782 74876 87788 74928
rect 87840 74876 87846 74928
rect 87984 74916 88012 74956
rect 88150 74944 88156 74996
rect 88208 74984 88214 74996
rect 88245 74987 88303 74993
rect 88245 74984 88257 74987
rect 88208 74956 88257 74984
rect 88208 74944 88214 74956
rect 88245 74953 88257 74956
rect 88291 74984 88303 74987
rect 88702 74984 88708 74996
rect 88291 74956 88708 74984
rect 88291 74953 88303 74956
rect 88245 74947 88303 74953
rect 88702 74944 88708 74956
rect 88760 74944 88766 74996
rect 89622 74944 89628 74996
rect 89680 74944 89686 74996
rect 89714 74944 89720 74996
rect 89772 74984 89778 74996
rect 90913 74987 90971 74993
rect 90913 74984 90925 74987
rect 89772 74956 90925 74984
rect 89772 74944 89778 74956
rect 90913 74953 90925 74956
rect 90959 74984 90971 74987
rect 91649 74987 91707 74993
rect 91649 74984 91661 74987
rect 90959 74956 91661 74984
rect 90959 74953 90971 74956
rect 90913 74947 90971 74953
rect 91649 74953 91661 74956
rect 91695 74984 91707 74987
rect 91830 74984 91836 74996
rect 91695 74956 91836 74984
rect 91695 74953 91707 74956
rect 91649 74947 91707 74953
rect 91830 74944 91836 74956
rect 91888 74984 91894 74996
rect 92201 74987 92259 74993
rect 92201 74984 92213 74987
rect 91888 74956 92213 74984
rect 91888 74944 91894 74956
rect 92201 74953 92213 74956
rect 92247 74984 92259 74987
rect 93302 74984 93308 74996
rect 92247 74956 93308 74984
rect 92247 74953 92259 74956
rect 92201 74947 92259 74953
rect 93302 74944 93308 74956
rect 93360 74944 93366 74996
rect 96890 74984 96896 74996
rect 94516 74956 96896 74984
rect 88334 74916 88340 74928
rect 87984 74888 88340 74916
rect 19886 74808 19892 74860
rect 19944 74808 19950 74860
rect 88076 74857 88104 74888
rect 88334 74876 88340 74888
rect 88392 74876 88398 74928
rect 93946 74916 93952 74928
rect 89824 74888 93952 74916
rect 89824 74857 89852 74888
rect 93946 74876 93952 74888
rect 94004 74876 94010 74928
rect 88061 74851 88119 74857
rect 88061 74817 88073 74851
rect 88107 74817 88119 74851
rect 89533 74851 89591 74857
rect 89533 74848 89545 74851
rect 88061 74811 88119 74817
rect 88536 74820 89545 74848
rect 18138 74740 18144 74792
rect 18196 74740 18202 74792
rect 19613 74783 19671 74789
rect 19613 74749 19625 74783
rect 19659 74780 19671 74783
rect 28534 74780 28540 74792
rect 19659 74752 28540 74780
rect 19659 74749 19671 74752
rect 19613 74743 19671 74749
rect 28534 74740 28540 74752
rect 28592 74740 28598 74792
rect 86037 74783 86095 74789
rect 86037 74749 86049 74783
rect 86083 74780 86095 74783
rect 88150 74780 88156 74792
rect 86083 74752 88156 74780
rect 86083 74749 86095 74752
rect 86037 74743 86095 74749
rect 88150 74740 88156 74752
rect 88208 74740 88214 74792
rect 85942 74604 85948 74656
rect 86000 74644 86006 74656
rect 88536 74644 88564 74820
rect 89533 74817 89545 74820
rect 89579 74848 89591 74851
rect 89809 74851 89867 74857
rect 89809 74848 89821 74851
rect 89579 74820 89821 74848
rect 89579 74817 89591 74820
rect 89533 74811 89591 74817
rect 89809 74817 89821 74820
rect 89855 74817 89867 74851
rect 89809 74811 89867 74817
rect 91189 74851 91247 74857
rect 91189 74817 91201 74851
rect 91235 74848 91247 74851
rect 91462 74848 91468 74860
rect 91235 74820 91468 74848
rect 91235 74817 91247 74820
rect 91189 74811 91247 74817
rect 91462 74808 91468 74820
rect 91520 74808 91526 74860
rect 91741 74851 91799 74857
rect 91741 74817 91753 74851
rect 91787 74817 91799 74851
rect 91741 74811 91799 74817
rect 89441 74783 89499 74789
rect 89441 74749 89453 74783
rect 89487 74780 89499 74783
rect 89898 74780 89904 74792
rect 89487 74752 89904 74780
rect 89487 74749 89499 74752
rect 89441 74743 89499 74749
rect 89898 74740 89904 74752
rect 89956 74780 89962 74792
rect 90726 74780 90732 74792
rect 89956 74752 90732 74780
rect 89956 74740 89962 74752
rect 90726 74740 90732 74752
rect 90784 74780 90790 74792
rect 91756 74780 91784 74811
rect 91830 74808 91836 74860
rect 91888 74808 91894 74860
rect 91925 74851 91983 74857
rect 91925 74817 91937 74851
rect 91971 74817 91983 74851
rect 91925 74811 91983 74817
rect 92109 74851 92167 74857
rect 92109 74817 92121 74851
rect 92155 74848 92167 74851
rect 92382 74848 92388 74860
rect 92155 74820 92388 74848
rect 92155 74817 92167 74820
rect 92109 74811 92167 74817
rect 91940 74780 91968 74811
rect 92382 74808 92388 74820
rect 92440 74808 92446 74860
rect 94038 74808 94044 74860
rect 94096 74848 94102 74860
rect 94409 74851 94467 74857
rect 94409 74848 94421 74851
rect 94096 74820 94421 74848
rect 94096 74808 94102 74820
rect 94409 74817 94421 74820
rect 94455 74817 94467 74851
rect 94409 74811 94467 74817
rect 94056 74780 94084 74808
rect 94516 74789 94544 74956
rect 96890 74944 96896 74956
rect 96948 74944 96954 74996
rect 96985 74987 97043 74993
rect 96985 74953 96997 74987
rect 97031 74984 97043 74987
rect 97442 74984 97448 74996
rect 97031 74956 97448 74984
rect 97031 74953 97043 74956
rect 96985 74947 97043 74953
rect 97442 74944 97448 74956
rect 97500 74944 97506 74996
rect 97902 74944 97908 74996
rect 97960 74984 97966 74996
rect 97960 74956 98684 74984
rect 97960 74944 97966 74956
rect 98273 74919 98331 74925
rect 96632 74888 98040 74916
rect 96632 74857 96660 74888
rect 96617 74851 96675 74857
rect 96617 74817 96629 74851
rect 96663 74817 96675 74851
rect 96617 74811 96675 74817
rect 97350 74808 97356 74860
rect 97408 74808 97414 74860
rect 97445 74851 97503 74857
rect 97445 74817 97457 74851
rect 97491 74817 97503 74851
rect 97445 74811 97503 74817
rect 90784 74752 94084 74780
rect 94501 74783 94559 74789
rect 90784 74740 90790 74752
rect 94501 74749 94513 74783
rect 94547 74749 94559 74783
rect 94501 74743 94559 74749
rect 96706 74740 96712 74792
rect 96764 74740 96770 74792
rect 97460 74780 97488 74811
rect 97534 74808 97540 74860
rect 97592 74808 97598 74860
rect 97718 74808 97724 74860
rect 97776 74808 97782 74860
rect 98012 74857 98040 74888
rect 98273 74885 98285 74919
rect 98319 74916 98331 74919
rect 98546 74916 98552 74928
rect 98319 74888 98552 74916
rect 98319 74885 98331 74888
rect 98273 74879 98331 74885
rect 98546 74876 98552 74888
rect 98604 74876 98610 74928
rect 97997 74851 98055 74857
rect 97997 74817 98009 74851
rect 98043 74848 98055 74851
rect 98362 74848 98368 74860
rect 98043 74820 98368 74848
rect 98043 74817 98055 74820
rect 97997 74811 98055 74817
rect 98362 74808 98368 74820
rect 98420 74808 98426 74860
rect 98457 74851 98515 74857
rect 98457 74817 98469 74851
rect 98503 74848 98515 74851
rect 98656 74848 98684 74956
rect 99098 74944 99104 74996
rect 99156 74984 99162 74996
rect 100021 74987 100079 74993
rect 99156 74956 99788 74984
rect 99156 74944 99162 74956
rect 99466 74916 99472 74928
rect 98748 74888 99472 74916
rect 98748 74857 98776 74888
rect 99466 74876 99472 74888
rect 99524 74876 99530 74928
rect 98503 74820 98684 74848
rect 98733 74851 98791 74857
rect 98503 74817 98515 74820
rect 98457 74811 98515 74817
rect 98733 74817 98745 74851
rect 98779 74817 98791 74851
rect 98733 74811 98791 74817
rect 99282 74808 99288 74860
rect 99340 74808 99346 74860
rect 99760 74857 99788 74956
rect 100021 74953 100033 74987
rect 100067 74984 100079 74987
rect 100110 74984 100116 74996
rect 100067 74956 100116 74984
rect 100067 74953 100079 74956
rect 100021 74947 100079 74953
rect 100110 74944 100116 74956
rect 100168 74944 100174 74996
rect 100938 74944 100944 74996
rect 100996 74993 101002 74996
rect 100996 74984 101005 74993
rect 100996 74956 101041 74984
rect 100996 74947 101005 74956
rect 100996 74944 101002 74947
rect 101214 74944 101220 74996
rect 101272 74984 101278 74996
rect 101858 74984 101864 74996
rect 101272 74956 101864 74984
rect 101272 74944 101278 74956
rect 101858 74944 101864 74956
rect 101916 74984 101922 74996
rect 101916 74956 102180 74984
rect 101916 74944 101922 74956
rect 101033 74919 101091 74925
rect 101033 74916 101045 74919
rect 100496 74888 101045 74916
rect 100496 74860 100524 74888
rect 101033 74885 101045 74888
rect 101079 74885 101091 74919
rect 101585 74919 101643 74925
rect 101585 74916 101597 74919
rect 101033 74879 101091 74885
rect 101140 74888 101597 74916
rect 101140 74860 101168 74888
rect 101585 74885 101597 74888
rect 101631 74885 101643 74919
rect 101585 74879 101643 74885
rect 99745 74851 99803 74857
rect 99745 74817 99757 74851
rect 99791 74817 99803 74851
rect 99745 74811 99803 74817
rect 99926 74808 99932 74860
rect 99984 74808 99990 74860
rect 100018 74808 100024 74860
rect 100076 74848 100082 74860
rect 100113 74851 100171 74857
rect 100113 74848 100125 74851
rect 100076 74820 100125 74848
rect 100076 74808 100082 74820
rect 100113 74817 100125 74820
rect 100159 74817 100171 74851
rect 100113 74811 100171 74817
rect 100202 74808 100208 74860
rect 100260 74808 100266 74860
rect 100294 74808 100300 74860
rect 100352 74808 100358 74860
rect 100478 74808 100484 74860
rect 100536 74808 100542 74860
rect 100573 74851 100631 74857
rect 100573 74817 100585 74851
rect 100619 74817 100631 74851
rect 100573 74811 100631 74817
rect 97902 74780 97908 74792
rect 97460 74752 97908 74780
rect 97902 74740 97908 74752
rect 97960 74740 97966 74792
rect 99190 74780 99196 74792
rect 98012 74752 99196 74780
rect 88702 74672 88708 74724
rect 88760 74712 88766 74724
rect 98012 74712 98040 74752
rect 99190 74740 99196 74752
rect 99248 74740 99254 74792
rect 99466 74740 99472 74792
rect 99524 74740 99530 74792
rect 99561 74783 99619 74789
rect 99561 74749 99573 74783
rect 99607 74749 99619 74783
rect 99561 74743 99619 74749
rect 88760 74684 98040 74712
rect 88760 74672 88766 74684
rect 98454 74672 98460 74724
rect 98512 74712 98518 74724
rect 99377 74715 99435 74721
rect 99377 74712 99389 74715
rect 98512 74684 99389 74712
rect 98512 74672 98518 74684
rect 99377 74681 99389 74684
rect 99423 74681 99435 74715
rect 99576 74712 99604 74743
rect 99834 74740 99840 74792
rect 99892 74780 99898 74792
rect 100220 74780 100248 74808
rect 99892 74752 100248 74780
rect 100588 74780 100616 74811
rect 100662 74808 100668 74860
rect 100720 74848 100726 74860
rect 100849 74851 100907 74857
rect 100849 74848 100861 74851
rect 100720 74820 100861 74848
rect 100720 74808 100726 74820
rect 100849 74817 100861 74820
rect 100895 74817 100907 74851
rect 100849 74811 100907 74817
rect 101122 74808 101128 74860
rect 101180 74808 101186 74860
rect 101398 74808 101404 74860
rect 101456 74808 101462 74860
rect 101769 74851 101827 74857
rect 101769 74817 101781 74851
rect 101815 74817 101827 74851
rect 101769 74811 101827 74817
rect 101140 74780 101168 74808
rect 100588 74752 101168 74780
rect 101784 74780 101812 74811
rect 101950 74808 101956 74860
rect 102008 74808 102014 74860
rect 102042 74808 102048 74860
rect 102100 74808 102106 74860
rect 102152 74857 102180 74956
rect 104066 74944 104072 74996
rect 104124 74944 104130 74996
rect 102962 74876 102968 74928
rect 103020 74916 103026 74928
rect 103790 74916 103796 74928
rect 103020 74888 103796 74916
rect 103020 74876 103026 74888
rect 102137 74851 102195 74857
rect 102137 74817 102149 74851
rect 102183 74817 102195 74851
rect 102137 74811 102195 74817
rect 102321 74851 102379 74857
rect 102321 74817 102333 74851
rect 102367 74817 102379 74851
rect 102321 74811 102379 74817
rect 102229 74783 102287 74789
rect 102229 74780 102241 74783
rect 101784 74752 102241 74780
rect 99892 74740 99898 74752
rect 102229 74749 102241 74752
rect 102275 74749 102287 74783
rect 102229 74743 102287 74749
rect 100202 74712 100208 74724
rect 99576 74684 100208 74712
rect 99377 74675 99435 74681
rect 100202 74672 100208 74684
rect 100260 74712 100266 74724
rect 101217 74715 101275 74721
rect 101217 74712 101229 74715
rect 100260 74684 101229 74712
rect 100260 74672 100266 74684
rect 101217 74681 101229 74684
rect 101263 74681 101275 74715
rect 102336 74712 102364 74811
rect 102502 74808 102508 74860
rect 102560 74848 102566 74860
rect 103057 74851 103115 74857
rect 103057 74848 103069 74851
rect 102560 74820 103069 74848
rect 102560 74808 102566 74820
rect 103057 74817 103069 74820
rect 103103 74817 103115 74851
rect 103057 74811 103115 74817
rect 103241 74851 103299 74857
rect 103241 74817 103253 74851
rect 103287 74817 103299 74851
rect 103241 74811 103299 74817
rect 103333 74851 103391 74857
rect 103333 74817 103345 74851
rect 103379 74848 103391 74851
rect 103422 74848 103428 74860
rect 103379 74820 103428 74848
rect 103379 74817 103391 74820
rect 103333 74811 103391 74817
rect 102870 74740 102876 74792
rect 102928 74780 102934 74792
rect 103149 74783 103207 74789
rect 103149 74780 103161 74783
rect 102928 74752 103161 74780
rect 102928 74740 102934 74752
rect 103149 74749 103161 74752
rect 103195 74749 103207 74783
rect 103256 74780 103284 74811
rect 103422 74808 103428 74820
rect 103480 74808 103486 74860
rect 103532 74857 103560 74888
rect 103790 74876 103796 74888
rect 103848 74876 103854 74928
rect 104434 74876 104440 74928
rect 104492 74876 104498 74928
rect 103517 74851 103575 74857
rect 103517 74817 103529 74851
rect 103563 74817 103575 74851
rect 103517 74811 103575 74817
rect 103701 74851 103759 74857
rect 103701 74817 103713 74851
rect 103747 74848 103759 74851
rect 103974 74848 103980 74860
rect 103747 74820 103980 74848
rect 103747 74817 103759 74820
rect 103701 74811 103759 74817
rect 103716 74780 103744 74811
rect 103974 74808 103980 74820
rect 104032 74808 104038 74860
rect 104066 74808 104072 74860
rect 104124 74848 104130 74860
rect 104802 74848 104808 74860
rect 104124 74820 104808 74848
rect 104124 74808 104130 74820
rect 104802 74808 104808 74820
rect 104860 74808 104866 74860
rect 105173 74851 105231 74857
rect 105173 74848 105185 74851
rect 104912 74820 105185 74848
rect 103256 74752 103744 74780
rect 103992 74780 104020 74808
rect 104618 74780 104624 74792
rect 103992 74752 104624 74780
rect 103149 74743 103207 74749
rect 104618 74740 104624 74752
rect 104676 74740 104682 74792
rect 104912 74789 104940 74820
rect 105173 74817 105185 74820
rect 105219 74817 105231 74851
rect 105173 74811 105231 74817
rect 104897 74783 104955 74789
rect 104897 74749 104909 74783
rect 104943 74749 104955 74783
rect 104897 74743 104955 74749
rect 104986 74740 104992 74792
rect 105044 74780 105050 74792
rect 105081 74783 105139 74789
rect 105081 74780 105093 74783
rect 105044 74752 105093 74780
rect 105044 74740 105050 74752
rect 105081 74749 105093 74752
rect 105127 74749 105139 74783
rect 105081 74743 105139 74749
rect 103698 74712 103704 74724
rect 102336 74684 103704 74712
rect 101217 74675 101275 74681
rect 103698 74672 103704 74684
rect 103756 74672 103762 74724
rect 104342 74672 104348 74724
rect 104400 74712 104406 74724
rect 104713 74715 104771 74721
rect 104713 74712 104725 74715
rect 104400 74684 104725 74712
rect 104400 74672 104406 74684
rect 104713 74681 104725 74684
rect 104759 74681 104771 74715
rect 104713 74675 104771 74681
rect 86000 74616 88564 74644
rect 86000 74604 86006 74616
rect 88978 74604 88984 74656
rect 89036 74604 89042 74656
rect 91278 74604 91284 74656
rect 91336 74604 91342 74656
rect 91462 74604 91468 74656
rect 91520 74644 91526 74656
rect 91833 74647 91891 74653
rect 91833 74644 91845 74647
rect 91520 74616 91845 74644
rect 91520 74604 91526 74616
rect 91833 74613 91845 74616
rect 91879 74613 91891 74647
rect 91833 74607 91891 74613
rect 94133 74647 94191 74653
rect 94133 74613 94145 74647
rect 94179 74644 94191 74647
rect 94406 74644 94412 74656
rect 94179 74616 94412 74644
rect 94179 74613 94191 74616
rect 94133 74607 94191 74613
rect 94406 74604 94412 74616
rect 94464 74604 94470 74656
rect 96890 74604 96896 74656
rect 96948 74644 96954 74656
rect 97077 74647 97135 74653
rect 97077 74644 97089 74647
rect 96948 74616 97089 74644
rect 96948 74604 96954 74616
rect 97077 74613 97089 74616
rect 97123 74613 97135 74647
rect 97077 74607 97135 74613
rect 97350 74604 97356 74656
rect 97408 74644 97414 74656
rect 97810 74644 97816 74656
rect 97408 74616 97816 74644
rect 97408 74604 97414 74616
rect 97810 74604 97816 74616
rect 97868 74604 97874 74656
rect 97902 74604 97908 74656
rect 97960 74644 97966 74656
rect 99101 74647 99159 74653
rect 99101 74644 99113 74647
rect 97960 74616 99113 74644
rect 97960 74604 97966 74616
rect 99101 74613 99113 74616
rect 99147 74613 99159 74647
rect 99101 74607 99159 74613
rect 99650 74604 99656 74656
rect 99708 74644 99714 74656
rect 100294 74644 100300 74656
rect 99708 74616 100300 74644
rect 99708 74604 99714 74616
rect 100294 74604 100300 74616
rect 100352 74604 100358 74656
rect 100754 74604 100760 74656
rect 100812 74604 100818 74656
rect 103146 74604 103152 74656
rect 103204 74644 103210 74656
rect 103422 74644 103428 74656
rect 103204 74616 103428 74644
rect 103204 74604 103210 74616
rect 103422 74604 103428 74616
rect 103480 74604 103486 74656
rect 103606 74604 103612 74656
rect 103664 74604 103670 74656
rect 103793 74647 103851 74653
rect 103793 74613 103805 74647
rect 103839 74644 103851 74647
rect 103974 74644 103980 74656
rect 103839 74616 103980 74644
rect 103839 74613 103851 74616
rect 103793 74607 103851 74613
rect 103974 74604 103980 74616
rect 104032 74604 104038 74656
rect 105354 74604 105360 74656
rect 105412 74644 105418 74656
rect 105449 74647 105507 74653
rect 105449 74644 105461 74647
rect 105412 74616 105461 74644
rect 105412 74604 105418 74616
rect 105449 74613 105461 74616
rect 105495 74613 105507 74647
rect 105449 74607 105507 74613
rect 1104 74554 108836 74576
rect 1104 74502 4214 74554
rect 4266 74502 4278 74554
rect 4330 74502 4342 74554
rect 4394 74502 4406 74554
rect 4458 74502 4470 74554
rect 4522 74502 34934 74554
rect 34986 74502 34998 74554
rect 35050 74502 35062 74554
rect 35114 74502 35126 74554
rect 35178 74502 35190 74554
rect 35242 74502 65654 74554
rect 65706 74502 65718 74554
rect 65770 74502 65782 74554
rect 65834 74502 65846 74554
rect 65898 74502 65910 74554
rect 65962 74502 96374 74554
rect 96426 74502 96438 74554
rect 96490 74502 96502 74554
rect 96554 74502 96566 74554
rect 96618 74502 96630 74554
rect 96682 74502 108836 74554
rect 1104 74480 108836 74502
rect 21729 74443 21787 74449
rect 21729 74409 21741 74443
rect 21775 74440 21787 74443
rect 23311 74443 23369 74449
rect 23311 74440 23323 74443
rect 21775 74412 23323 74440
rect 21775 74409 21787 74412
rect 21729 74403 21787 74409
rect 23311 74409 23323 74412
rect 23357 74440 23369 74443
rect 35434 74440 35440 74452
rect 23357 74412 35440 74440
rect 23357 74409 23369 74412
rect 23311 74403 23369 74409
rect 35434 74400 35440 74412
rect 35492 74400 35498 74452
rect 74721 74443 74779 74449
rect 74721 74409 74733 74443
rect 74767 74440 74779 74443
rect 75086 74440 75092 74452
rect 74767 74412 75092 74440
rect 74767 74409 74779 74412
rect 74721 74403 74779 74409
rect 75086 74400 75092 74412
rect 75144 74440 75150 74452
rect 82538 74440 82544 74452
rect 75144 74412 82544 74440
rect 75144 74400 75150 74412
rect 82538 74400 82544 74412
rect 82596 74400 82602 74452
rect 85666 74400 85672 74452
rect 85724 74400 85730 74452
rect 85942 74400 85948 74452
rect 86000 74400 86006 74452
rect 87138 74400 87144 74452
rect 87196 74440 87202 74452
rect 87509 74443 87567 74449
rect 87509 74440 87521 74443
rect 87196 74412 87521 74440
rect 87196 74400 87202 74412
rect 87509 74409 87521 74412
rect 87555 74440 87567 74443
rect 88150 74440 88156 74452
rect 87555 74412 88156 74440
rect 87555 74409 87567 74412
rect 87509 74403 87567 74409
rect 88150 74400 88156 74412
rect 88208 74440 88214 74452
rect 91186 74440 91192 74452
rect 88208 74412 91192 74440
rect 88208 74400 88214 74412
rect 91186 74400 91192 74412
rect 91244 74400 91250 74452
rect 91557 74443 91615 74449
rect 91557 74409 91569 74443
rect 91603 74440 91615 74443
rect 93026 74440 93032 74452
rect 91603 74412 93032 74440
rect 91603 74409 91615 74412
rect 91557 74403 91615 74409
rect 93026 74400 93032 74412
rect 93084 74400 93090 74452
rect 96706 74400 96712 74452
rect 96764 74400 96770 74452
rect 98362 74400 98368 74452
rect 98420 74440 98426 74452
rect 99282 74440 99288 74452
rect 98420 74412 99288 74440
rect 98420 74400 98426 74412
rect 99282 74400 99288 74412
rect 99340 74440 99346 74452
rect 99929 74443 99987 74449
rect 99929 74440 99941 74443
rect 99340 74412 99941 74440
rect 99340 74400 99346 74412
rect 99929 74409 99941 74412
rect 99975 74409 99987 74443
rect 99929 74403 99987 74409
rect 101769 74443 101827 74449
rect 101769 74409 101781 74443
rect 101815 74440 101827 74443
rect 101950 74440 101956 74452
rect 101815 74412 101956 74440
rect 101815 74409 101827 74412
rect 101769 74403 101827 74409
rect 101950 74400 101956 74412
rect 102008 74400 102014 74452
rect 102873 74443 102931 74449
rect 102873 74409 102885 74443
rect 102919 74440 102931 74443
rect 103422 74440 103428 74452
rect 102919 74412 103428 74440
rect 102919 74409 102931 74412
rect 102873 74403 102931 74409
rect 103422 74400 103428 74412
rect 103480 74400 103486 74452
rect 842 74332 848 74384
rect 900 74372 906 74384
rect 1489 74375 1547 74381
rect 1489 74372 1501 74375
rect 900 74344 1501 74372
rect 900 74332 906 74344
rect 1489 74341 1501 74344
rect 1535 74341 1547 74375
rect 1489 74335 1547 74341
rect 84286 74332 84292 74384
rect 84344 74372 84350 74384
rect 90085 74375 90143 74381
rect 84344 74344 88472 74372
rect 84344 74332 84350 74344
rect 21821 74307 21879 74313
rect 21821 74273 21833 74307
rect 21867 74273 21879 74307
rect 28169 74307 28227 74313
rect 28169 74304 28181 74307
rect 21821 74267 21879 74273
rect 22204 74276 28181 74304
rect 1673 74239 1731 74245
rect 1673 74205 1685 74239
rect 1719 74236 1731 74239
rect 1857 74239 1915 74245
rect 1857 74236 1869 74239
rect 1719 74208 1869 74236
rect 1719 74205 1731 74208
rect 1673 74199 1731 74205
rect 1857 74205 1869 74208
rect 1903 74236 1915 74239
rect 21836 74236 21864 74267
rect 1903 74208 21864 74236
rect 22204 74222 22232 74276
rect 28169 74273 28181 74276
rect 28215 74273 28227 74307
rect 28169 74267 28227 74273
rect 88334 74264 88340 74316
rect 88392 74264 88398 74316
rect 88444 74304 88472 74344
rect 90085 74341 90097 74375
rect 90131 74372 90143 74375
rect 90269 74375 90327 74381
rect 90269 74372 90281 74375
rect 90131 74344 90281 74372
rect 90131 74341 90143 74344
rect 90085 74335 90143 74341
rect 90269 74341 90281 74344
rect 90315 74372 90327 74375
rect 98638 74372 98644 74384
rect 90315 74344 98644 74372
rect 90315 74341 90327 74344
rect 90269 74335 90327 74341
rect 98638 74332 98644 74344
rect 98696 74332 98702 74384
rect 100386 74332 100392 74384
rect 100444 74332 100450 74384
rect 101493 74375 101551 74381
rect 101493 74341 101505 74375
rect 101539 74372 101551 74375
rect 102042 74372 102048 74384
rect 101539 74344 102048 74372
rect 101539 74341 101551 74344
rect 101493 74335 101551 74341
rect 102042 74332 102048 74344
rect 102100 74332 102106 74384
rect 102134 74332 102140 74384
rect 102192 74372 102198 74384
rect 104158 74372 104164 74384
rect 102192 74344 104164 74372
rect 102192 74332 102198 74344
rect 104158 74332 104164 74344
rect 104216 74332 104222 74384
rect 104437 74375 104495 74381
rect 104437 74341 104449 74375
rect 104483 74372 104495 74375
rect 104526 74372 104532 74384
rect 104483 74344 104532 74372
rect 104483 74341 104495 74344
rect 104437 74335 104495 74341
rect 104526 74332 104532 74344
rect 104584 74332 104590 74384
rect 88613 74307 88671 74313
rect 88613 74304 88625 74307
rect 88444 74276 88625 74304
rect 88613 74273 88625 74276
rect 88659 74273 88671 74307
rect 88613 74267 88671 74273
rect 96798 74264 96804 74316
rect 96856 74304 96862 74316
rect 96893 74307 96951 74313
rect 96893 74304 96905 74307
rect 96856 74276 96905 74304
rect 96856 74264 96862 74276
rect 96893 74273 96905 74276
rect 96939 74273 96951 74307
rect 96893 74267 96951 74273
rect 97994 74264 98000 74316
rect 98052 74304 98058 74316
rect 99926 74304 99932 74316
rect 98052 74276 98132 74304
rect 98052 74264 98058 74276
rect 23569 74239 23627 74245
rect 1903 74205 1915 74208
rect 1857 74199 1915 74205
rect 21836 74100 21864 74208
rect 23569 74205 23581 74239
rect 23615 74236 23627 74239
rect 24581 74239 24639 74245
rect 23615 74208 23980 74236
rect 23615 74205 23627 74208
rect 23569 74199 23627 74205
rect 23382 74128 23388 74180
rect 23440 74168 23446 74180
rect 23952 74177 23980 74208
rect 24581 74205 24593 74239
rect 24627 74236 24639 74239
rect 24762 74236 24768 74248
rect 24627 74208 24768 74236
rect 24627 74205 24639 74208
rect 24581 74199 24639 74205
rect 24762 74196 24768 74208
rect 24820 74236 24826 74248
rect 28258 74236 28264 74248
rect 24820 74208 28264 74236
rect 24820 74196 24826 74208
rect 28258 74196 28264 74208
rect 28316 74236 28322 74248
rect 28445 74239 28503 74245
rect 28445 74236 28457 74239
rect 28316 74208 28457 74236
rect 28316 74196 28322 74208
rect 28445 74205 28457 74208
rect 28491 74236 28503 74239
rect 29733 74239 29791 74245
rect 29733 74236 29745 74239
rect 28491 74208 29745 74236
rect 28491 74205 28503 74208
rect 28445 74199 28503 74205
rect 29733 74205 29745 74208
rect 29779 74236 29791 74239
rect 29779 74208 29960 74236
rect 29779 74205 29791 74208
rect 29733 74199 29791 74205
rect 23937 74171 23995 74177
rect 23440 74140 23796 74168
rect 23440 74128 23446 74140
rect 23661 74103 23719 74109
rect 23661 74100 23673 74103
rect 21836 74072 23673 74100
rect 23661 74069 23673 74072
rect 23707 74069 23719 74103
rect 23768 74100 23796 74140
rect 23937 74137 23949 74171
rect 23983 74168 23995 74171
rect 25038 74168 25044 74180
rect 23983 74140 25044 74168
rect 23983 74137 23995 74140
rect 23937 74131 23995 74137
rect 25038 74128 25044 74140
rect 25096 74128 25102 74180
rect 24489 74103 24547 74109
rect 24489 74100 24501 74103
rect 23768 74072 24501 74100
rect 23661 74063 23719 74069
rect 24489 74069 24501 74072
rect 24535 74069 24547 74103
rect 24489 74063 24547 74069
rect 29638 74060 29644 74112
rect 29696 74060 29702 74112
rect 29932 74109 29960 74208
rect 74166 74196 74172 74248
rect 74224 74236 74230 74248
rect 74905 74239 74963 74245
rect 74905 74236 74917 74239
rect 74224 74208 74917 74236
rect 74224 74196 74230 74208
rect 74905 74205 74917 74208
rect 74951 74236 74963 74239
rect 78766 74236 78772 74248
rect 74951 74208 78772 74236
rect 74951 74205 74963 74208
rect 74905 74199 74963 74205
rect 78766 74196 78772 74208
rect 78824 74196 78830 74248
rect 85114 74196 85120 74248
rect 85172 74236 85178 74248
rect 85577 74239 85635 74245
rect 85577 74236 85589 74239
rect 85172 74208 85589 74236
rect 85172 74196 85178 74208
rect 85577 74205 85589 74208
rect 85623 74236 85635 74239
rect 85942 74236 85948 74248
rect 85623 74208 85948 74236
rect 85623 74205 85635 74208
rect 85577 74199 85635 74205
rect 85942 74196 85948 74208
rect 86000 74196 86006 74248
rect 87138 74196 87144 74248
rect 87196 74196 87202 74248
rect 91186 74196 91192 74248
rect 91244 74236 91250 74248
rect 91465 74239 91523 74245
rect 91465 74236 91477 74239
rect 91244 74208 91477 74236
rect 91244 74196 91250 74208
rect 91465 74205 91477 74208
rect 91511 74236 91523 74239
rect 91741 74239 91799 74245
rect 91741 74236 91753 74239
rect 91511 74208 91753 74236
rect 91511 74205 91523 74208
rect 91465 74199 91523 74205
rect 91741 74205 91753 74208
rect 91787 74205 91799 74239
rect 91741 74199 91799 74205
rect 96985 74239 97043 74245
rect 96985 74205 96997 74239
rect 97031 74236 97043 74239
rect 97442 74236 97448 74248
rect 97031 74208 97448 74236
rect 97031 74205 97043 74208
rect 96985 74199 97043 74205
rect 97442 74196 97448 74208
rect 97500 74196 97506 74248
rect 97902 74245 97908 74248
rect 97900 74236 97908 74245
rect 97863 74208 97908 74236
rect 97900 74199 97908 74208
rect 97902 74196 97908 74199
rect 97960 74196 97966 74248
rect 98104 74245 98132 74276
rect 98288 74276 99932 74304
rect 98288 74248 98316 74276
rect 99926 74264 99932 74276
rect 99984 74264 99990 74316
rect 100754 74304 100760 74316
rect 100128 74276 100760 74304
rect 98089 74239 98147 74245
rect 98089 74205 98101 74239
rect 98135 74205 98147 74239
rect 98270 74236 98276 74248
rect 98231 74208 98276 74236
rect 98089 74199 98147 74205
rect 98270 74196 98276 74208
rect 98328 74196 98334 74248
rect 98365 74239 98423 74245
rect 98365 74205 98377 74239
rect 98411 74236 98423 74239
rect 98638 74236 98644 74248
rect 98411 74208 98644 74236
rect 98411 74205 98423 74208
rect 98365 74199 98423 74205
rect 98638 74196 98644 74208
rect 98696 74196 98702 74248
rect 100128 74245 100156 74276
rect 100113 74239 100171 74245
rect 100113 74205 100125 74239
rect 100159 74205 100171 74239
rect 100113 74199 100171 74205
rect 100202 74196 100208 74248
rect 100260 74196 100266 74248
rect 100392 74245 100420 74276
rect 100754 74264 100760 74276
rect 100812 74264 100818 74316
rect 101858 74264 101864 74316
rect 101916 74304 101922 74316
rect 101953 74307 102011 74313
rect 101953 74304 101965 74307
rect 101916 74276 101965 74304
rect 101916 74264 101922 74276
rect 101953 74273 101965 74276
rect 101999 74273 102011 74307
rect 101953 74267 102011 74273
rect 102781 74307 102839 74313
rect 102781 74273 102793 74307
rect 102827 74304 102839 74307
rect 103054 74304 103060 74316
rect 102827 74276 103060 74304
rect 102827 74273 102839 74276
rect 102781 74267 102839 74273
rect 103054 74264 103060 74276
rect 103112 74264 103118 74316
rect 103514 74304 103520 74316
rect 103164 74276 103520 74304
rect 100377 74239 100435 74245
rect 100377 74205 100389 74239
rect 100423 74205 100435 74239
rect 100377 74199 100435 74205
rect 100570 74196 100576 74248
rect 100628 74196 100634 74248
rect 101306 74196 101312 74248
rect 101364 74196 101370 74248
rect 101674 74196 101680 74248
rect 101732 74236 101738 74248
rect 102045 74239 102103 74245
rect 102045 74236 102057 74239
rect 101732 74208 102057 74236
rect 101732 74196 101738 74208
rect 102045 74205 102057 74208
rect 102091 74205 102103 74239
rect 102045 74199 102103 74205
rect 102873 74239 102931 74245
rect 102873 74205 102885 74239
rect 102919 74236 102931 74239
rect 103164 74236 103192 74276
rect 103514 74264 103520 74276
rect 103572 74264 103578 74316
rect 105354 74264 105360 74316
rect 105412 74264 105418 74316
rect 105446 74264 105452 74316
rect 105504 74264 105510 74316
rect 102919 74208 103192 74236
rect 102919 74205 102931 74208
rect 102873 74199 102931 74205
rect 103238 74196 103244 74248
rect 103296 74196 103302 74248
rect 104434 74196 104440 74248
rect 104492 74196 104498 74248
rect 104713 74239 104771 74245
rect 104713 74205 104725 74239
rect 104759 74236 104771 74239
rect 104894 74236 104900 74248
rect 104759 74208 104900 74236
rect 104759 74205 104771 74208
rect 104713 74199 104771 74205
rect 104894 74196 104900 74208
rect 104952 74196 104958 74248
rect 105262 74196 105268 74248
rect 105320 74196 105326 74248
rect 108209 74239 108267 74245
rect 108209 74236 108221 74239
rect 108040 74208 108221 74236
rect 87233 74171 87291 74177
rect 87233 74137 87245 74171
rect 87279 74168 87291 74171
rect 97997 74171 98055 74177
rect 87279 74140 87736 74168
rect 87279 74137 87291 74140
rect 87233 74131 87291 74137
rect 29917 74103 29975 74109
rect 29917 74069 29929 74103
rect 29963 74100 29975 74103
rect 36170 74100 36176 74112
rect 29963 74072 36176 74100
rect 29963 74069 29975 74072
rect 29917 74063 29975 74069
rect 36170 74060 36176 74072
rect 36228 74060 36234 74112
rect 87708 74100 87736 74140
rect 88720 74140 89102 74168
rect 90008 74140 97856 74168
rect 88720 74100 88748 74140
rect 87708 74072 88748 74100
rect 88794 74060 88800 74112
rect 88852 74100 88858 74112
rect 90008 74100 90036 74140
rect 88852 74072 90036 74100
rect 90453 74103 90511 74109
rect 88852 74060 88858 74072
rect 90453 74069 90465 74103
rect 90499 74100 90511 74103
rect 91370 74100 91376 74112
rect 90499 74072 91376 74100
rect 90499 74069 90511 74072
rect 90453 74063 90511 74069
rect 91370 74060 91376 74072
rect 91428 74060 91434 74112
rect 97718 74060 97724 74112
rect 97776 74060 97782 74112
rect 97828 74100 97856 74140
rect 97997 74137 98009 74171
rect 98043 74168 98055 74171
rect 99190 74168 99196 74180
rect 98043 74140 99196 74168
rect 98043 74137 98055 74140
rect 97997 74131 98055 74137
rect 99190 74128 99196 74140
rect 99248 74128 99254 74180
rect 99742 74128 99748 74180
rect 99800 74168 99806 74180
rect 99800 74140 104296 74168
rect 99800 74128 99806 74140
rect 98914 74100 98920 74112
rect 97828 74072 98920 74100
rect 98914 74060 98920 74072
rect 98972 74060 98978 74112
rect 99926 74060 99932 74112
rect 99984 74100 99990 74112
rect 101582 74100 101588 74112
rect 99984 74072 101588 74100
rect 99984 74060 99990 74072
rect 101582 74060 101588 74072
rect 101640 74060 101646 74112
rect 101950 74060 101956 74112
rect 102008 74100 102014 74112
rect 102505 74103 102563 74109
rect 102505 74100 102517 74103
rect 102008 74072 102517 74100
rect 102008 74060 102014 74072
rect 102505 74069 102517 74072
rect 102551 74069 102563 74103
rect 102505 74063 102563 74069
rect 102870 74060 102876 74112
rect 102928 74100 102934 74112
rect 103057 74103 103115 74109
rect 103057 74100 103069 74103
rect 102928 74072 103069 74100
rect 102928 74060 102934 74072
rect 103057 74069 103069 74072
rect 103103 74069 103115 74103
rect 104268 74100 104296 74140
rect 104342 74128 104348 74180
rect 104400 74168 104406 74180
rect 108040 74177 108068 74208
rect 108209 74205 108221 74208
rect 108255 74205 108267 74239
rect 108209 74199 108267 74205
rect 104621 74171 104679 74177
rect 104621 74168 104633 74171
rect 104400 74140 104633 74168
rect 104400 74128 104406 74140
rect 104621 74137 104633 74140
rect 104667 74137 104679 74171
rect 108025 74171 108083 74177
rect 108025 74168 108037 74171
rect 104621 74131 104679 74137
rect 104820 74140 108037 74168
rect 104820 74100 104848 74140
rect 108025 74137 108037 74140
rect 108071 74137 108083 74171
rect 108025 74131 108083 74137
rect 104268 74072 104848 74100
rect 104897 74103 104955 74109
rect 103057 74063 103115 74069
rect 104897 74069 104909 74103
rect 104943 74100 104955 74103
rect 104986 74100 104992 74112
rect 104943 74072 104992 74100
rect 104943 74069 104955 74072
rect 104897 74063 104955 74069
rect 104986 74060 104992 74072
rect 105044 74060 105050 74112
rect 108390 74060 108396 74112
rect 108448 74060 108454 74112
rect 1104 74010 108836 74032
rect 1104 73958 4874 74010
rect 4926 73958 4938 74010
rect 4990 73958 5002 74010
rect 5054 73958 5066 74010
rect 5118 73958 5130 74010
rect 5182 73958 35594 74010
rect 35646 73958 35658 74010
rect 35710 73958 35722 74010
rect 35774 73958 35786 74010
rect 35838 73958 35850 74010
rect 35902 73958 66314 74010
rect 66366 73958 66378 74010
rect 66430 73958 66442 74010
rect 66494 73958 66506 74010
rect 66558 73958 66570 74010
rect 66622 73958 97034 74010
rect 97086 73958 97098 74010
rect 97150 73958 97162 74010
rect 97214 73958 97226 74010
rect 97278 73958 97290 74010
rect 97342 73958 108836 74010
rect 1104 73936 108836 73958
rect 9582 73856 9588 73908
rect 9640 73896 9646 73908
rect 35529 73899 35587 73905
rect 9640 73868 31754 73896
rect 9640 73856 9646 73868
rect 23382 73828 23388 73840
rect 18262 73800 23388 73828
rect 23382 73788 23388 73800
rect 23440 73788 23446 73840
rect 29638 73828 29644 73840
rect 24334 73800 29644 73828
rect 29638 73788 29644 73800
rect 29696 73788 29702 73840
rect 31726 73828 31754 73868
rect 35529 73865 35541 73899
rect 35575 73896 35587 73899
rect 39850 73896 39856 73908
rect 35575 73868 39856 73896
rect 35575 73865 35587 73868
rect 35529 73859 35587 73865
rect 39850 73856 39856 73868
rect 39908 73856 39914 73908
rect 68462 73856 68468 73908
rect 68520 73856 68526 73908
rect 68925 73899 68983 73905
rect 68925 73865 68937 73899
rect 68971 73865 68983 73899
rect 68925 73859 68983 73865
rect 68940 73828 68968 73859
rect 70118 73856 70124 73908
rect 70176 73856 70182 73908
rect 74445 73899 74503 73905
rect 74445 73865 74457 73899
rect 74491 73896 74503 73899
rect 74534 73896 74540 73908
rect 74491 73868 74540 73896
rect 74491 73865 74503 73868
rect 74445 73859 74503 73865
rect 74534 73856 74540 73868
rect 74592 73856 74598 73908
rect 75086 73896 75092 73908
rect 74828 73868 75092 73896
rect 74718 73828 74724 73840
rect 31726 73800 41414 73828
rect 68940 73800 74724 73828
rect 1673 73763 1731 73769
rect 1673 73729 1685 73763
rect 1719 73760 1731 73763
rect 11609 73763 11667 73769
rect 11609 73760 11621 73763
rect 1719 73732 1900 73760
rect 1719 73729 1731 73732
rect 1673 73723 1731 73729
rect 842 73584 848 73636
rect 900 73624 906 73636
rect 1489 73627 1547 73633
rect 1489 73624 1501 73627
rect 900 73596 1501 73624
rect 900 73584 906 73596
rect 1489 73593 1501 73596
rect 1535 73593 1547 73627
rect 1489 73587 1547 73593
rect 1872 73568 1900 73732
rect 11256 73732 11621 73760
rect 1854 73516 1860 73568
rect 1912 73516 1918 73568
rect 6178 73516 6184 73568
rect 6236 73556 6242 73568
rect 11256 73565 11284 73732
rect 11609 73729 11621 73732
rect 11655 73729 11667 73763
rect 11609 73723 11667 73729
rect 18966 73720 18972 73772
rect 19024 73720 19030 73772
rect 27985 73763 28043 73769
rect 27985 73729 27997 73763
rect 28031 73760 28043 73763
rect 28169 73763 28227 73769
rect 28169 73760 28181 73763
rect 28031 73732 28181 73760
rect 28031 73729 28043 73732
rect 27985 73723 28043 73729
rect 28169 73729 28181 73732
rect 28215 73760 28227 73763
rect 28258 73760 28264 73772
rect 28215 73732 28264 73760
rect 28215 73729 28227 73732
rect 28169 73723 28227 73729
rect 28258 73720 28264 73732
rect 28316 73720 28322 73772
rect 35437 73763 35495 73769
rect 35437 73729 35449 73763
rect 35483 73760 35495 73763
rect 38838 73760 38844 73772
rect 35483 73732 38844 73760
rect 35483 73729 35495 73732
rect 35437 73723 35495 73729
rect 38838 73720 38844 73732
rect 38896 73720 38902 73772
rect 41386 73760 41414 73800
rect 74718 73788 74724 73800
rect 74776 73788 74782 73840
rect 55217 73763 55275 73769
rect 55217 73760 55229 73763
rect 41386 73732 55229 73760
rect 55217 73729 55229 73732
rect 55263 73760 55275 73763
rect 55309 73763 55367 73769
rect 55309 73760 55321 73763
rect 55263 73732 55321 73760
rect 55263 73729 55275 73732
rect 55217 73723 55275 73729
rect 55309 73729 55321 73732
rect 55355 73729 55367 73763
rect 55309 73723 55367 73729
rect 68554 73720 68560 73772
rect 68612 73720 68618 73772
rect 69014 73720 69020 73772
rect 69072 73760 69078 73772
rect 70213 73763 70271 73769
rect 70213 73760 70225 73763
rect 69072 73732 70225 73760
rect 69072 73720 69078 73732
rect 70213 73729 70225 73732
rect 70259 73729 70271 73763
rect 70213 73723 70271 73729
rect 73801 73763 73859 73769
rect 73801 73729 73813 73763
rect 73847 73760 73859 73763
rect 74166 73760 74172 73772
rect 73847 73732 74172 73760
rect 73847 73729 73859 73732
rect 73801 73723 73859 73729
rect 74166 73720 74172 73732
rect 74224 73720 74230 73772
rect 74534 73720 74540 73772
rect 74592 73720 74598 73772
rect 11698 73652 11704 73704
rect 11756 73692 11762 73704
rect 13357 73695 13415 73701
rect 11756 73664 12434 73692
rect 11756 73652 11762 73664
rect 11241 73559 11299 73565
rect 11241 73556 11253 73559
rect 6236 73528 11253 73556
rect 6236 73516 6242 73528
rect 11241 73525 11253 73528
rect 11287 73525 11299 73559
rect 12406 73556 12434 73664
rect 13357 73661 13369 73695
rect 13403 73661 13415 73695
rect 13357 73655 13415 73661
rect 18693 73695 18751 73701
rect 18693 73661 18705 73695
rect 18739 73692 18751 73695
rect 24670 73692 24676 73704
rect 18739 73664 24676 73692
rect 18739 73661 18751 73664
rect 18693 73655 18751 73661
rect 13372 73624 13400 73655
rect 24670 73652 24676 73664
rect 24728 73652 24734 73704
rect 24762 73652 24768 73704
rect 24820 73652 24826 73704
rect 25038 73652 25044 73704
rect 25096 73692 25102 73704
rect 25409 73695 25467 73701
rect 25409 73692 25421 73695
rect 25096 73664 25421 73692
rect 25096 73652 25102 73664
rect 25409 73661 25421 73664
rect 25455 73692 25467 73695
rect 31754 73692 31760 73704
rect 25455 73664 31760 73692
rect 25455 73661 25467 73664
rect 25409 73655 25467 73661
rect 31754 73652 31760 73664
rect 31812 73652 31818 73704
rect 33042 73652 33048 73704
rect 33100 73692 33106 73704
rect 35621 73695 35679 73701
rect 35621 73692 35633 73695
rect 33100 73664 35633 73692
rect 33100 73652 33106 73664
rect 35621 73661 35633 73664
rect 35667 73692 35679 73695
rect 35897 73695 35955 73701
rect 35897 73692 35909 73695
rect 35667 73664 35909 73692
rect 35667 73661 35679 73664
rect 35621 73655 35679 73661
rect 35897 73661 35909 73664
rect 35943 73692 35955 73695
rect 37918 73692 37924 73704
rect 35943 73664 37924 73692
rect 35943 73661 35955 73664
rect 35897 73655 35955 73661
rect 37918 73652 37924 73664
rect 37976 73652 37982 73704
rect 68278 73652 68284 73704
rect 68336 73692 68342 73704
rect 69109 73695 69167 73701
rect 69109 73692 69121 73695
rect 68336 73664 69121 73692
rect 68336 73652 68342 73664
rect 69109 73661 69121 73664
rect 69155 73692 69167 73695
rect 69937 73695 69995 73701
rect 69937 73692 69949 73695
rect 69155 73664 69949 73692
rect 69155 73661 69167 73664
rect 69109 73655 69167 73661
rect 69937 73661 69949 73664
rect 69983 73692 69995 73695
rect 70673 73695 70731 73701
rect 70673 73692 70685 73695
rect 69983 73664 70685 73692
rect 69983 73661 69995 73664
rect 69937 73655 69995 73661
rect 70673 73661 70685 73664
rect 70719 73692 70731 73695
rect 72418 73692 72424 73704
rect 70719 73664 72424 73692
rect 70719 73661 70731 73664
rect 70673 73655 70731 73661
rect 72418 73652 72424 73664
rect 72476 73692 72482 73704
rect 73525 73695 73583 73701
rect 73525 73692 73537 73695
rect 72476 73664 73537 73692
rect 72476 73652 72482 73664
rect 73525 73661 73537 73664
rect 73571 73692 73583 73695
rect 73893 73695 73951 73701
rect 73893 73692 73905 73695
rect 73571 73664 73905 73692
rect 73571 73661 73583 73664
rect 73525 73655 73583 73661
rect 73893 73661 73905 73664
rect 73939 73661 73951 73695
rect 73893 73655 73951 73661
rect 74353 73695 74411 73701
rect 74353 73661 74365 73695
rect 74399 73692 74411 73695
rect 74828 73692 74856 73868
rect 75086 73856 75092 73868
rect 75144 73856 75150 73908
rect 84841 73899 84899 73905
rect 79336 73868 80054 73896
rect 74902 73788 74908 73840
rect 74960 73828 74966 73840
rect 79336 73828 79364 73868
rect 74960 73800 79364 73828
rect 80026 73828 80054 73868
rect 84841 73865 84853 73899
rect 84887 73896 84899 73899
rect 87417 73899 87475 73905
rect 84887 73868 86080 73896
rect 84887 73865 84899 73868
rect 84841 73859 84899 73865
rect 85945 73831 86003 73837
rect 85945 73828 85957 73831
rect 80026 73800 85957 73828
rect 74960 73788 74966 73800
rect 85945 73797 85957 73800
rect 85991 73797 86003 73831
rect 86052 73828 86080 73868
rect 87417 73865 87429 73899
rect 87463 73896 87475 73899
rect 87601 73899 87659 73905
rect 87601 73896 87613 73899
rect 87463 73868 87613 73896
rect 87463 73865 87475 73868
rect 87417 73859 87475 73865
rect 87601 73865 87613 73868
rect 87647 73896 87659 73899
rect 88702 73896 88708 73908
rect 87647 73868 88708 73896
rect 87647 73865 87659 73868
rect 87601 73859 87659 73865
rect 88702 73856 88708 73868
rect 88760 73856 88766 73908
rect 91370 73896 91376 73908
rect 88812 73868 91376 73896
rect 86052 73800 86434 73828
rect 85945 73791 86003 73797
rect 84286 73760 84292 73772
rect 74399 73664 74856 73692
rect 74920 73732 84292 73760
rect 74399 73661 74411 73664
rect 74353 73655 74411 73661
rect 13541 73627 13599 73633
rect 13541 73624 13553 73627
rect 13372 73596 13553 73624
rect 13541 73593 13553 73596
rect 13587 73624 13599 73627
rect 13814 73624 13820 73636
rect 13587 73596 13820 73624
rect 13587 73593 13599 73596
rect 13541 73587 13599 73593
rect 13814 73584 13820 73596
rect 13872 73624 13878 73636
rect 17129 73627 17187 73633
rect 17129 73624 17141 73627
rect 13872 73596 17141 73624
rect 13872 73584 13878 73596
rect 17129 73593 17141 73596
rect 17175 73624 17187 73627
rect 73154 73624 73160 73636
rect 17175 73596 17356 73624
rect 17175 73593 17187 73596
rect 17129 73587 17187 73593
rect 17221 73559 17279 73565
rect 17221 73556 17233 73559
rect 12406 73528 17233 73556
rect 11241 73519 11299 73525
rect 17221 73525 17233 73528
rect 17267 73525 17279 73559
rect 17328 73556 17356 73596
rect 64846 73596 73160 73624
rect 18966 73556 18972 73568
rect 17328 73528 18972 73556
rect 17221 73519 17279 73525
rect 18966 73516 18972 73528
rect 19024 73516 19030 73568
rect 22922 73516 22928 73568
rect 22980 73556 22986 73568
rect 23293 73559 23351 73565
rect 23293 73556 23305 73559
rect 22980 73528 23305 73556
rect 22980 73516 22986 73528
rect 23293 73525 23305 73528
rect 23339 73556 23351 73559
rect 25133 73559 25191 73565
rect 25133 73556 25145 73559
rect 23339 73528 25145 73556
rect 23339 73525 23351 73528
rect 23293 73519 23351 73525
rect 25133 73525 25145 73528
rect 25179 73525 25191 73559
rect 25133 73519 25191 73525
rect 27890 73516 27896 73568
rect 27948 73516 27954 73568
rect 29362 73516 29368 73568
rect 29420 73556 29426 73568
rect 35069 73559 35127 73565
rect 35069 73556 35081 73559
rect 29420 73528 35081 73556
rect 29420 73516 29426 73528
rect 35069 73525 35081 73528
rect 35115 73525 35127 73559
rect 35069 73519 35127 73525
rect 56134 73516 56140 73568
rect 56192 73556 56198 73568
rect 56781 73559 56839 73565
rect 56781 73556 56793 73559
rect 56192 73528 56793 73556
rect 56192 73516 56198 73528
rect 56781 73525 56793 73528
rect 56827 73556 56839 73559
rect 57241 73559 57299 73565
rect 57241 73556 57253 73559
rect 56827 73528 57253 73556
rect 56827 73525 56839 73528
rect 56781 73519 56839 73525
rect 57241 73525 57253 73528
rect 57287 73556 57299 73559
rect 64846 73556 64874 73596
rect 73154 73584 73160 73596
rect 73212 73624 73218 73636
rect 73798 73624 73804 73636
rect 73212 73596 73804 73624
rect 73212 73584 73218 73596
rect 73798 73584 73804 73596
rect 73856 73584 73862 73636
rect 74920 73633 74948 73732
rect 84286 73720 84292 73732
rect 84344 73720 84350 73772
rect 84933 73763 84991 73769
rect 84933 73729 84945 73763
rect 84979 73760 84991 73763
rect 85114 73760 85120 73772
rect 84979 73732 85120 73760
rect 84979 73729 84991 73732
rect 84933 73723 84991 73729
rect 85114 73720 85120 73732
rect 85172 73720 85178 73772
rect 88812 73769 88840 73868
rect 91370 73856 91376 73868
rect 91428 73856 91434 73908
rect 93302 73856 93308 73908
rect 93360 73856 93366 73908
rect 98178 73896 98184 73908
rect 93688 73868 98184 73896
rect 89530 73788 89536 73840
rect 89588 73788 89594 73840
rect 90805 73831 90863 73837
rect 90805 73797 90817 73831
rect 90851 73828 90863 73831
rect 90851 73800 90956 73828
rect 90851 73797 90863 73800
rect 90805 73791 90863 73797
rect 88797 73763 88855 73769
rect 88797 73729 88809 73763
rect 88843 73729 88855 73763
rect 90928 73760 90956 73800
rect 91002 73788 91008 73840
rect 91060 73788 91066 73840
rect 91189 73831 91247 73837
rect 91189 73797 91201 73831
rect 91235 73828 91247 73831
rect 93688 73828 93716 73868
rect 98178 73856 98184 73868
rect 98236 73856 98242 73908
rect 98822 73856 98828 73908
rect 98880 73856 98886 73908
rect 98914 73856 98920 73908
rect 98972 73896 98978 73908
rect 99742 73896 99748 73908
rect 98972 73868 99748 73896
rect 98972 73856 98978 73868
rect 99742 73856 99748 73868
rect 99800 73856 99806 73908
rect 99926 73856 99932 73908
rect 99984 73896 99990 73908
rect 100294 73896 100300 73908
rect 99984 73868 100300 73896
rect 99984 73856 99990 73868
rect 100294 73856 100300 73868
rect 100352 73856 100358 73908
rect 101953 73899 102011 73905
rect 101953 73896 101965 73899
rect 101416 73868 101965 73896
rect 91235 73800 93716 73828
rect 91235 73797 91247 73800
rect 91189 73791 91247 73797
rect 91278 73760 91284 73772
rect 90928 73732 91284 73760
rect 88797 73723 88855 73729
rect 91278 73720 91284 73732
rect 91336 73720 91342 73772
rect 78582 73652 78588 73704
rect 78640 73692 78646 73704
rect 85574 73692 85580 73704
rect 78640 73664 85580 73692
rect 78640 73652 78646 73664
rect 85574 73652 85580 73664
rect 85632 73652 85638 73704
rect 85669 73695 85727 73701
rect 85669 73661 85681 73695
rect 85715 73661 85727 73695
rect 85669 73655 85727 73661
rect 74905 73627 74963 73633
rect 74905 73593 74917 73627
rect 74951 73593 74963 73627
rect 74905 73587 74963 73593
rect 57287 73528 64874 73556
rect 57287 73525 57299 73528
rect 57241 73519 57299 73525
rect 70578 73516 70584 73568
rect 70636 73516 70642 73568
rect 85577 73559 85635 73565
rect 85577 73525 85589 73559
rect 85623 73556 85635 73559
rect 85684 73556 85712 73655
rect 89070 73652 89076 73704
rect 89128 73652 89134 73704
rect 90545 73695 90603 73701
rect 90545 73661 90557 73695
rect 90591 73692 90603 73695
rect 91388 73692 91416 73800
rect 97810 73788 97816 73840
rect 97868 73828 97874 73840
rect 98270 73828 98276 73840
rect 97868 73800 98276 73828
rect 97868 73788 97874 73800
rect 98270 73788 98276 73800
rect 98328 73788 98334 73840
rect 99116 73800 100156 73828
rect 93302 73720 93308 73772
rect 93360 73760 93366 73772
rect 93489 73763 93547 73769
rect 93489 73760 93501 73763
rect 93360 73732 93501 73760
rect 93360 73720 93366 73732
rect 93489 73729 93501 73732
rect 93535 73729 93547 73763
rect 93489 73723 93547 73729
rect 93673 73763 93731 73769
rect 93673 73729 93685 73763
rect 93719 73729 93731 73763
rect 93673 73723 93731 73729
rect 90591 73664 91416 73692
rect 90591 73661 90603 73664
rect 90545 73655 90603 73661
rect 90637 73627 90695 73633
rect 90637 73624 90649 73627
rect 90192 73596 90649 73624
rect 86034 73556 86040 73568
rect 85623 73528 86040 73556
rect 85623 73525 85635 73528
rect 85577 73519 85635 73525
rect 86034 73516 86040 73528
rect 86092 73516 86098 73568
rect 89622 73516 89628 73568
rect 89680 73556 89686 73568
rect 90192 73556 90220 73596
rect 90637 73593 90649 73596
rect 90683 73593 90695 73627
rect 91462 73624 91468 73636
rect 90637 73587 90695 73593
rect 90836 73596 91468 73624
rect 90836 73565 90864 73596
rect 91462 73584 91468 73596
rect 91520 73584 91526 73636
rect 93504 73624 93532 73723
rect 93688 73692 93716 73723
rect 93854 73720 93860 73772
rect 93912 73760 93918 73772
rect 94133 73763 94191 73769
rect 94133 73760 94145 73763
rect 93912 73732 94145 73760
rect 93912 73720 93918 73732
rect 94133 73729 94145 73732
rect 94179 73729 94191 73763
rect 94133 73723 94191 73729
rect 94406 73720 94412 73772
rect 94464 73720 94470 73772
rect 94593 73763 94651 73769
rect 94593 73729 94605 73763
rect 94639 73729 94651 73763
rect 94593 73723 94651 73729
rect 94424 73692 94452 73720
rect 93688 73664 94452 73692
rect 94608 73624 94636 73723
rect 97442 73720 97448 73772
rect 97500 73760 97506 73772
rect 98454 73760 98460 73772
rect 97500 73732 98460 73760
rect 97500 73720 97506 73732
rect 98454 73720 98460 73732
rect 98512 73760 98518 73772
rect 98641 73763 98699 73769
rect 98641 73760 98653 73763
rect 98512 73732 98653 73760
rect 98512 73720 98518 73732
rect 98641 73729 98653 73732
rect 98687 73729 98699 73763
rect 98641 73723 98699 73729
rect 98917 73763 98975 73769
rect 98917 73729 98929 73763
rect 98963 73760 98975 73763
rect 99006 73760 99012 73772
rect 98963 73732 99012 73760
rect 98963 73729 98975 73732
rect 98917 73723 98975 73729
rect 99006 73720 99012 73732
rect 99064 73720 99070 73772
rect 99116 73769 99144 73800
rect 99101 73763 99159 73769
rect 99101 73729 99113 73763
rect 99147 73729 99159 73763
rect 99101 73723 99159 73729
rect 98362 73652 98368 73704
rect 98420 73692 98426 73704
rect 99116 73692 99144 73723
rect 99282 73720 99288 73772
rect 99340 73720 99346 73772
rect 99374 73720 99380 73772
rect 99432 73760 99438 73772
rect 100021 73763 100079 73769
rect 100021 73760 100033 73763
rect 99432 73732 100033 73760
rect 99432 73720 99438 73732
rect 100021 73729 100033 73732
rect 100067 73729 100079 73763
rect 100128 73766 100156 73800
rect 100570 73788 100576 73840
rect 100628 73828 100634 73840
rect 101122 73828 101128 73840
rect 100628 73800 101128 73828
rect 100628 73788 100634 73800
rect 101122 73788 101128 73800
rect 101180 73828 101186 73840
rect 101416 73828 101444 73868
rect 101953 73865 101965 73868
rect 101999 73896 102011 73899
rect 102134 73896 102140 73908
rect 101999 73868 102140 73896
rect 101999 73865 102011 73868
rect 101953 73859 102011 73865
rect 102134 73856 102140 73868
rect 102192 73856 102198 73908
rect 103422 73856 103428 73908
rect 103480 73896 103486 73908
rect 104434 73896 104440 73908
rect 103480 73868 104440 73896
rect 103480 73856 103486 73868
rect 104434 73856 104440 73868
rect 104492 73896 104498 73908
rect 104897 73899 104955 73905
rect 104897 73896 104909 73899
rect 104492 73868 104909 73896
rect 104492 73856 104498 73868
rect 104897 73865 104909 73868
rect 104943 73865 104955 73899
rect 104897 73859 104955 73865
rect 105265 73899 105323 73905
rect 105265 73865 105277 73899
rect 105311 73896 105323 73899
rect 105446 73896 105452 73908
rect 105311 73868 105452 73896
rect 105311 73865 105323 73868
rect 105265 73859 105323 73865
rect 105446 73856 105452 73868
rect 105504 73856 105510 73908
rect 105906 73896 105912 73908
rect 105648 73868 105912 73896
rect 101180 73800 101444 73828
rect 101180 73788 101186 73800
rect 101582 73788 101588 73840
rect 101640 73828 101646 73840
rect 102505 73831 102563 73837
rect 102505 73828 102517 73831
rect 101640 73800 102517 73828
rect 101640 73788 101646 73800
rect 102505 73797 102517 73800
rect 102551 73828 102563 73831
rect 102870 73828 102876 73840
rect 102551 73800 102876 73828
rect 102551 73797 102563 73800
rect 102505 73791 102563 73797
rect 102870 73788 102876 73800
rect 102928 73788 102934 73840
rect 103514 73828 103520 73840
rect 103164 73800 103520 73828
rect 100128 73760 100340 73766
rect 100478 73760 100484 73772
rect 100128 73738 100484 73760
rect 100312 73732 100484 73738
rect 100021 73723 100079 73729
rect 100478 73720 100484 73732
rect 100536 73720 100542 73772
rect 100665 73763 100723 73769
rect 100665 73729 100677 73763
rect 100711 73760 100723 73763
rect 100754 73760 100760 73772
rect 100711 73732 100760 73760
rect 100711 73729 100723 73732
rect 100665 73723 100723 73729
rect 100754 73720 100760 73732
rect 100812 73720 100818 73772
rect 101766 73720 101772 73772
rect 101824 73760 101830 73772
rect 101861 73763 101919 73769
rect 101861 73760 101873 73763
rect 101824 73732 101873 73760
rect 101824 73720 101830 73732
rect 101861 73729 101873 73732
rect 101907 73729 101919 73763
rect 102321 73763 102379 73769
rect 102321 73760 102333 73763
rect 101861 73723 101919 73729
rect 101968 73732 102333 73760
rect 99561 73695 99619 73701
rect 99561 73692 99573 73695
rect 98420 73664 99144 73692
rect 99208 73664 99573 73692
rect 98420 73652 98426 73664
rect 93504 73596 94636 73624
rect 98638 73584 98644 73636
rect 98696 73584 98702 73636
rect 98730 73584 98736 73636
rect 98788 73624 98794 73636
rect 99208 73624 99236 73664
rect 99561 73661 99573 73664
rect 99607 73661 99619 73695
rect 99561 73655 99619 73661
rect 99650 73652 99656 73704
rect 99708 73692 99714 73704
rect 99837 73695 99895 73701
rect 99837 73692 99849 73695
rect 99708 73664 99849 73692
rect 99708 73652 99714 73664
rect 99837 73661 99849 73664
rect 99883 73661 99895 73695
rect 99837 73655 99895 73661
rect 100205 73695 100263 73701
rect 100205 73661 100217 73695
rect 100251 73661 100263 73695
rect 100205 73655 100263 73661
rect 98788 73596 99236 73624
rect 98788 73584 98794 73596
rect 99466 73584 99472 73636
rect 99524 73584 99530 73636
rect 100220 73624 100248 73655
rect 100294 73652 100300 73704
rect 100352 73652 100358 73704
rect 100386 73652 100392 73704
rect 100444 73652 100450 73704
rect 101306 73624 101312 73636
rect 100220 73596 101312 73624
rect 101306 73584 101312 73596
rect 101364 73584 101370 73636
rect 89680 73528 90220 73556
rect 90821 73559 90879 73565
rect 89680 73516 89686 73528
rect 90821 73525 90833 73559
rect 90867 73525 90879 73559
rect 90821 73519 90879 73525
rect 91370 73516 91376 73568
rect 91428 73556 91434 73568
rect 91830 73556 91836 73568
rect 91428 73528 91836 73556
rect 91428 73516 91434 73528
rect 91830 73516 91836 73528
rect 91888 73516 91894 73568
rect 93578 73516 93584 73568
rect 93636 73516 93642 73568
rect 93946 73516 93952 73568
rect 94004 73516 94010 73568
rect 99377 73559 99435 73565
rect 99377 73525 99389 73559
rect 99423 73556 99435 73559
rect 100110 73556 100116 73568
rect 99423 73528 100116 73556
rect 99423 73525 99435 73528
rect 99377 73519 99435 73525
rect 100110 73516 100116 73528
rect 100168 73516 100174 73568
rect 100294 73516 100300 73568
rect 100352 73556 100358 73568
rect 101968 73556 101996 73732
rect 102321 73729 102333 73732
rect 102367 73760 102379 73763
rect 102778 73760 102784 73772
rect 102367 73732 102784 73760
rect 102367 73729 102379 73732
rect 102321 73723 102379 73729
rect 102778 73720 102784 73732
rect 102836 73720 102842 73772
rect 102965 73763 103023 73769
rect 102965 73729 102977 73763
rect 103011 73760 103023 73763
rect 103054 73760 103060 73772
rect 103011 73732 103060 73760
rect 103011 73729 103023 73732
rect 102965 73723 103023 73729
rect 103054 73720 103060 73732
rect 103112 73720 103118 73772
rect 103164 73769 103192 73800
rect 103514 73788 103520 73800
rect 103572 73788 103578 73840
rect 104618 73788 104624 73840
rect 104676 73788 104682 73840
rect 105648 73837 105676 73868
rect 105906 73856 105912 73868
rect 105964 73896 105970 73908
rect 108301 73899 108359 73905
rect 108301 73896 108313 73899
rect 105964 73868 108313 73896
rect 105964 73856 105970 73868
rect 108301 73865 108313 73868
rect 108347 73865 108359 73899
rect 108301 73859 108359 73865
rect 105633 73831 105691 73837
rect 105633 73797 105645 73831
rect 105679 73797 105691 73831
rect 105633 73791 105691 73797
rect 103149 73763 103207 73769
rect 103149 73729 103161 73763
rect 103195 73729 103207 73763
rect 103149 73723 103207 73729
rect 103422 73720 103428 73772
rect 103480 73720 103486 73772
rect 104253 73763 104311 73769
rect 104253 73729 104265 73763
rect 104299 73729 104311 73763
rect 104253 73723 104311 73729
rect 104346 73763 104404 73769
rect 104346 73729 104358 73763
rect 104392 73729 104404 73763
rect 104346 73723 104404 73729
rect 104529 73763 104587 73769
rect 104529 73729 104541 73763
rect 104575 73760 104587 73763
rect 104575 73732 104648 73760
rect 104575 73729 104587 73732
rect 104529 73723 104587 73729
rect 102689 73695 102747 73701
rect 102689 73661 102701 73695
rect 102735 73692 102747 73695
rect 103606 73692 103612 73704
rect 102735 73664 103612 73692
rect 102735 73661 102747 73664
rect 102689 73655 102747 73661
rect 103606 73652 103612 73664
rect 103664 73692 103670 73704
rect 104268 73692 104296 73723
rect 103664 73664 104296 73692
rect 103664 73652 103670 73664
rect 103790 73584 103796 73636
rect 103848 73624 103854 73636
rect 104360 73624 104388 73723
rect 104620 73636 104648 73732
rect 104710 73720 104716 73772
rect 104768 73769 104774 73772
rect 104768 73760 104776 73769
rect 104768 73732 104813 73760
rect 104768 73723 104776 73732
rect 104768 73720 104774 73723
rect 105170 73720 105176 73772
rect 105228 73720 105234 73772
rect 105354 73720 105360 73772
rect 105412 73720 105418 73772
rect 105538 73720 105544 73772
rect 105596 73760 105602 73772
rect 105817 73763 105875 73769
rect 105817 73760 105829 73763
rect 105596 73732 105829 73760
rect 105596 73720 105602 73732
rect 105817 73729 105829 73732
rect 105863 73729 105875 73763
rect 105817 73723 105875 73729
rect 108209 73763 108267 73769
rect 108209 73729 108221 73763
rect 108255 73760 108267 73763
rect 108482 73760 108488 73772
rect 108255 73732 108488 73760
rect 108255 73729 108267 73732
rect 108209 73723 108267 73729
rect 108482 73720 108488 73732
rect 108540 73720 108546 73772
rect 104894 73652 104900 73704
rect 104952 73692 104958 73704
rect 105449 73695 105507 73701
rect 105449 73692 105461 73695
rect 104952 73664 105461 73692
rect 104952 73652 104958 73664
rect 105449 73661 105461 73664
rect 105495 73661 105507 73695
rect 105449 73655 105507 73661
rect 103848 73596 104388 73624
rect 103848 73584 103854 73596
rect 104618 73584 104624 73636
rect 104676 73624 104682 73636
rect 105262 73624 105268 73636
rect 104676 73596 105268 73624
rect 104676 73584 104682 73596
rect 105262 73584 105268 73596
rect 105320 73584 105326 73636
rect 100352 73528 101996 73556
rect 100352 73516 100358 73528
rect 103514 73516 103520 73568
rect 103572 73556 103578 73568
rect 103609 73559 103667 73565
rect 103609 73556 103621 73559
rect 103572 73528 103621 73556
rect 103572 73516 103578 73528
rect 103609 73525 103621 73528
rect 103655 73525 103667 73559
rect 103609 73519 103667 73525
rect 1104 73466 108836 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 34934 73466
rect 34986 73414 34998 73466
rect 35050 73414 35062 73466
rect 35114 73414 35126 73466
rect 35178 73414 35190 73466
rect 35242 73414 65654 73466
rect 65706 73414 65718 73466
rect 65770 73414 65782 73466
rect 65834 73414 65846 73466
rect 65898 73414 65910 73466
rect 65962 73414 96374 73466
rect 96426 73414 96438 73466
rect 96490 73414 96502 73466
rect 96554 73414 96566 73466
rect 96618 73414 96630 73466
rect 96682 73414 108836 73466
rect 1104 73392 108836 73414
rect 1854 73312 1860 73364
rect 1912 73352 1918 73364
rect 21453 73355 21511 73361
rect 21453 73352 21465 73355
rect 1912 73324 21465 73352
rect 1912 73312 1918 73324
rect 21453 73321 21465 73324
rect 21499 73352 21511 73355
rect 23293 73355 23351 73361
rect 23293 73352 23305 73355
rect 21499 73324 23305 73352
rect 21499 73321 21511 73324
rect 21453 73315 21511 73321
rect 23293 73321 23305 73324
rect 23339 73321 23351 73355
rect 23293 73315 23351 73321
rect 23569 73355 23627 73361
rect 23569 73321 23581 73355
rect 23615 73352 23627 73355
rect 25038 73352 25044 73364
rect 23615 73324 25044 73352
rect 23615 73321 23627 73324
rect 23569 73315 23627 73321
rect 1857 73219 1915 73225
rect 1857 73185 1869 73219
rect 1903 73216 1915 73219
rect 22922 73216 22928 73228
rect 1903 73188 22928 73216
rect 1903 73185 1915 73188
rect 1857 73179 1915 73185
rect 1673 73151 1731 73157
rect 1673 73117 1685 73151
rect 1719 73148 1731 73151
rect 1872 73148 1900 73179
rect 22922 73176 22928 73188
rect 22980 73176 22986 73228
rect 23201 73219 23259 73225
rect 23201 73185 23213 73219
rect 23247 73216 23259 73219
rect 23584 73216 23612 73315
rect 25038 73312 25044 73324
rect 25096 73312 25102 73364
rect 70578 73312 70584 73364
rect 70636 73352 70642 73364
rect 78582 73352 78588 73364
rect 70636 73324 78588 73352
rect 70636 73312 70642 73324
rect 78582 73312 78588 73324
rect 78640 73312 78646 73364
rect 78692 73324 80192 73352
rect 69106 73244 69112 73296
rect 69164 73284 69170 73296
rect 70489 73287 70547 73293
rect 70489 73284 70501 73287
rect 69164 73256 70501 73284
rect 69164 73244 69170 73256
rect 70489 73253 70501 73256
rect 70535 73284 70547 73287
rect 70535 73256 72924 73284
rect 70535 73253 70547 73256
rect 70489 73247 70547 73253
rect 72896 73228 72924 73256
rect 29362 73216 29368 73228
rect 23247 73188 23612 73216
rect 23676 73188 29368 73216
rect 23247 73185 23259 73188
rect 23201 73179 23259 73185
rect 1719 73120 1900 73148
rect 1719 73117 1731 73120
rect 1673 73111 1731 73117
rect 22925 73083 22983 73089
rect 22494 73052 22876 73080
rect 842 72972 848 73024
rect 900 73012 906 73024
rect 1489 73015 1547 73021
rect 1489 73012 1501 73015
rect 900 72984 1501 73012
rect 900 72972 906 72984
rect 1489 72981 1501 72984
rect 1535 72981 1547 73015
rect 22848 73012 22876 73052
rect 22925 73049 22937 73083
rect 22971 73080 22983 73083
rect 23676 73080 23704 73188
rect 29362 73176 29368 73188
rect 29420 73176 29426 73228
rect 37918 73176 37924 73228
rect 37976 73216 37982 73228
rect 38197 73219 38255 73225
rect 38197 73216 38209 73219
rect 37976 73188 38209 73216
rect 37976 73176 37982 73188
rect 38197 73185 38209 73188
rect 38243 73216 38255 73219
rect 40405 73219 40463 73225
rect 40405 73216 40417 73219
rect 38243 73188 40417 73216
rect 38243 73185 38255 73188
rect 38197 73179 38255 73185
rect 40405 73185 40417 73188
rect 40451 73216 40463 73219
rect 40681 73219 40739 73225
rect 40681 73216 40693 73219
rect 40451 73188 40693 73216
rect 40451 73185 40463 73188
rect 40405 73179 40463 73185
rect 40681 73185 40693 73188
rect 40727 73216 40739 73219
rect 68278 73216 68284 73228
rect 40727 73188 68284 73216
rect 40727 73185 40739 73188
rect 40681 73179 40739 73185
rect 68278 73176 68284 73188
rect 68336 73176 68342 73228
rect 72418 73176 72424 73228
rect 72476 73216 72482 73228
rect 72476 73188 72832 73216
rect 72476 73176 72482 73188
rect 24762 73108 24768 73160
rect 24820 73148 24826 73160
rect 40313 73151 40371 73157
rect 24820 73120 39896 73148
rect 24820 73108 24826 73120
rect 22971 73052 23704 73080
rect 22971 73049 22983 73052
rect 22925 73043 22983 73049
rect 27890 73012 27896 73024
rect 22848 72984 27896 73012
rect 1489 72975 1547 72981
rect 27890 72972 27896 72984
rect 27948 72972 27954 73024
rect 35434 72972 35440 73024
rect 35492 73012 35498 73024
rect 37369 73015 37427 73021
rect 37369 73012 37381 73015
rect 35492 72984 37381 73012
rect 35492 72972 35498 72984
rect 37369 72981 37381 72984
rect 37415 72981 37427 73015
rect 37369 72975 37427 72981
rect 37734 72972 37740 73024
rect 37792 72972 37798 73024
rect 37826 72972 37832 73024
rect 37884 72972 37890 73024
rect 39868 73021 39896 73120
rect 40313 73117 40325 73151
rect 40359 73148 40371 73151
rect 45462 73148 45468 73160
rect 40359 73120 45468 73148
rect 40359 73117 40371 73120
rect 40313 73111 40371 73117
rect 45462 73108 45468 73120
rect 45520 73108 45526 73160
rect 68922 73108 68928 73160
rect 68980 73148 68986 73160
rect 72605 73151 72663 73157
rect 72605 73148 72617 73151
rect 68980 73120 72617 73148
rect 68980 73108 68986 73120
rect 72605 73117 72617 73120
rect 72651 73117 72663 73151
rect 72804 73148 72832 73188
rect 72878 73176 72884 73228
rect 72936 73216 72942 73228
rect 78692 73225 78720 73324
rect 78766 73244 78772 73296
rect 78824 73244 78830 73296
rect 80164 73225 80192 73324
rect 88150 73312 88156 73364
rect 88208 73312 88214 73364
rect 93302 73312 93308 73364
rect 93360 73352 93366 73364
rect 93765 73355 93823 73361
rect 93765 73352 93777 73355
rect 93360 73324 93777 73352
rect 93360 73312 93366 73324
rect 93765 73321 93777 73324
rect 93811 73321 93823 73355
rect 93765 73315 93823 73321
rect 98546 73312 98552 73364
rect 98604 73312 98610 73364
rect 98733 73355 98791 73361
rect 98733 73321 98745 73355
rect 98779 73352 98791 73355
rect 99282 73352 99288 73364
rect 98779 73324 99288 73352
rect 98779 73321 98791 73324
rect 98733 73315 98791 73321
rect 99282 73312 99288 73324
rect 99340 73312 99346 73364
rect 99558 73312 99564 73364
rect 99616 73352 99622 73364
rect 100294 73352 100300 73364
rect 99616 73324 100300 73352
rect 99616 73312 99622 73324
rect 100294 73312 100300 73324
rect 100352 73312 100358 73364
rect 100386 73312 100392 73364
rect 100444 73352 100450 73364
rect 100573 73355 100631 73361
rect 100573 73352 100585 73355
rect 100444 73324 100585 73352
rect 100444 73312 100450 73324
rect 100573 73321 100585 73324
rect 100619 73321 100631 73355
rect 100573 73315 100631 73321
rect 100757 73355 100815 73361
rect 100757 73321 100769 73355
rect 100803 73321 100815 73355
rect 100757 73315 100815 73321
rect 101677 73355 101735 73361
rect 101677 73321 101689 73355
rect 101723 73352 101735 73355
rect 101858 73352 101864 73364
rect 101723 73324 101864 73352
rect 101723 73321 101735 73324
rect 101677 73315 101735 73321
rect 78677 73219 78735 73225
rect 78677 73216 78689 73219
rect 72936 73188 78689 73216
rect 72936 73176 72942 73188
rect 78677 73185 78689 73188
rect 78723 73185 78735 73219
rect 78677 73179 78735 73185
rect 80149 73219 80207 73225
rect 80149 73185 80161 73219
rect 80195 73185 80207 73219
rect 88168 73216 88196 73312
rect 97718 73284 97724 73296
rect 97092 73256 97724 73284
rect 80149 73179 80207 73185
rect 87800 73188 88196 73216
rect 87800 73157 87828 73188
rect 93854 73176 93860 73228
rect 93912 73216 93918 73228
rect 95513 73219 95571 73225
rect 95513 73216 95525 73219
rect 93912 73188 95525 73216
rect 93912 73176 93918 73188
rect 95513 73185 95525 73188
rect 95559 73185 95571 73219
rect 95513 73179 95571 73185
rect 95881 73219 95939 73225
rect 95881 73185 95893 73219
rect 95927 73216 95939 73219
rect 97092 73216 97120 73256
rect 97718 73244 97724 73256
rect 97776 73244 97782 73296
rect 98454 73244 98460 73296
rect 98512 73284 98518 73296
rect 100110 73284 100116 73296
rect 98512 73256 100116 73284
rect 98512 73244 98518 73256
rect 100110 73244 100116 73256
rect 100168 73244 100174 73296
rect 100772 73284 100800 73315
rect 101858 73312 101864 73324
rect 101916 73312 101922 73364
rect 102965 73355 103023 73361
rect 102965 73321 102977 73355
rect 103011 73321 103023 73355
rect 102965 73315 103023 73321
rect 101582 73284 101588 73296
rect 100312 73256 101588 73284
rect 95927 73188 97120 73216
rect 95927 73185 95939 73188
rect 95881 73179 95939 73185
rect 73157 73151 73215 73157
rect 73157 73148 73169 73151
rect 72804 73120 73169 73148
rect 72605 73111 72663 73117
rect 73157 73117 73169 73120
rect 73203 73117 73215 73151
rect 73157 73111 73215 73117
rect 87785 73151 87843 73157
rect 87785 73117 87797 73151
rect 87831 73117 87843 73151
rect 87785 73111 87843 73117
rect 87877 73151 87935 73157
rect 87877 73117 87889 73151
rect 87923 73148 87935 73151
rect 89530 73148 89536 73160
rect 87923 73120 89536 73148
rect 87923 73117 87935 73120
rect 87877 73111 87935 73117
rect 89530 73108 89536 73120
rect 89588 73108 89594 73160
rect 95697 73151 95755 73157
rect 95697 73117 95709 73151
rect 95743 73148 95755 73151
rect 96890 73148 96896 73160
rect 95743 73120 96896 73148
rect 95743 73117 95755 73120
rect 95697 73111 95755 73117
rect 96890 73108 96896 73120
rect 96948 73148 96954 73160
rect 97092 73157 97120 73188
rect 97353 73219 97411 73225
rect 97353 73185 97365 73219
rect 97399 73216 97411 73219
rect 97905 73219 97963 73225
rect 97905 73216 97917 73219
rect 97399 73188 97917 73216
rect 97399 73185 97411 73188
rect 97353 73179 97411 73185
rect 97905 73185 97917 73188
rect 97951 73216 97963 73219
rect 99926 73216 99932 73228
rect 97951 73188 99932 73216
rect 97951 73185 97963 73188
rect 97905 73179 97963 73185
rect 99926 73176 99932 73188
rect 99984 73176 99990 73228
rect 100312 73216 100340 73256
rect 101582 73244 101588 73256
rect 101640 73284 101646 73296
rect 101766 73284 101772 73296
rect 101640 73256 101772 73284
rect 101640 73244 101646 73256
rect 101766 73244 101772 73256
rect 101824 73284 101830 73296
rect 102980 73284 103008 73315
rect 103330 73312 103336 73364
rect 103388 73312 103394 73364
rect 103793 73355 103851 73361
rect 103793 73321 103805 73355
rect 103839 73352 103851 73355
rect 104618 73352 104624 73364
rect 103839 73324 104624 73352
rect 103839 73321 103851 73324
rect 103793 73315 103851 73321
rect 103146 73284 103152 73296
rect 101824 73256 103152 73284
rect 101824 73244 101830 73256
rect 103146 73244 103152 73256
rect 103204 73284 103210 73296
rect 103808 73284 103836 73315
rect 104618 73312 104624 73324
rect 104676 73312 104682 73364
rect 103204 73256 103836 73284
rect 103204 73244 103210 73256
rect 103974 73244 103980 73296
rect 104032 73284 104038 73296
rect 105446 73284 105452 73296
rect 104032 73256 105452 73284
rect 104032 73244 104038 73256
rect 105446 73244 105452 73256
rect 105504 73244 105510 73296
rect 106185 73287 106243 73293
rect 106185 73284 106197 73287
rect 105556 73256 106197 73284
rect 100128 73188 100340 73216
rect 100389 73219 100447 73225
rect 96985 73151 97043 73157
rect 96985 73148 96997 73151
rect 96948 73120 96997 73148
rect 96948 73108 96954 73120
rect 96985 73117 96997 73120
rect 97031 73117 97043 73151
rect 96985 73111 97043 73117
rect 97077 73151 97135 73157
rect 97077 73117 97089 73151
rect 97123 73117 97135 73151
rect 97077 73111 97135 73117
rect 97169 73151 97227 73157
rect 97169 73117 97181 73151
rect 97215 73148 97227 73151
rect 97534 73148 97540 73160
rect 97215 73120 97540 73148
rect 97215 73117 97227 73120
rect 97169 73111 97227 73117
rect 40221 73083 40279 73089
rect 40221 73049 40233 73083
rect 40267 73080 40279 73083
rect 70121 73083 70179 73089
rect 40267 73052 41414 73080
rect 40267 73049 40279 73052
rect 40221 73043 40279 73049
rect 39853 73015 39911 73021
rect 39853 72981 39865 73015
rect 39899 72981 39911 73015
rect 41386 73012 41414 73052
rect 70121 73049 70133 73083
rect 70167 73080 70179 73083
rect 70210 73080 70216 73092
rect 70167 73052 70216 73080
rect 70167 73049 70179 73052
rect 70121 73043 70179 73049
rect 70210 73040 70216 73052
rect 70268 73040 70274 73092
rect 70394 73040 70400 73092
rect 70452 73080 70458 73092
rect 72697 73083 72755 73089
rect 72697 73080 72709 73083
rect 70452 73052 72709 73080
rect 70452 73040 70458 73052
rect 72697 73049 72709 73052
rect 72743 73049 72755 73083
rect 72697 73043 72755 73049
rect 79904 73083 79962 73089
rect 79904 73049 79916 73083
rect 79950 73080 79962 73083
rect 81986 73080 81992 73092
rect 79950 73052 81992 73080
rect 79950 73049 79962 73052
rect 79904 73043 79962 73049
rect 81986 73040 81992 73052
rect 82044 73040 82050 73092
rect 97000 73080 97028 73111
rect 97534 73108 97540 73120
rect 97592 73108 97598 73160
rect 97629 73151 97687 73157
rect 97629 73117 97641 73151
rect 97675 73117 97687 73151
rect 97629 73111 97687 73117
rect 97644 73080 97672 73111
rect 97718 73108 97724 73160
rect 97776 73108 97782 73160
rect 97813 73151 97871 73157
rect 97813 73117 97825 73151
rect 97859 73117 97871 73151
rect 97813 73111 97871 73117
rect 97828 73080 97856 73111
rect 98086 73108 98092 73160
rect 98144 73108 98150 73160
rect 98178 73108 98184 73160
rect 98236 73108 98242 73160
rect 98365 73151 98423 73157
rect 98365 73117 98377 73151
rect 98411 73117 98423 73151
rect 98365 73111 98423 73117
rect 98641 73151 98699 73157
rect 98641 73117 98653 73151
rect 98687 73117 98699 73151
rect 98641 73111 98699 73117
rect 99469 73151 99527 73157
rect 99469 73117 99481 73151
rect 99515 73117 99527 73151
rect 99469 73111 99527 73117
rect 97000 73052 97672 73080
rect 97736 73052 97856 73080
rect 42702 73012 42708 73024
rect 41386 72984 42708 73012
rect 39853 72975 39911 72981
rect 42702 72972 42708 72984
rect 42760 72972 42766 73024
rect 68833 73015 68891 73021
rect 68833 72981 68845 73015
rect 68879 73012 68891 73015
rect 69106 73012 69112 73024
rect 68879 72984 69112 73012
rect 68879 72981 68891 72984
rect 68833 72975 68891 72981
rect 69106 72972 69112 72984
rect 69164 72972 69170 73024
rect 73062 72972 73068 73024
rect 73120 72972 73126 73024
rect 96154 72972 96160 73024
rect 96212 73012 96218 73024
rect 96801 73015 96859 73021
rect 96801 73012 96813 73015
rect 96212 72984 96813 73012
rect 96212 72972 96218 72984
rect 96801 72981 96813 72984
rect 96847 72981 96859 73015
rect 96801 72975 96859 72981
rect 97442 72972 97448 73024
rect 97500 72972 97506 73024
rect 97534 72972 97540 73024
rect 97592 73012 97598 73024
rect 97736 73012 97764 73052
rect 97902 73040 97908 73092
rect 97960 73080 97966 73092
rect 98380 73080 98408 73111
rect 97960 73052 98408 73080
rect 97960 73040 97966 73052
rect 97592 72984 97764 73012
rect 97592 72972 97598 72984
rect 98270 72972 98276 73024
rect 98328 73012 98334 73024
rect 98656 73012 98684 73111
rect 99484 73080 99512 73111
rect 99650 73108 99656 73160
rect 99708 73148 99714 73160
rect 99745 73151 99803 73157
rect 99745 73148 99757 73151
rect 99708 73120 99757 73148
rect 99708 73108 99714 73120
rect 99745 73117 99757 73120
rect 99791 73117 99803 73151
rect 99745 73111 99803 73117
rect 100128 73080 100156 73188
rect 100389 73185 100401 73219
rect 100435 73216 100447 73219
rect 100435 73188 101076 73216
rect 100435 73185 100447 73188
rect 100389 73179 100447 73185
rect 100202 73108 100208 73160
rect 100260 73148 100266 73160
rect 100297 73151 100355 73157
rect 100297 73148 100309 73151
rect 100260 73120 100309 73148
rect 100260 73108 100266 73120
rect 100297 73117 100309 73120
rect 100343 73117 100355 73151
rect 100297 73111 100355 73117
rect 100481 73151 100539 73157
rect 100481 73117 100493 73151
rect 100527 73148 100539 73151
rect 100662 73148 100668 73160
rect 100527 73120 100668 73148
rect 100527 73117 100539 73120
rect 100481 73111 100539 73117
rect 100662 73108 100668 73120
rect 100720 73108 100726 73160
rect 101048 73157 101076 73188
rect 101858 73176 101864 73228
rect 101916 73216 101922 73228
rect 102229 73219 102287 73225
rect 102229 73216 102241 73219
rect 101916 73188 102241 73216
rect 101916 73176 101922 73188
rect 102229 73185 102241 73188
rect 102275 73185 102287 73219
rect 102229 73179 102287 73185
rect 102778 73176 102784 73228
rect 102836 73176 102842 73228
rect 103609 73219 103667 73225
rect 103609 73185 103621 73219
rect 103655 73216 103667 73219
rect 103790 73216 103796 73228
rect 103655 73188 103796 73216
rect 103655 73185 103667 73188
rect 103609 73179 103667 73185
rect 103790 73176 103796 73188
rect 103848 73176 103854 73228
rect 104434 73176 104440 73228
rect 104492 73216 104498 73228
rect 104529 73219 104587 73225
rect 104529 73216 104541 73219
rect 104492 73188 104541 73216
rect 104492 73176 104498 73188
rect 104529 73185 104541 73188
rect 104575 73185 104587 73219
rect 104529 73179 104587 73185
rect 101033 73151 101091 73157
rect 101033 73117 101045 73151
rect 101079 73117 101091 73151
rect 101033 73111 101091 73117
rect 102965 73151 103023 73157
rect 102965 73117 102977 73151
rect 103011 73148 103023 73151
rect 103238 73148 103244 73160
rect 103011 73120 103244 73148
rect 103011 73117 103023 73120
rect 102965 73111 103023 73117
rect 103238 73108 103244 73120
rect 103296 73108 103302 73160
rect 103885 73151 103943 73157
rect 103885 73117 103897 73151
rect 103931 73148 103943 73151
rect 104069 73151 104127 73157
rect 104069 73148 104081 73151
rect 103931 73120 104081 73148
rect 103931 73117 103943 73120
rect 103885 73111 103943 73117
rect 104069 73117 104081 73120
rect 104115 73117 104127 73151
rect 104069 73111 104127 73117
rect 99484 73052 100156 73080
rect 100941 73083 100999 73089
rect 100941 73049 100953 73083
rect 100987 73049 100999 73083
rect 100941 73043 100999 73049
rect 98328 72984 98684 73012
rect 98328 72972 98334 72984
rect 99190 72972 99196 73024
rect 99248 72972 99254 73024
rect 100478 72972 100484 73024
rect 100536 73012 100542 73024
rect 100731 73015 100789 73021
rect 100731 73012 100743 73015
rect 100536 72984 100743 73012
rect 100536 72972 100542 72984
rect 100731 72981 100743 72984
rect 100777 72981 100789 73015
rect 100956 73012 100984 73043
rect 101214 73040 101220 73092
rect 101272 73040 101278 73092
rect 101401 73083 101459 73089
rect 101401 73049 101413 73083
rect 101447 73080 101459 73083
rect 102045 73083 102103 73089
rect 102045 73080 102057 73083
rect 101447 73052 102057 73080
rect 101447 73049 101459 73052
rect 101401 73043 101459 73049
rect 102045 73049 102057 73052
rect 102091 73049 102103 73083
rect 102045 73043 102103 73049
rect 102502 73040 102508 73092
rect 102560 73040 102566 73092
rect 103900 73080 103928 73111
rect 104618 73108 104624 73160
rect 104676 73148 104682 73160
rect 105556 73148 105584 73256
rect 106185 73253 106197 73256
rect 106231 73253 106243 73287
rect 106185 73247 106243 73253
rect 106200 73188 106412 73216
rect 104676 73120 105584 73148
rect 104676 73108 104682 73120
rect 105630 73108 105636 73160
rect 105688 73108 105694 73160
rect 106001 73151 106059 73157
rect 106001 73117 106013 73151
rect 106047 73148 106059 73151
rect 106200 73148 106228 73188
rect 106047 73120 106228 73148
rect 106277 73151 106335 73157
rect 106047 73117 106059 73120
rect 106001 73111 106059 73117
rect 106277 73117 106289 73151
rect 106323 73117 106335 73151
rect 106384 73148 106412 73188
rect 108114 73148 108120 73160
rect 106384 73120 108120 73148
rect 106277 73111 106335 73117
rect 103164 73052 103928 73080
rect 104161 73083 104219 73089
rect 101490 73012 101496 73024
rect 100956 72984 101496 73012
rect 100731 72975 100789 72981
rect 101490 72972 101496 72984
rect 101548 72972 101554 73024
rect 101766 72972 101772 73024
rect 101824 73012 101830 73024
rect 103164 73021 103192 73052
rect 104161 73049 104173 73083
rect 104207 73080 104219 73083
rect 106292 73080 106320 73111
rect 108114 73108 108120 73120
rect 108172 73108 108178 73160
rect 108209 73151 108267 73157
rect 108209 73117 108221 73151
rect 108255 73148 108267 73151
rect 108482 73148 108488 73160
rect 108255 73120 108488 73148
rect 108255 73117 108267 73120
rect 108209 73111 108267 73117
rect 108482 73108 108488 73120
rect 108540 73108 108546 73160
rect 104207 73052 108344 73080
rect 104207 73049 104219 73052
rect 104161 73043 104219 73049
rect 102137 73015 102195 73021
rect 102137 73012 102149 73015
rect 101824 72984 102149 73012
rect 101824 72972 101830 72984
rect 102137 72981 102149 72984
rect 102183 72981 102195 73015
rect 102137 72975 102195 72981
rect 103149 73015 103207 73021
rect 103149 72981 103161 73015
rect 103195 72981 103207 73015
rect 103149 72975 103207 72981
rect 104250 72972 104256 73024
rect 104308 72972 104314 73024
rect 105262 72972 105268 73024
rect 105320 73012 105326 73024
rect 105449 73015 105507 73021
rect 105449 73012 105461 73015
rect 105320 72984 105461 73012
rect 105320 72972 105326 72984
rect 105449 72981 105461 72984
rect 105495 72981 105507 73015
rect 105449 72975 105507 72981
rect 105630 72972 105636 73024
rect 105688 73012 105694 73024
rect 108316 73021 108344 73052
rect 105817 73015 105875 73021
rect 105817 73012 105829 73015
rect 105688 72984 105829 73012
rect 105688 72972 105694 72984
rect 105817 72981 105829 72984
rect 105863 72981 105875 73015
rect 105817 72975 105875 72981
rect 108301 73015 108359 73021
rect 108301 72981 108313 73015
rect 108347 72981 108359 73015
rect 108301 72975 108359 72981
rect 1104 72922 108836 72944
rect 1104 72870 4874 72922
rect 4926 72870 4938 72922
rect 4990 72870 5002 72922
rect 5054 72870 5066 72922
rect 5118 72870 5130 72922
rect 5182 72870 35594 72922
rect 35646 72870 35658 72922
rect 35710 72870 35722 72922
rect 35774 72870 35786 72922
rect 35838 72870 35850 72922
rect 35902 72870 66314 72922
rect 66366 72870 66378 72922
rect 66430 72870 66442 72922
rect 66494 72870 66506 72922
rect 66558 72870 66570 72922
rect 66622 72870 97034 72922
rect 97086 72870 97098 72922
rect 97150 72870 97162 72922
rect 97214 72870 97226 72922
rect 97278 72870 97290 72922
rect 97342 72870 108836 72922
rect 1104 72848 108836 72870
rect 37826 72768 37832 72820
rect 37884 72808 37890 72820
rect 42886 72808 42892 72820
rect 37884 72780 42892 72808
rect 37884 72768 37890 72780
rect 42886 72768 42892 72780
rect 42944 72768 42950 72820
rect 69106 72808 69112 72820
rect 68848 72780 69112 72808
rect 37734 72700 37740 72752
rect 37792 72740 37798 72752
rect 42426 72740 42432 72752
rect 37792 72712 42432 72740
rect 37792 72700 37798 72712
rect 42426 72700 42432 72712
rect 42484 72700 42490 72752
rect 1673 72675 1731 72681
rect 1673 72641 1685 72675
rect 1719 72672 1731 72675
rect 1857 72675 1915 72681
rect 1857 72672 1869 72675
rect 1719 72644 1869 72672
rect 1719 72641 1731 72644
rect 1673 72635 1731 72641
rect 1857 72641 1869 72644
rect 1903 72672 1915 72675
rect 11698 72672 11704 72684
rect 1903 72644 11704 72672
rect 1903 72641 1915 72644
rect 1857 72635 1915 72641
rect 11698 72632 11704 72644
rect 11756 72632 11762 72684
rect 68848 72681 68876 72780
rect 69106 72768 69112 72780
rect 69164 72768 69170 72820
rect 73062 72768 73068 72820
rect 73120 72808 73126 72820
rect 73120 72780 80054 72808
rect 73120 72768 73126 72780
rect 68833 72675 68891 72681
rect 68833 72641 68845 72675
rect 68879 72641 68891 72675
rect 80026 72672 80054 72780
rect 85574 72768 85580 72820
rect 85632 72808 85638 72820
rect 86221 72811 86279 72817
rect 86221 72808 86233 72811
rect 85632 72780 86233 72808
rect 85632 72768 85638 72780
rect 86221 72777 86233 72780
rect 86267 72808 86279 72811
rect 86678 72808 86684 72820
rect 86267 72780 86684 72808
rect 86267 72777 86279 72780
rect 86221 72771 86279 72777
rect 86678 72768 86684 72780
rect 86736 72768 86742 72820
rect 88153 72811 88211 72817
rect 88153 72777 88165 72811
rect 88199 72777 88211 72811
rect 88153 72771 88211 72777
rect 97727 72811 97785 72817
rect 97727 72777 97739 72811
rect 97773 72808 97785 72811
rect 97902 72808 97908 72820
rect 97773 72780 97908 72808
rect 97773 72777 97785 72780
rect 97727 72771 97785 72777
rect 85482 72700 85488 72752
rect 85540 72740 85546 72752
rect 88168 72740 88196 72771
rect 97902 72768 97908 72780
rect 97960 72768 97966 72820
rect 98178 72768 98184 72820
rect 98236 72808 98242 72820
rect 98365 72811 98423 72817
rect 98365 72808 98377 72811
rect 98236 72780 98377 72808
rect 98236 72768 98242 72780
rect 98365 72777 98377 72780
rect 98411 72777 98423 72811
rect 98365 72771 98423 72777
rect 100018 72768 100024 72820
rect 100076 72768 100082 72820
rect 100846 72768 100852 72820
rect 100904 72808 100910 72820
rect 101214 72808 101220 72820
rect 100904 72780 101220 72808
rect 100904 72768 100910 72780
rect 101214 72768 101220 72780
rect 101272 72768 101278 72820
rect 103790 72768 103796 72820
rect 103848 72808 103854 72820
rect 104618 72808 104624 72820
rect 103848 72780 104624 72808
rect 103848 72768 103854 72780
rect 104618 72768 104624 72780
rect 104676 72768 104682 72820
rect 104805 72811 104863 72817
rect 104805 72777 104817 72811
rect 104851 72808 104863 72811
rect 105170 72808 105176 72820
rect 104851 72780 105176 72808
rect 104851 72777 104863 72780
rect 104805 72771 104863 72777
rect 105170 72768 105176 72780
rect 105228 72768 105234 72820
rect 105354 72768 105360 72820
rect 105412 72768 105418 72820
rect 105446 72768 105452 72820
rect 105504 72808 105510 72820
rect 105998 72808 106004 72820
rect 105504 72780 106004 72808
rect 105504 72768 105510 72780
rect 105998 72768 106004 72780
rect 106056 72768 106062 72820
rect 88337 72743 88395 72749
rect 88337 72740 88349 72743
rect 85540 72712 87170 72740
rect 88168 72712 88349 72740
rect 85540 72700 85546 72712
rect 88337 72709 88349 72712
rect 88383 72740 88395 72743
rect 94498 72740 94504 72752
rect 88383 72712 94504 72740
rect 88383 72709 88395 72712
rect 88337 72703 88395 72709
rect 94498 72700 94504 72712
rect 94556 72700 94562 72752
rect 96062 72700 96068 72752
rect 96120 72740 96126 72752
rect 97626 72740 97632 72752
rect 96120 72712 97632 72740
rect 96120 72700 96126 72712
rect 97626 72700 97632 72712
rect 97684 72700 97690 72752
rect 96433 72675 96491 72681
rect 80026 72644 86172 72672
rect 68833 72635 68891 72641
rect 842 72428 848 72480
rect 900 72468 906 72480
rect 1489 72471 1547 72477
rect 1489 72468 1501 72471
rect 900 72440 1501 72468
rect 900 72428 906 72440
rect 1489 72437 1501 72440
rect 1535 72437 1547 72471
rect 1489 72431 1547 72437
rect 86034 72428 86040 72480
rect 86092 72428 86098 72480
rect 86144 72468 86172 72644
rect 96433 72641 96445 72675
rect 96479 72672 96491 72675
rect 97718 72672 97724 72684
rect 96479 72644 97724 72672
rect 96479 72641 96491 72644
rect 96433 72635 96491 72641
rect 97718 72632 97724 72644
rect 97776 72632 97782 72684
rect 97813 72675 97871 72681
rect 97813 72641 97825 72675
rect 97859 72641 97871 72675
rect 97813 72635 97871 72641
rect 97905 72675 97963 72681
rect 97905 72641 97917 72675
rect 97951 72672 97963 72675
rect 98196 72672 98224 72768
rect 98454 72700 98460 72752
rect 98512 72740 98518 72752
rect 98549 72743 98607 72749
rect 98549 72740 98561 72743
rect 98512 72712 98561 72740
rect 98512 72700 98518 72712
rect 98549 72709 98561 72712
rect 98595 72740 98607 72743
rect 99101 72743 99159 72749
rect 99101 72740 99113 72743
rect 98595 72712 99113 72740
rect 98595 72709 98607 72712
rect 98549 72703 98607 72709
rect 99101 72709 99113 72712
rect 99147 72709 99159 72743
rect 99101 72703 99159 72709
rect 100588 72712 101904 72740
rect 97951 72644 98224 72672
rect 98273 72675 98331 72681
rect 97951 72641 97963 72644
rect 97905 72635 97963 72641
rect 98273 72641 98285 72675
rect 98319 72672 98331 72675
rect 98362 72672 98368 72684
rect 98319 72644 98368 72672
rect 98319 72641 98331 72644
rect 98273 72635 98331 72641
rect 86218 72564 86224 72616
rect 86276 72604 86282 72616
rect 86405 72607 86463 72613
rect 86405 72604 86417 72607
rect 86276 72576 86417 72604
rect 86276 72564 86282 72576
rect 86405 72573 86417 72576
rect 86451 72573 86463 72607
rect 86405 72567 86463 72573
rect 86678 72564 86684 72616
rect 86736 72564 86742 72616
rect 96525 72607 96583 72613
rect 96525 72573 96537 72607
rect 96571 72604 96583 72607
rect 97828 72604 97856 72635
rect 98362 72632 98368 72644
rect 98420 72632 98426 72684
rect 98730 72632 98736 72684
rect 98788 72632 98794 72684
rect 99285 72675 99343 72681
rect 99285 72641 99297 72675
rect 99331 72672 99343 72675
rect 99331 72644 100064 72672
rect 99331 72641 99343 72644
rect 99285 72635 99343 72641
rect 100036 72616 100064 72644
rect 100386 72632 100392 72684
rect 100444 72632 100450 72684
rect 98086 72604 98092 72616
rect 96571 72576 96752 72604
rect 96571 72573 96583 72576
rect 96525 72567 96583 72573
rect 89070 72468 89076 72480
rect 86144 72440 89076 72468
rect 89070 72428 89076 72440
rect 89128 72428 89134 72480
rect 96724 72468 96752 72576
rect 96816 72576 98092 72604
rect 96816 72545 96844 72576
rect 98086 72564 98092 72576
rect 98144 72604 98150 72616
rect 98546 72604 98552 72616
rect 98144 72576 98552 72604
rect 98144 72564 98150 72576
rect 98546 72564 98552 72576
rect 98604 72564 98610 72616
rect 99469 72607 99527 72613
rect 99469 72573 99481 72607
rect 99515 72604 99527 72607
rect 99558 72604 99564 72616
rect 99515 72576 99564 72604
rect 99515 72573 99527 72576
rect 99469 72567 99527 72573
rect 99558 72564 99564 72576
rect 99616 72564 99622 72616
rect 100018 72564 100024 72616
rect 100076 72604 100082 72616
rect 100588 72613 100616 72712
rect 101876 72684 101904 72712
rect 102778 72700 102784 72752
rect 102836 72700 102842 72752
rect 102965 72743 103023 72749
rect 102965 72709 102977 72743
rect 103011 72740 103023 72743
rect 104526 72740 104532 72752
rect 103011 72712 104532 72740
rect 103011 72709 103023 72712
rect 102965 72703 103023 72709
rect 100662 72632 100668 72684
rect 100720 72672 100726 72684
rect 101033 72675 101091 72681
rect 101033 72672 101045 72675
rect 100720 72644 101045 72672
rect 100720 72632 100726 72644
rect 101033 72641 101045 72644
rect 101079 72641 101091 72675
rect 101033 72635 101091 72641
rect 101122 72632 101128 72684
rect 101180 72632 101186 72684
rect 101582 72632 101588 72684
rect 101640 72632 101646 72684
rect 101769 72675 101827 72681
rect 101769 72641 101781 72675
rect 101815 72641 101827 72675
rect 101769 72635 101827 72641
rect 100481 72607 100539 72613
rect 100481 72604 100493 72607
rect 100076 72576 100493 72604
rect 100076 72564 100082 72576
rect 100481 72573 100493 72576
rect 100527 72573 100539 72607
rect 100481 72567 100539 72573
rect 100573 72607 100631 72613
rect 100573 72573 100585 72607
rect 100619 72573 100631 72607
rect 100573 72567 100631 72573
rect 96801 72539 96859 72545
rect 96801 72505 96813 72539
rect 96847 72505 96859 72539
rect 98270 72536 98276 72548
rect 96801 72499 96859 72505
rect 96908 72508 98276 72536
rect 96908 72468 96936 72508
rect 98270 72496 98276 72508
rect 98328 72496 98334 72548
rect 96724 72440 96936 72468
rect 97626 72428 97632 72480
rect 97684 72468 97690 72480
rect 98089 72471 98147 72477
rect 98089 72468 98101 72471
rect 97684 72440 98101 72468
rect 97684 72428 97690 72440
rect 98089 72437 98101 72440
rect 98135 72468 98147 72471
rect 100588 72468 100616 72567
rect 101490 72564 101496 72616
rect 101548 72604 101554 72616
rect 101784 72604 101812 72635
rect 101858 72632 101864 72684
rect 101916 72632 101922 72684
rect 102796 72672 102824 72700
rect 103517 72675 103575 72681
rect 103517 72672 103529 72675
rect 102796 72644 103529 72672
rect 103517 72641 103529 72644
rect 103563 72672 103575 72675
rect 103606 72672 103612 72684
rect 103563 72644 103612 72672
rect 103563 72641 103575 72644
rect 103517 72635 103575 72641
rect 103606 72632 103612 72644
rect 103664 72632 103670 72684
rect 103716 72681 103744 72712
rect 104526 72700 104532 72712
rect 104584 72700 104590 72752
rect 104636 72740 104664 72768
rect 104989 72743 105047 72749
rect 104989 72740 105001 72743
rect 104636 72712 105001 72740
rect 104989 72709 105001 72712
rect 105035 72709 105047 72743
rect 105372 72740 105400 72768
rect 105372 72712 105768 72740
rect 104989 72703 105047 72709
rect 103701 72675 103759 72681
rect 103701 72641 103713 72675
rect 103747 72641 103759 72675
rect 103701 72635 103759 72641
rect 103790 72632 103796 72684
rect 103848 72632 103854 72684
rect 104345 72675 104403 72681
rect 104345 72641 104357 72675
rect 104391 72672 104403 72675
rect 104544 72672 104572 72700
rect 104391 72644 104572 72672
rect 104621 72675 104679 72681
rect 104391 72641 104403 72644
rect 104345 72635 104403 72641
rect 104621 72641 104633 72675
rect 104667 72641 104679 72675
rect 104621 72635 104679 72641
rect 103330 72604 103336 72616
rect 101548 72576 103336 72604
rect 101548 72564 101554 72576
rect 103330 72564 103336 72576
rect 103388 72564 103394 72616
rect 103422 72564 103428 72616
rect 103480 72604 103486 72616
rect 104250 72604 104256 72616
rect 103480 72576 104256 72604
rect 103480 72564 103486 72576
rect 104250 72564 104256 72576
rect 104308 72604 104314 72616
rect 104529 72607 104587 72613
rect 104529 72604 104541 72607
rect 104308 72576 104541 72604
rect 104308 72564 104314 72576
rect 104529 72573 104541 72576
rect 104575 72573 104587 72607
rect 104529 72567 104587 72573
rect 101306 72496 101312 72548
rect 101364 72536 101370 72548
rect 101585 72539 101643 72545
rect 101585 72536 101597 72539
rect 101364 72508 101597 72536
rect 101364 72496 101370 72508
rect 101585 72505 101597 72508
rect 101631 72505 101643 72539
rect 101585 72499 101643 72505
rect 103514 72496 103520 72548
rect 103572 72536 103578 72548
rect 104437 72539 104495 72545
rect 104437 72536 104449 72539
rect 103572 72508 104449 72536
rect 103572 72496 103578 72508
rect 104437 72505 104449 72508
rect 104483 72505 104495 72539
rect 104636 72536 104664 72635
rect 104802 72632 104808 72684
rect 104860 72672 104866 72684
rect 104897 72675 104955 72681
rect 104897 72672 104909 72675
rect 104860 72644 104909 72672
rect 104860 72632 104866 72644
rect 104897 72641 104909 72644
rect 104943 72641 104955 72675
rect 104897 72635 104955 72641
rect 105173 72675 105231 72681
rect 105173 72641 105185 72675
rect 105219 72641 105231 72675
rect 105173 72635 105231 72641
rect 104710 72564 104716 72616
rect 104768 72604 104774 72616
rect 105188 72604 105216 72635
rect 105446 72632 105452 72684
rect 105504 72632 105510 72684
rect 105740 72681 105768 72712
rect 105924 72712 106320 72740
rect 105924 72684 105952 72712
rect 105725 72675 105783 72681
rect 105725 72641 105737 72675
rect 105771 72641 105783 72675
rect 105725 72635 105783 72641
rect 104768 72576 105216 72604
rect 105740 72604 105768 72635
rect 105906 72632 105912 72684
rect 105964 72632 105970 72684
rect 106292 72681 106320 72712
rect 106001 72675 106059 72681
rect 106001 72641 106013 72675
rect 106047 72641 106059 72675
rect 106001 72635 106059 72641
rect 106277 72675 106335 72681
rect 106277 72641 106289 72675
rect 106323 72641 106335 72675
rect 106277 72635 106335 72641
rect 108209 72675 108267 72681
rect 108209 72641 108221 72675
rect 108255 72672 108267 72675
rect 108482 72672 108488 72684
rect 108255 72644 108488 72672
rect 108255 72641 108267 72644
rect 108209 72635 108267 72641
rect 106016 72604 106044 72635
rect 108482 72632 108488 72644
rect 108540 72632 108546 72684
rect 105740 72576 106044 72604
rect 106093 72607 106151 72613
rect 104768 72564 104774 72576
rect 106093 72573 106105 72607
rect 106139 72573 106151 72607
rect 106093 72567 106151 72573
rect 104437 72499 104495 72505
rect 104544 72508 104664 72536
rect 98135 72440 100616 72468
rect 102597 72471 102655 72477
rect 98135 72437 98147 72440
rect 98089 72431 98147 72437
rect 102597 72437 102609 72471
rect 102643 72468 102655 72471
rect 103054 72468 103060 72480
rect 102643 72440 103060 72468
rect 102643 72437 102655 72440
rect 102597 72431 102655 72437
rect 103054 72428 103060 72440
rect 103112 72428 103118 72480
rect 103146 72428 103152 72480
rect 103204 72468 103210 72480
rect 103609 72471 103667 72477
rect 103609 72468 103621 72471
rect 103204 72440 103621 72468
rect 103204 72428 103210 72440
rect 103609 72437 103621 72440
rect 103655 72437 103667 72471
rect 103609 72431 103667 72437
rect 103698 72428 103704 72480
rect 103756 72468 103762 72480
rect 103977 72471 104035 72477
rect 103977 72468 103989 72471
rect 103756 72440 103989 72468
rect 103756 72428 103762 72440
rect 103977 72437 103989 72440
rect 104023 72468 104035 72471
rect 104544 72468 104572 72508
rect 105170 72496 105176 72548
rect 105228 72536 105234 72548
rect 105587 72539 105645 72545
rect 105587 72536 105599 72539
rect 105228 72508 105599 72536
rect 105228 72496 105234 72508
rect 105587 72505 105599 72508
rect 105633 72536 105645 72539
rect 106108 72536 106136 72567
rect 105633 72508 106136 72536
rect 105633 72505 105645 72508
rect 105587 72499 105645 72505
rect 104023 72440 104572 72468
rect 104023 72437 104035 72440
rect 103977 72431 104035 72437
rect 105814 72428 105820 72480
rect 105872 72428 105878 72480
rect 105998 72428 106004 72480
rect 106056 72428 106062 72480
rect 106090 72428 106096 72480
rect 106148 72468 106154 72480
rect 106461 72471 106519 72477
rect 106461 72468 106473 72471
rect 106148 72440 106473 72468
rect 106148 72428 106154 72440
rect 106461 72437 106473 72440
rect 106507 72437 106519 72471
rect 106461 72431 106519 72437
rect 108298 72428 108304 72480
rect 108356 72428 108362 72480
rect 1104 72378 108836 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 34934 72378
rect 34986 72326 34998 72378
rect 35050 72326 35062 72378
rect 35114 72326 35126 72378
rect 35178 72326 35190 72378
rect 35242 72326 65654 72378
rect 65706 72326 65718 72378
rect 65770 72326 65782 72378
rect 65834 72326 65846 72378
rect 65898 72326 65910 72378
rect 65962 72326 96374 72378
rect 96426 72326 96438 72378
rect 96490 72326 96502 72378
rect 96554 72326 96566 72378
rect 96618 72326 96630 72378
rect 96682 72326 108836 72378
rect 1104 72304 108836 72326
rect 81986 72224 81992 72276
rect 82044 72224 82050 72276
rect 85482 72224 85488 72276
rect 85540 72224 85546 72276
rect 88150 72224 88156 72276
rect 88208 72264 88214 72276
rect 88705 72267 88763 72273
rect 88705 72264 88717 72267
rect 88208 72236 88717 72264
rect 88208 72224 88214 72236
rect 85114 72156 85120 72208
rect 85172 72196 85178 72208
rect 85669 72199 85727 72205
rect 85669 72196 85681 72199
rect 85172 72168 85681 72196
rect 85172 72156 85178 72168
rect 85206 72128 85212 72140
rect 83292 72100 85212 72128
rect 83113 72063 83171 72069
rect 83113 72029 83125 72063
rect 83159 72060 83171 72063
rect 83292 72060 83320 72100
rect 85206 72088 85212 72100
rect 85264 72088 85270 72140
rect 85408 72072 85436 72168
rect 85669 72165 85681 72168
rect 85715 72165 85727 72199
rect 85669 72159 85727 72165
rect 83159 72032 83320 72060
rect 83369 72063 83427 72069
rect 83159 72029 83171 72032
rect 83113 72023 83171 72029
rect 83369 72029 83381 72063
rect 83415 72060 83427 72063
rect 83415 72032 83504 72060
rect 83415 72029 83427 72032
rect 83369 72023 83427 72029
rect 83476 71936 83504 72032
rect 85390 72020 85396 72072
rect 85448 72020 85454 72072
rect 88444 72069 88472 72236
rect 88705 72233 88717 72236
rect 88751 72264 88763 72267
rect 89714 72264 89720 72276
rect 88751 72236 89720 72264
rect 88751 72233 88763 72236
rect 88705 72227 88763 72233
rect 89714 72224 89720 72236
rect 89772 72224 89778 72276
rect 94498 72224 94504 72276
rect 94556 72264 94562 72276
rect 99009 72267 99067 72273
rect 94556 72236 98592 72264
rect 94556 72224 94562 72236
rect 93946 72156 93952 72208
rect 94004 72156 94010 72208
rect 97626 72196 97632 72208
rect 97460 72168 97632 72196
rect 93964 72128 93992 72156
rect 93412 72100 93992 72128
rect 93412 72069 93440 72100
rect 96798 72088 96804 72140
rect 96856 72088 96862 72140
rect 97460 72137 97488 72168
rect 97626 72156 97632 72168
rect 97684 72156 97690 72208
rect 98454 72156 98460 72208
rect 98512 72156 98518 72208
rect 98564 72196 98592 72236
rect 99009 72233 99021 72267
rect 99055 72264 99067 72267
rect 99098 72264 99104 72276
rect 99055 72236 99104 72264
rect 99055 72233 99067 72236
rect 99009 72227 99067 72233
rect 99098 72224 99104 72236
rect 99156 72224 99162 72276
rect 101217 72267 101275 72273
rect 101217 72233 101229 72267
rect 101263 72264 101275 72267
rect 101766 72264 101772 72276
rect 101263 72236 101772 72264
rect 101263 72233 101275 72236
rect 101217 72227 101275 72233
rect 101766 72224 101772 72236
rect 101824 72224 101830 72276
rect 103238 72224 103244 72276
rect 103296 72264 103302 72276
rect 104345 72267 104403 72273
rect 104345 72264 104357 72267
rect 103296 72236 104357 72264
rect 103296 72224 103302 72236
rect 104345 72233 104357 72236
rect 104391 72264 104403 72267
rect 104710 72264 104716 72276
rect 104391 72236 104716 72264
rect 104391 72233 104403 72236
rect 104345 72227 104403 72233
rect 104710 72224 104716 72236
rect 104768 72224 104774 72276
rect 104066 72196 104072 72208
rect 98564 72168 104072 72196
rect 104066 72156 104072 72168
rect 104124 72156 104130 72208
rect 107286 72196 107292 72208
rect 104176 72168 107292 72196
rect 97077 72131 97135 72137
rect 97077 72097 97089 72131
rect 97123 72097 97135 72131
rect 97077 72091 97135 72097
rect 97445 72131 97503 72137
rect 97445 72097 97457 72131
rect 97491 72097 97503 72131
rect 97445 72091 97503 72097
rect 98365 72131 98423 72137
rect 98365 72097 98377 72131
rect 98411 72128 98423 72131
rect 98730 72128 98736 72140
rect 98411 72100 98736 72128
rect 98411 72097 98423 72100
rect 98365 72091 98423 72097
rect 93578 72069 93584 72072
rect 88429 72063 88487 72069
rect 88429 72029 88441 72063
rect 88475 72029 88487 72063
rect 88429 72023 88487 72029
rect 93397 72063 93455 72069
rect 93397 72029 93409 72063
rect 93443 72029 93455 72063
rect 93397 72023 93455 72029
rect 93545 72063 93584 72069
rect 93545 72029 93557 72063
rect 93545 72023 93584 72029
rect 93578 72020 93584 72023
rect 93636 72020 93642 72072
rect 93903 72063 93961 72069
rect 93903 72029 93915 72063
rect 93949 72060 93961 72063
rect 94314 72060 94320 72072
rect 93949 72032 94320 72060
rect 93949 72029 93961 72032
rect 93903 72023 93961 72029
rect 94314 72020 94320 72032
rect 94372 72020 94378 72072
rect 96706 72020 96712 72072
rect 96764 72020 96770 72072
rect 97092 72060 97120 72091
rect 98730 72088 98736 72100
rect 98788 72128 98794 72140
rect 99561 72131 99619 72137
rect 99561 72128 99573 72131
rect 98788 72100 99573 72128
rect 98788 72088 98794 72100
rect 99561 72097 99573 72100
rect 99607 72097 99619 72131
rect 100846 72128 100852 72140
rect 99561 72091 99619 72097
rect 99760 72100 100852 72128
rect 97537 72063 97595 72069
rect 97537 72060 97549 72063
rect 97092 72032 97549 72060
rect 97537 72029 97549 72032
rect 97583 72029 97595 72063
rect 97537 72023 97595 72029
rect 97629 72063 97687 72069
rect 97629 72029 97641 72063
rect 97675 72060 97687 72063
rect 97994 72060 98000 72072
rect 97675 72032 98000 72060
rect 97675 72029 97687 72032
rect 97629 72023 97687 72029
rect 97994 72020 98000 72032
rect 98052 72020 98058 72072
rect 98086 72020 98092 72072
rect 98144 72020 98150 72072
rect 98273 72063 98331 72069
rect 98273 72029 98285 72063
rect 98319 72029 98331 72063
rect 98273 72023 98331 72029
rect 88521 71995 88579 72001
rect 88521 71961 88533 71995
rect 88567 71992 88579 71995
rect 90082 71992 90088 72004
rect 88567 71964 90088 71992
rect 88567 71961 88579 71964
rect 88521 71955 88579 71961
rect 90082 71952 90088 71964
rect 90140 71952 90146 72004
rect 93673 71995 93731 72001
rect 93673 71961 93685 71995
rect 93719 71961 93731 71995
rect 93673 71955 93731 71961
rect 83458 71884 83464 71936
rect 83516 71884 83522 71936
rect 93688 71924 93716 71955
rect 93762 71952 93768 72004
rect 93820 71952 93826 72004
rect 98288 71992 98316 72023
rect 98546 72020 98552 72072
rect 98604 72020 98610 72072
rect 99760 72069 99788 72100
rect 100846 72088 100852 72100
rect 100904 72088 100910 72140
rect 102318 72088 102324 72140
rect 102376 72128 102382 72140
rect 103974 72128 103980 72140
rect 102376 72100 103980 72128
rect 102376 72088 102382 72100
rect 103974 72088 103980 72100
rect 104032 72088 104038 72140
rect 99745 72063 99803 72069
rect 99745 72029 99757 72063
rect 99791 72029 99803 72063
rect 99745 72023 99803 72029
rect 100018 72020 100024 72072
rect 100076 72020 100082 72072
rect 100205 72063 100263 72069
rect 100205 72029 100217 72063
rect 100251 72029 100263 72063
rect 100205 72023 100263 72029
rect 98012 71964 98316 71992
rect 93854 71924 93860 71936
rect 93688 71896 93860 71924
rect 93854 71884 93860 71896
rect 93912 71884 93918 71936
rect 94041 71927 94099 71933
rect 94041 71893 94053 71927
rect 94087 71924 94099 71927
rect 95050 71924 95056 71936
rect 94087 71896 95056 71924
rect 94087 71893 94099 71896
rect 94041 71887 94099 71893
rect 95050 71884 95056 71896
rect 95108 71884 95114 71936
rect 98012 71933 98040 71964
rect 98362 71952 98368 72004
rect 98420 71992 98426 72004
rect 98733 71995 98791 72001
rect 98733 71992 98745 71995
rect 98420 71964 98745 71992
rect 98420 71952 98426 71964
rect 98733 71961 98745 71964
rect 98779 71961 98791 71995
rect 98733 71955 98791 71961
rect 99190 71952 99196 72004
rect 99248 71952 99254 72004
rect 99558 71952 99564 72004
rect 99616 71992 99622 72004
rect 100220 71992 100248 72023
rect 100294 72020 100300 72072
rect 100352 72060 100358 72072
rect 101125 72063 101183 72069
rect 101125 72060 101137 72063
rect 100352 72032 101137 72060
rect 100352 72020 100358 72032
rect 101125 72029 101137 72032
rect 101171 72029 101183 72063
rect 101125 72023 101183 72029
rect 101214 72020 101220 72072
rect 101272 72060 101278 72072
rect 101309 72063 101367 72069
rect 101309 72060 101321 72063
rect 101272 72032 101321 72060
rect 101272 72020 101278 72032
rect 101309 72029 101321 72032
rect 101355 72060 101367 72063
rect 102229 72063 102287 72069
rect 102229 72060 102241 72063
rect 101355 72032 102241 72060
rect 101355 72029 101367 72032
rect 101309 72023 101367 72029
rect 102229 72029 102241 72032
rect 102275 72060 102287 72063
rect 102502 72060 102508 72072
rect 102275 72032 102508 72060
rect 102275 72029 102287 72032
rect 102229 72023 102287 72029
rect 102502 72020 102508 72032
rect 102560 72020 102566 72072
rect 103054 72020 103060 72072
rect 103112 72020 103118 72072
rect 103146 72020 103152 72072
rect 103204 72020 103210 72072
rect 103422 72020 103428 72072
rect 103480 72020 103486 72072
rect 103514 72020 103520 72072
rect 103572 72020 103578 72072
rect 104176 72069 104204 72168
rect 107286 72156 107292 72168
rect 107344 72156 107350 72208
rect 105998 72128 106004 72140
rect 104820 72100 106004 72128
rect 104161 72063 104219 72069
rect 104161 72029 104173 72063
rect 104207 72029 104219 72063
rect 104161 72023 104219 72029
rect 104526 72020 104532 72072
rect 104584 72020 104590 72072
rect 104820 72069 104848 72100
rect 105998 72088 106004 72100
rect 106056 72088 106062 72140
rect 104805 72063 104863 72069
rect 104805 72029 104817 72063
rect 104851 72029 104863 72063
rect 104805 72023 104863 72029
rect 105262 72020 105268 72072
rect 105320 72020 105326 72072
rect 105354 72020 105360 72072
rect 105412 72060 105418 72072
rect 105541 72063 105599 72069
rect 105541 72060 105553 72063
rect 105412 72032 105553 72060
rect 105412 72020 105418 72032
rect 105541 72029 105553 72032
rect 105587 72029 105599 72063
rect 105541 72023 105599 72029
rect 99616 71964 100248 71992
rect 99616 71952 99622 71964
rect 101398 71952 101404 72004
rect 101456 71992 101462 72004
rect 103241 71995 103299 72001
rect 103241 71992 103253 71995
rect 101456 71964 103253 71992
rect 101456 71952 101462 71964
rect 103241 71961 103253 71964
rect 103287 71961 103299 71995
rect 103241 71955 103299 71961
rect 103330 71952 103336 72004
rect 103388 71992 103394 72004
rect 104894 71992 104900 72004
rect 103388 71964 104900 71992
rect 103388 71952 103394 71964
rect 104894 71952 104900 71964
rect 104952 71952 104958 72004
rect 105449 71995 105507 72001
rect 105449 71992 105461 71995
rect 105004 71964 105461 71992
rect 97997 71927 98055 71933
rect 97997 71893 98009 71927
rect 98043 71893 98055 71927
rect 97997 71887 98055 71893
rect 98638 71884 98644 71936
rect 98696 71924 98702 71936
rect 99006 71933 99012 71936
rect 98825 71927 98883 71933
rect 98825 71924 98837 71927
rect 98696 71896 98837 71924
rect 98696 71884 98702 71896
rect 98825 71893 98837 71896
rect 98871 71893 98883 71927
rect 98825 71887 98883 71893
rect 98993 71927 99012 71933
rect 98993 71893 99005 71927
rect 98993 71887 99012 71893
rect 99006 71884 99012 71887
rect 99064 71884 99070 71936
rect 100570 71884 100576 71936
rect 100628 71924 100634 71936
rect 102318 71924 102324 71936
rect 100628 71896 102324 71924
rect 100628 71884 100634 71896
rect 102318 71884 102324 71896
rect 102376 71884 102382 71936
rect 102778 71884 102784 71936
rect 102836 71924 102842 71936
rect 102873 71927 102931 71933
rect 102873 71924 102885 71927
rect 102836 71896 102885 71924
rect 102836 71884 102842 71896
rect 102873 71893 102885 71896
rect 102919 71893 102931 71927
rect 102873 71887 102931 71893
rect 103514 71884 103520 71936
rect 103572 71924 103578 71936
rect 103790 71924 103796 71936
rect 103572 71896 103796 71924
rect 103572 71884 103578 71896
rect 103790 71884 103796 71896
rect 103848 71924 103854 71936
rect 103885 71927 103943 71933
rect 103885 71924 103897 71927
rect 103848 71896 103897 71924
rect 103848 71884 103854 71896
rect 103885 71893 103897 71896
rect 103931 71924 103943 71927
rect 104434 71924 104440 71936
rect 103931 71896 104440 71924
rect 103931 71893 103943 71896
rect 103885 71887 103943 71893
rect 104434 71884 104440 71896
rect 104492 71924 104498 71936
rect 104802 71924 104808 71936
rect 104492 71896 104808 71924
rect 104492 71884 104498 71896
rect 104802 71884 104808 71896
rect 104860 71884 104866 71936
rect 105004 71933 105032 71964
rect 105449 71961 105461 71964
rect 105495 71961 105507 71995
rect 105556 71992 105584 72023
rect 105630 72020 105636 72072
rect 105688 72020 105694 72072
rect 105725 72063 105783 72069
rect 105725 72029 105737 72063
rect 105771 72060 105783 72063
rect 105814 72060 105820 72072
rect 105771 72032 105820 72060
rect 105771 72029 105783 72032
rect 105725 72023 105783 72029
rect 105814 72020 105820 72032
rect 105872 72060 105878 72072
rect 106185 72063 106243 72069
rect 106185 72060 106197 72063
rect 105872 72032 106197 72060
rect 105872 72020 105878 72032
rect 106185 72029 106197 72032
rect 106231 72029 106243 72063
rect 106185 72023 106243 72029
rect 105909 71995 105967 72001
rect 105909 71992 105921 71995
rect 105556 71964 105921 71992
rect 105449 71955 105507 71961
rect 105909 71961 105921 71964
rect 105955 71992 105967 71995
rect 106090 71992 106096 72004
rect 105955 71964 106096 71992
rect 105955 71961 105967 71964
rect 105909 71955 105967 71961
rect 106090 71952 106096 71964
rect 106148 71952 106154 72004
rect 104989 71927 105047 71933
rect 104989 71893 105001 71927
rect 105035 71893 105047 71927
rect 104989 71887 105047 71893
rect 105081 71927 105139 71933
rect 105081 71893 105093 71927
rect 105127 71924 105139 71927
rect 105538 71924 105544 71936
rect 105127 71896 105544 71924
rect 105127 71893 105139 71896
rect 105081 71887 105139 71893
rect 105538 71884 105544 71896
rect 105596 71884 105602 71936
rect 105814 71884 105820 71936
rect 105872 71884 105878 71936
rect 105998 71884 106004 71936
rect 106056 71884 106062 71936
rect 1104 71834 108836 71856
rect 1104 71782 4874 71834
rect 4926 71782 4938 71834
rect 4990 71782 5002 71834
rect 5054 71782 5066 71834
rect 5118 71782 5130 71834
rect 5182 71782 35594 71834
rect 35646 71782 35658 71834
rect 35710 71782 35722 71834
rect 35774 71782 35786 71834
rect 35838 71782 35850 71834
rect 35902 71782 66314 71834
rect 66366 71782 66378 71834
rect 66430 71782 66442 71834
rect 66494 71782 66506 71834
rect 66558 71782 66570 71834
rect 66622 71782 97034 71834
rect 97086 71782 97098 71834
rect 97150 71782 97162 71834
rect 97214 71782 97226 71834
rect 97278 71782 97290 71834
rect 97342 71782 108836 71834
rect 1104 71760 108836 71782
rect 91557 71723 91615 71729
rect 91557 71720 91569 71723
rect 91388 71692 91569 71720
rect 89622 71612 89628 71664
rect 89680 71612 89686 71664
rect 90082 71612 90088 71664
rect 90140 71612 90146 71664
rect 91388 71661 91416 71692
rect 91557 71689 91569 71692
rect 91603 71720 91615 71723
rect 92474 71720 92480 71732
rect 91603 71692 92480 71720
rect 91603 71689 91615 71692
rect 91557 71683 91615 71689
rect 92474 71680 92480 71692
rect 92532 71680 92538 71732
rect 96798 71680 96804 71732
rect 96856 71720 96862 71732
rect 96893 71723 96951 71729
rect 96893 71720 96905 71723
rect 96856 71692 96905 71720
rect 96856 71680 96862 71692
rect 96893 71689 96905 71692
rect 96939 71689 96951 71723
rect 96893 71683 96951 71689
rect 98086 71680 98092 71732
rect 98144 71720 98150 71732
rect 98181 71723 98239 71729
rect 98181 71720 98193 71723
rect 98144 71692 98193 71720
rect 98144 71680 98150 71692
rect 98181 71689 98193 71692
rect 98227 71689 98239 71723
rect 98181 71683 98239 71689
rect 98914 71680 98920 71732
rect 98972 71720 98978 71732
rect 100294 71720 100300 71732
rect 98972 71692 100300 71720
rect 98972 71680 98978 71692
rect 100294 71680 100300 71692
rect 100352 71680 100358 71732
rect 100386 71680 100392 71732
rect 100444 71720 100450 71732
rect 100481 71723 100539 71729
rect 100481 71720 100493 71723
rect 100444 71692 100493 71720
rect 100444 71680 100450 71692
rect 100481 71689 100493 71692
rect 100527 71689 100539 71723
rect 100481 71683 100539 71689
rect 101398 71680 101404 71732
rect 101456 71680 101462 71732
rect 104526 71720 104532 71732
rect 102612 71692 104532 71720
rect 91373 71655 91431 71661
rect 91373 71621 91385 71655
rect 91419 71621 91431 71655
rect 91373 71615 91431 71621
rect 96154 71612 96160 71664
rect 96212 71612 96218 71664
rect 98546 71652 98552 71664
rect 97184 71624 98552 71652
rect 1210 71544 1216 71596
rect 1268 71584 1274 71596
rect 97184 71593 97212 71624
rect 98546 71612 98552 71624
rect 98604 71612 98610 71664
rect 99190 71652 99196 71664
rect 98748 71624 99196 71652
rect 1489 71587 1547 71593
rect 1489 71584 1501 71587
rect 1268 71556 1501 71584
rect 1268 71544 1274 71556
rect 1489 71553 1501 71556
rect 1535 71584 1547 71587
rect 1949 71587 2007 71593
rect 1949 71584 1961 71587
rect 1535 71556 1961 71584
rect 1535 71553 1547 71556
rect 1489 71547 1547 71553
rect 1949 71553 1961 71556
rect 1995 71553 2007 71587
rect 1949 71547 2007 71553
rect 97168 71587 97226 71593
rect 97168 71553 97180 71587
rect 97214 71553 97226 71587
rect 97168 71547 97226 71553
rect 97261 71587 97319 71593
rect 97261 71553 97273 71587
rect 97307 71584 97319 71587
rect 97534 71584 97540 71596
rect 97307 71556 97540 71584
rect 97307 71553 97319 71556
rect 97261 71547 97319 71553
rect 97534 71544 97540 71556
rect 97592 71544 97598 71596
rect 97813 71587 97871 71593
rect 97813 71553 97825 71587
rect 97859 71553 97871 71587
rect 97813 71547 97871 71553
rect 89349 71519 89407 71525
rect 89349 71516 89361 71519
rect 89180 71488 89361 71516
rect 1673 71451 1731 71457
rect 1673 71417 1685 71451
rect 1719 71448 1731 71451
rect 1857 71451 1915 71457
rect 1857 71448 1869 71451
rect 1719 71420 1869 71448
rect 1719 71417 1731 71420
rect 1673 71411 1731 71417
rect 1857 71417 1869 71420
rect 1903 71448 1915 71451
rect 1903 71420 6914 71448
rect 1903 71417 1915 71420
rect 1857 71411 1915 71417
rect 6886 71380 6914 71420
rect 89180 71392 89208 71488
rect 89349 71485 89361 71488
rect 89395 71485 89407 71519
rect 97828 71516 97856 71547
rect 97902 71544 97908 71596
rect 97960 71584 97966 71596
rect 97997 71587 98055 71593
rect 97997 71584 98009 71587
rect 97960 71556 98009 71584
rect 97960 71544 97966 71556
rect 97997 71553 98009 71556
rect 98043 71553 98055 71587
rect 97997 71547 98055 71553
rect 98362 71544 98368 71596
rect 98420 71584 98426 71596
rect 98748 71593 98776 71624
rect 99190 71612 99196 71624
rect 99248 71652 99254 71664
rect 102612 71661 102640 71692
rect 104526 71680 104532 71692
rect 104584 71720 104590 71732
rect 108301 71723 108359 71729
rect 108301 71720 108313 71723
rect 104584 71692 108313 71720
rect 104584 71680 104590 71692
rect 108301 71689 108313 71692
rect 108347 71689 108359 71723
rect 108301 71683 108359 71689
rect 102597 71655 102655 71661
rect 99248 71624 99880 71652
rect 99248 71612 99254 71624
rect 99852 71596 99880 71624
rect 101324 71624 102180 71652
rect 98457 71587 98515 71593
rect 98457 71584 98469 71587
rect 98420 71556 98469 71584
rect 98420 71544 98426 71556
rect 98457 71553 98469 71556
rect 98503 71553 98515 71587
rect 98457 71547 98515 71553
rect 98733 71587 98791 71593
rect 98733 71553 98745 71587
rect 98779 71553 98791 71587
rect 99469 71587 99527 71593
rect 99469 71584 99481 71587
rect 98733 71547 98791 71553
rect 99346 71556 99481 71584
rect 98086 71516 98092 71528
rect 97828 71488 98092 71516
rect 89349 71479 89407 71485
rect 98086 71476 98092 71488
rect 98144 71476 98150 71528
rect 98472 71516 98500 71547
rect 99006 71516 99012 71528
rect 98472 71488 99012 71516
rect 99006 71476 99012 71488
rect 99064 71516 99070 71528
rect 99346 71516 99374 71556
rect 99469 71553 99481 71556
rect 99515 71553 99527 71587
rect 99469 71547 99527 71553
rect 99561 71587 99619 71593
rect 99561 71553 99573 71587
rect 99607 71553 99619 71587
rect 99561 71547 99619 71553
rect 99064 71488 99374 71516
rect 99064 71476 99070 71488
rect 94314 71408 94320 71460
rect 94372 71448 94378 71460
rect 95881 71451 95939 71457
rect 94372 71420 95832 71448
rect 94372 71408 94378 71420
rect 23474 71380 23480 71392
rect 6886 71352 23480 71380
rect 23474 71340 23480 71352
rect 23532 71340 23538 71392
rect 36170 71340 36176 71392
rect 36228 71380 36234 71392
rect 84838 71380 84844 71392
rect 36228 71352 84844 71380
rect 36228 71340 36234 71352
rect 84838 71340 84844 71352
rect 84896 71340 84902 71392
rect 89162 71340 89168 71392
rect 89220 71340 89226 71392
rect 95694 71340 95700 71392
rect 95752 71340 95758 71392
rect 95804 71380 95832 71420
rect 95881 71417 95893 71451
rect 95927 71448 95939 71451
rect 97442 71448 97448 71460
rect 95927 71420 97448 71448
rect 95927 71417 95939 71420
rect 95881 71411 95939 71417
rect 97442 71408 97448 71420
rect 97500 71408 97506 71460
rect 97626 71408 97632 71460
rect 97684 71448 97690 71460
rect 97684 71420 98316 71448
rect 97684 71408 97690 71420
rect 97902 71380 97908 71392
rect 95804 71352 97908 71380
rect 97902 71340 97908 71352
rect 97960 71340 97966 71392
rect 98288 71380 98316 71420
rect 98546 71408 98552 71460
rect 98604 71448 98610 71460
rect 99098 71448 99104 71460
rect 98604 71420 99104 71448
rect 98604 71408 98610 71420
rect 99098 71408 99104 71420
rect 99156 71448 99162 71460
rect 99576 71448 99604 71547
rect 99742 71544 99748 71596
rect 99800 71544 99806 71596
rect 99834 71544 99840 71596
rect 99892 71544 99898 71596
rect 100846 71544 100852 71596
rect 100904 71544 100910 71596
rect 101324 71593 101352 71624
rect 102152 71596 102180 71624
rect 102597 71621 102609 71655
rect 102643 71621 102655 71655
rect 104345 71655 104403 71661
rect 104345 71652 104357 71655
rect 102597 71615 102655 71621
rect 103440 71624 104357 71652
rect 101309 71587 101367 71593
rect 101309 71553 101321 71587
rect 101355 71553 101367 71587
rect 101309 71547 101367 71553
rect 101766 71544 101772 71596
rect 101824 71544 101830 71596
rect 102134 71544 102140 71596
rect 102192 71584 102198 71596
rect 102229 71587 102287 71593
rect 102229 71584 102241 71587
rect 102192 71556 102241 71584
rect 102192 71544 102198 71556
rect 102229 71553 102241 71556
rect 102275 71553 102287 71587
rect 102229 71547 102287 71553
rect 102778 71544 102784 71596
rect 102836 71544 102842 71596
rect 102965 71587 103023 71593
rect 102965 71553 102977 71587
rect 103011 71584 103023 71587
rect 103238 71584 103244 71596
rect 103011 71556 103244 71584
rect 103011 71553 103023 71556
rect 102965 71547 103023 71553
rect 103238 71544 103244 71556
rect 103296 71544 103302 71596
rect 103440 71593 103468 71624
rect 104345 71621 104357 71624
rect 104391 71621 104403 71655
rect 104345 71615 104403 71621
rect 104894 71612 104900 71664
rect 104952 71652 104958 71664
rect 104952 71624 105676 71652
rect 104952 71612 104958 71624
rect 103425 71587 103483 71593
rect 103425 71553 103437 71587
rect 103471 71553 103483 71587
rect 103425 71547 103483 71553
rect 103517 71587 103575 71593
rect 103517 71553 103529 71587
rect 103563 71553 103575 71587
rect 103517 71547 103575 71553
rect 103701 71587 103759 71593
rect 103701 71553 103713 71587
rect 103747 71553 103759 71587
rect 103701 71547 103759 71553
rect 99156 71420 99604 71448
rect 99760 71448 99788 71544
rect 100294 71476 100300 71528
rect 100352 71516 100358 71528
rect 100757 71519 100815 71525
rect 100757 71516 100769 71519
rect 100352 71488 100769 71516
rect 100352 71476 100358 71488
rect 100757 71485 100769 71488
rect 100803 71485 100815 71519
rect 100757 71479 100815 71485
rect 101861 71519 101919 71525
rect 101861 71485 101873 71519
rect 101907 71516 101919 71519
rect 102873 71519 102931 71525
rect 101907 71488 102088 71516
rect 101907 71485 101919 71488
rect 101861 71479 101919 71485
rect 100570 71448 100576 71460
rect 99760 71420 100576 71448
rect 99156 71408 99162 71420
rect 100570 71408 100576 71420
rect 100628 71408 100634 71460
rect 98914 71380 98920 71392
rect 98288 71352 98920 71380
rect 98914 71340 98920 71352
rect 98972 71340 98978 71392
rect 99285 71383 99343 71389
rect 99285 71349 99297 71383
rect 99331 71380 99343 71383
rect 99374 71380 99380 71392
rect 99331 71352 99380 71380
rect 99331 71349 99343 71352
rect 99285 71343 99343 71349
rect 99374 71340 99380 71352
rect 99432 71380 99438 71392
rect 100662 71380 100668 71392
rect 99432 71352 100668 71380
rect 99432 71340 99438 71352
rect 100662 71340 100668 71352
rect 100720 71340 100726 71392
rect 102060 71380 102088 71488
rect 102873 71485 102885 71519
rect 102919 71516 102931 71519
rect 103532 71516 103560 71547
rect 102919 71488 103560 71516
rect 102919 71485 102931 71488
rect 102873 71479 102931 71485
rect 102137 71451 102195 71457
rect 102137 71417 102149 71451
rect 102183 71448 102195 71451
rect 103422 71448 103428 71460
rect 102183 71420 103428 71448
rect 102183 71417 102195 71420
rect 102137 71411 102195 71417
rect 103422 71408 103428 71420
rect 103480 71448 103486 71460
rect 103716 71448 103744 71547
rect 103790 71544 103796 71596
rect 103848 71544 103854 71596
rect 104253 71587 104311 71593
rect 104253 71553 104265 71587
rect 104299 71553 104311 71587
rect 104253 71547 104311 71553
rect 104268 71516 104296 71547
rect 104434 71544 104440 71596
rect 104492 71544 104498 71596
rect 104529 71587 104587 71593
rect 104529 71553 104541 71587
rect 104575 71584 104587 71587
rect 104618 71584 104624 71596
rect 104575 71556 104624 71584
rect 104575 71553 104587 71556
rect 104529 71547 104587 71553
rect 104618 71544 104624 71556
rect 104676 71544 104682 71596
rect 104710 71544 104716 71596
rect 104768 71544 104774 71596
rect 104986 71544 104992 71596
rect 105044 71544 105050 71596
rect 105354 71544 105360 71596
rect 105412 71544 105418 71596
rect 105648 71593 105676 71624
rect 105633 71587 105691 71593
rect 105633 71553 105645 71587
rect 105679 71584 105691 71587
rect 105722 71584 105728 71596
rect 105679 71556 105728 71584
rect 105679 71553 105691 71556
rect 105633 71547 105691 71553
rect 105722 71544 105728 71556
rect 105780 71544 105786 71596
rect 107749 71587 107807 71593
rect 107749 71553 107761 71587
rect 107795 71584 107807 71587
rect 108298 71584 108304 71596
rect 107795 71556 108304 71584
rect 107795 71553 107807 71556
rect 107749 71547 107807 71553
rect 108298 71544 108304 71556
rect 108356 71544 108362 71596
rect 108482 71544 108488 71596
rect 108540 71544 108546 71596
rect 105004 71516 105032 71544
rect 103480 71420 103744 71448
rect 103808 71488 105032 71516
rect 105541 71519 105599 71525
rect 103480 71408 103486 71420
rect 103808 71380 103836 71488
rect 105541 71485 105553 71519
rect 105587 71516 105599 71519
rect 105998 71516 106004 71528
rect 105587 71488 106004 71516
rect 105587 71485 105599 71488
rect 105541 71479 105599 71485
rect 105998 71476 106004 71488
rect 106056 71476 106062 71528
rect 108209 71519 108267 71525
rect 108209 71485 108221 71519
rect 108255 71516 108267 71519
rect 108500 71516 108528 71544
rect 108255 71488 108528 71516
rect 108255 71485 108267 71488
rect 108209 71479 108267 71485
rect 104621 71451 104679 71457
rect 104621 71417 104633 71451
rect 104667 71448 104679 71451
rect 104986 71448 104992 71460
rect 104667 71420 104992 71448
rect 104667 71417 104679 71420
rect 104621 71411 104679 71417
rect 104986 71408 104992 71420
rect 105044 71408 105050 71460
rect 102060 71352 103836 71380
rect 103882 71340 103888 71392
rect 103940 71380 103946 71392
rect 103977 71383 104035 71389
rect 103977 71380 103989 71383
rect 103940 71352 103989 71380
rect 103940 71340 103946 71352
rect 103977 71349 103989 71352
rect 104023 71349 104035 71383
rect 103977 71343 104035 71349
rect 104894 71340 104900 71392
rect 104952 71380 104958 71392
rect 105173 71383 105231 71389
rect 105173 71380 105185 71383
rect 104952 71352 105185 71380
rect 104952 71340 104958 71352
rect 105173 71349 105185 71352
rect 105219 71349 105231 71383
rect 105173 71343 105231 71349
rect 105354 71340 105360 71392
rect 105412 71380 105418 71392
rect 105817 71383 105875 71389
rect 105817 71380 105829 71383
rect 105412 71352 105829 71380
rect 105412 71340 105418 71352
rect 105817 71349 105829 71352
rect 105863 71349 105875 71383
rect 105817 71343 105875 71349
rect 106274 71340 106280 71392
rect 106332 71380 106338 71392
rect 107657 71383 107715 71389
rect 107657 71380 107669 71383
rect 106332 71352 107669 71380
rect 106332 71340 106338 71352
rect 107657 71349 107669 71352
rect 107703 71349 107715 71383
rect 107657 71343 107715 71349
rect 1104 71290 108836 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 34934 71290
rect 34986 71238 34998 71290
rect 35050 71238 35062 71290
rect 35114 71238 35126 71290
rect 35178 71238 35190 71290
rect 35242 71238 65654 71290
rect 65706 71238 65718 71290
rect 65770 71238 65782 71290
rect 65834 71238 65846 71290
rect 65898 71238 65910 71290
rect 65962 71238 96374 71290
rect 96426 71238 96438 71290
rect 96490 71238 96502 71290
rect 96554 71238 96566 71290
rect 96618 71238 96630 71290
rect 96682 71238 108836 71290
rect 1104 71216 108836 71238
rect 31573 71179 31631 71185
rect 31573 71145 31585 71179
rect 31619 71176 31631 71179
rect 31754 71176 31760 71188
rect 31619 71148 31760 71176
rect 31619 71145 31631 71148
rect 31573 71139 31631 71145
rect 31754 71136 31760 71148
rect 31812 71176 31818 71188
rect 33137 71179 33195 71185
rect 33137 71176 33149 71179
rect 31812 71148 33149 71176
rect 31812 71136 31818 71148
rect 33137 71145 33149 71148
rect 33183 71145 33195 71179
rect 33137 71139 33195 71145
rect 48593 71179 48651 71185
rect 48593 71145 48605 71179
rect 48639 71176 48651 71179
rect 55122 71176 55128 71188
rect 48639 71148 55128 71176
rect 48639 71145 48651 71148
rect 48593 71139 48651 71145
rect 33045 71043 33103 71049
rect 33045 71040 33057 71043
rect 32876 71012 33057 71040
rect 32876 70981 32904 71012
rect 33045 71009 33057 71012
rect 33091 71040 33103 71043
rect 48133 71043 48191 71049
rect 48133 71040 48145 71043
rect 33091 71012 41414 71040
rect 33091 71009 33103 71012
rect 33045 71003 33103 71009
rect 32861 70975 32919 70981
rect 22066 70944 31754 70972
rect 5258 70864 5264 70916
rect 5316 70904 5322 70916
rect 22066 70904 22094 70944
rect 5316 70876 22094 70904
rect 31726 70904 31754 70944
rect 32861 70941 32873 70975
rect 32907 70941 32919 70975
rect 41386 70972 41414 71012
rect 45526 71012 48145 71040
rect 45526 70972 45554 71012
rect 48133 71009 48145 71012
rect 48179 71040 48191 71043
rect 48608 71040 48636 71139
rect 55122 71136 55128 71148
rect 55180 71136 55186 71188
rect 74261 71179 74319 71185
rect 74261 71145 74273 71179
rect 74307 71176 74319 71179
rect 84010 71176 84016 71188
rect 74307 71148 84016 71176
rect 74307 71145 74319 71148
rect 74261 71139 74319 71145
rect 84010 71136 84016 71148
rect 84068 71136 84074 71188
rect 85206 71136 85212 71188
rect 85264 71176 85270 71188
rect 86310 71176 86316 71188
rect 85264 71148 86316 71176
rect 85264 71136 85270 71148
rect 86310 71136 86316 71148
rect 86368 71136 86374 71188
rect 92661 71179 92719 71185
rect 92661 71145 92673 71179
rect 92707 71176 92719 71179
rect 93302 71176 93308 71188
rect 92707 71148 93308 71176
rect 92707 71145 92719 71148
rect 92661 71139 92719 71145
rect 93302 71136 93308 71148
rect 93360 71176 93366 71188
rect 96525 71179 96583 71185
rect 93360 71148 94176 71176
rect 93360 71136 93366 71148
rect 85390 71068 85396 71120
rect 85448 71108 85454 71120
rect 85669 71111 85727 71117
rect 85669 71108 85681 71111
rect 85448 71080 85681 71108
rect 85448 71068 85454 71080
rect 85669 71077 85681 71080
rect 85715 71077 85727 71111
rect 85669 71071 85727 71077
rect 92474 71068 92480 71120
rect 92532 71108 92538 71120
rect 94148 71117 94176 71148
rect 96525 71145 96537 71179
rect 96571 71176 96583 71179
rect 96706 71176 96712 71188
rect 96571 71148 96712 71176
rect 96571 71145 96583 71148
rect 96525 71139 96583 71145
rect 96706 71136 96712 71148
rect 96764 71136 96770 71188
rect 98822 71176 98828 71188
rect 97828 71148 98828 71176
rect 92753 71111 92811 71117
rect 92753 71108 92765 71111
rect 92532 71080 92765 71108
rect 92532 71068 92538 71080
rect 92753 71077 92765 71080
rect 92799 71077 92811 71111
rect 92753 71071 92811 71077
rect 94133 71111 94191 71117
rect 94133 71077 94145 71111
rect 94179 71077 94191 71111
rect 97629 71111 97687 71117
rect 97629 71108 97641 71111
rect 94133 71071 94191 71077
rect 96724 71080 97641 71108
rect 48179 71012 48636 71040
rect 72605 71043 72663 71049
rect 48179 71009 48191 71012
rect 48133 71003 48191 71009
rect 72605 71009 72617 71043
rect 72651 71040 72663 71043
rect 72878 71040 72884 71052
rect 72651 71012 72884 71040
rect 72651 71009 72663 71012
rect 72605 71003 72663 71009
rect 72878 71000 72884 71012
rect 72936 71000 72942 71052
rect 85945 71043 86003 71049
rect 85945 71040 85957 71043
rect 83476 71012 85957 71040
rect 83476 70984 83504 71012
rect 85945 71009 85957 71012
rect 85991 71040 86003 71043
rect 86034 71040 86040 71052
rect 85991 71012 86040 71040
rect 85991 71009 86003 71012
rect 85945 71003 86003 71009
rect 86034 71000 86040 71012
rect 86092 71040 86098 71052
rect 88061 71043 88119 71049
rect 88061 71040 88073 71043
rect 86092 71012 88073 71040
rect 86092 71000 86098 71012
rect 88061 71009 88073 71012
rect 88107 71040 88119 71043
rect 89162 71040 89168 71052
rect 88107 71012 89168 71040
rect 88107 71009 88119 71012
rect 88061 71003 88119 71009
rect 89162 71000 89168 71012
rect 89220 71000 89226 71052
rect 92768 71040 92796 71071
rect 93121 71043 93179 71049
rect 93121 71040 93133 71043
rect 92768 71012 93133 71040
rect 93121 71009 93133 71012
rect 93167 71040 93179 71043
rect 93854 71040 93860 71052
rect 93167 71012 93860 71040
rect 93167 71009 93179 71012
rect 93121 71003 93179 71009
rect 93854 71000 93860 71012
rect 93912 71040 93918 71052
rect 94225 71043 94283 71049
rect 94225 71040 94237 71043
rect 93912 71012 94237 71040
rect 93912 71000 93918 71012
rect 94225 71009 94237 71012
rect 94271 71040 94283 71043
rect 94866 71040 94872 71052
rect 94271 71012 94872 71040
rect 94271 71009 94283 71012
rect 94225 71003 94283 71009
rect 94866 71000 94872 71012
rect 94924 71000 94930 71052
rect 41386 70944 45554 70972
rect 47305 70975 47363 70981
rect 32861 70935 32919 70941
rect 47305 70941 47317 70975
rect 47351 70972 47363 70975
rect 47351 70944 48452 70972
rect 47351 70941 47363 70944
rect 47305 70935 47363 70941
rect 47320 70904 47348 70935
rect 48424 70913 48452 70944
rect 68646 70932 68652 70984
rect 68704 70972 68710 70984
rect 79229 70975 79287 70981
rect 79229 70972 79241 70975
rect 68704 70944 79241 70972
rect 68704 70932 68710 70944
rect 79229 70941 79241 70944
rect 79275 70941 79287 70975
rect 79229 70935 79287 70941
rect 79413 70975 79471 70981
rect 79413 70941 79425 70975
rect 79459 70972 79471 70975
rect 79502 70972 79508 70984
rect 79459 70944 79508 70972
rect 79459 70941 79471 70944
rect 79413 70935 79471 70941
rect 31726 70876 47348 70904
rect 48409 70907 48467 70913
rect 5316 70864 5322 70876
rect 48409 70873 48421 70907
rect 48455 70904 48467 70907
rect 73126 70907 73184 70913
rect 73126 70904 73138 70907
rect 48455 70876 55214 70904
rect 48455 70873 48467 70876
rect 48409 70867 48467 70873
rect 30282 70796 30288 70848
rect 30340 70836 30346 70848
rect 34514 70836 34520 70848
rect 30340 70808 34520 70836
rect 30340 70796 30346 70808
rect 34514 70796 34520 70808
rect 34572 70796 34578 70848
rect 55186 70836 55214 70876
rect 72712 70876 73138 70904
rect 72712 70848 72740 70876
rect 73126 70873 73138 70876
rect 73172 70873 73184 70907
rect 79244 70904 79272 70935
rect 79502 70932 79508 70944
rect 79560 70972 79566 70984
rect 81069 70975 81127 70981
rect 81069 70972 81081 70975
rect 79560 70944 81081 70972
rect 79560 70932 79566 70944
rect 81069 70941 81081 70944
rect 81115 70972 81127 70975
rect 81158 70972 81164 70984
rect 81115 70944 81164 70972
rect 81115 70941 81127 70944
rect 81069 70935 81127 70941
rect 81158 70932 81164 70944
rect 81216 70972 81222 70984
rect 83458 70972 83464 70984
rect 81216 70944 83464 70972
rect 81216 70932 81222 70944
rect 83458 70932 83464 70944
rect 83516 70932 83522 70984
rect 85390 70932 85396 70984
rect 85448 70932 85454 70984
rect 93213 70975 93271 70981
rect 93213 70941 93225 70975
rect 93259 70941 93271 70975
rect 93213 70935 93271 70941
rect 79658 70907 79716 70913
rect 79658 70904 79670 70907
rect 79244 70876 79670 70904
rect 73126 70867 73184 70873
rect 79658 70873 79670 70876
rect 79704 70873 79716 70907
rect 79658 70867 79716 70873
rect 85485 70907 85543 70913
rect 85485 70873 85497 70907
rect 85531 70904 85543 70907
rect 85531 70876 86618 70904
rect 85531 70873 85543 70876
rect 85485 70867 85543 70873
rect 87782 70864 87788 70916
rect 87840 70864 87846 70916
rect 93228 70904 93256 70935
rect 93302 70932 93308 70984
rect 93360 70932 93366 70984
rect 93394 70932 93400 70984
rect 93452 70972 93458 70984
rect 96724 70981 96752 71080
rect 97629 71077 97641 71080
rect 97675 71108 97687 71111
rect 97718 71108 97724 71120
rect 97675 71080 97724 71108
rect 97675 71077 97687 71080
rect 97629 71071 97687 71077
rect 97718 71068 97724 71080
rect 97776 71068 97782 71120
rect 93765 70975 93823 70981
rect 93765 70972 93777 70975
rect 93452 70944 93777 70972
rect 93452 70932 93458 70944
rect 93765 70941 93777 70944
rect 93811 70972 93823 70975
rect 94409 70975 94467 70981
rect 94409 70972 94421 70975
rect 93811 70944 94421 70972
rect 93811 70941 93823 70944
rect 93765 70935 93823 70941
rect 94409 70941 94421 70944
rect 94455 70941 94467 70975
rect 94409 70935 94467 70941
rect 96709 70975 96767 70981
rect 96709 70941 96721 70975
rect 96755 70941 96767 70975
rect 96709 70935 96767 70941
rect 96798 70932 96804 70984
rect 96856 70972 96862 70984
rect 96985 70975 97043 70981
rect 96985 70972 96997 70975
rect 96856 70944 96997 70972
rect 96856 70932 96862 70944
rect 96985 70941 96997 70944
rect 97031 70941 97043 70975
rect 96985 70935 97043 70941
rect 97629 70975 97687 70981
rect 97629 70941 97641 70975
rect 97675 70972 97687 70975
rect 97718 70972 97724 70984
rect 97675 70944 97724 70972
rect 97675 70941 97687 70944
rect 97629 70935 97687 70941
rect 93949 70907 94007 70913
rect 93949 70904 93961 70907
rect 93228 70876 93961 70904
rect 93949 70873 93961 70876
rect 93995 70904 94007 70907
rect 94038 70904 94044 70916
rect 93995 70876 94044 70904
rect 93995 70873 94007 70876
rect 93949 70867 94007 70873
rect 94038 70864 94044 70876
rect 94096 70864 94102 70916
rect 97000 70904 97028 70935
rect 97718 70932 97724 70944
rect 97776 70932 97782 70984
rect 97828 70981 97856 71148
rect 98822 71136 98828 71148
rect 98880 71136 98886 71188
rect 99009 71179 99067 71185
rect 99009 71145 99021 71179
rect 99055 71176 99067 71179
rect 99374 71176 99380 71188
rect 99055 71148 99380 71176
rect 99055 71145 99067 71148
rect 99009 71139 99067 71145
rect 99374 71136 99380 71148
rect 99432 71136 99438 71188
rect 99561 71179 99619 71185
rect 99561 71145 99573 71179
rect 99607 71176 99619 71179
rect 100018 71176 100024 71188
rect 99607 71148 100024 71176
rect 99607 71145 99619 71148
rect 99561 71139 99619 71145
rect 98546 71068 98552 71120
rect 98604 71068 98610 71120
rect 97994 71000 98000 71052
rect 98052 71040 98058 71052
rect 98270 71040 98276 71052
rect 98052 71012 98276 71040
rect 98052 71000 98058 71012
rect 98270 71000 98276 71012
rect 98328 71040 98334 71052
rect 99650 71040 99656 71052
rect 98328 71012 98500 71040
rect 98328 71000 98334 71012
rect 98472 70981 98500 71012
rect 98656 71012 99656 71040
rect 98656 70984 98684 71012
rect 99650 71000 99656 71012
rect 99708 71000 99714 71052
rect 99944 71049 99972 71148
rect 100018 71136 100024 71148
rect 100076 71136 100082 71188
rect 100294 71136 100300 71188
rect 100352 71136 100358 71188
rect 105814 71136 105820 71188
rect 105872 71136 105878 71188
rect 107286 71136 107292 71188
rect 107344 71176 107350 71188
rect 108301 71179 108359 71185
rect 108301 71176 108313 71179
rect 107344 71148 108313 71176
rect 107344 71136 107350 71148
rect 108301 71145 108313 71148
rect 108347 71145 108359 71179
rect 108301 71139 108359 71145
rect 101858 71068 101864 71120
rect 101916 71068 101922 71120
rect 105998 71068 106004 71120
rect 106056 71108 106062 71120
rect 106369 71111 106427 71117
rect 106369 71108 106381 71111
rect 106056 71080 106381 71108
rect 106056 71068 106062 71080
rect 106369 71077 106381 71080
rect 106415 71077 106427 71111
rect 106369 71071 106427 71077
rect 99929 71043 99987 71049
rect 99929 71009 99941 71043
rect 99975 71009 99987 71043
rect 101876 71040 101904 71068
rect 103606 71040 103612 71052
rect 101876 71012 102087 71040
rect 99929 71003 99987 71009
rect 97813 70975 97871 70981
rect 97813 70941 97825 70975
rect 97859 70941 97871 70975
rect 97813 70935 97871 70941
rect 98089 70975 98147 70981
rect 98089 70941 98101 70975
rect 98135 70972 98147 70975
rect 98457 70975 98515 70981
rect 98135 70944 98408 70972
rect 98135 70941 98147 70944
rect 98089 70935 98147 70941
rect 98380 70904 98408 70944
rect 98457 70941 98469 70975
rect 98503 70941 98515 70975
rect 98457 70935 98515 70941
rect 98638 70932 98644 70984
rect 98696 70932 98702 70984
rect 98730 70932 98736 70984
rect 98788 70972 98794 70984
rect 99466 70981 99472 70984
rect 98917 70975 98975 70981
rect 98917 70972 98929 70975
rect 98788 70944 98929 70972
rect 98788 70932 98794 70944
rect 98917 70941 98929 70944
rect 98963 70941 98975 70975
rect 98917 70935 98975 70941
rect 99436 70975 99472 70981
rect 99436 70941 99448 70975
rect 99436 70935 99472 70941
rect 99466 70932 99472 70935
rect 99524 70932 99530 70984
rect 100018 70932 100024 70984
rect 100076 70932 100082 70984
rect 101030 70932 101036 70984
rect 101088 70932 101094 70984
rect 101861 70975 101919 70981
rect 101861 70941 101873 70975
rect 101907 70972 101919 70975
rect 101950 70972 101956 70984
rect 101907 70944 101956 70972
rect 101907 70941 101919 70944
rect 101861 70935 101919 70941
rect 101950 70932 101956 70944
rect 102008 70932 102014 70984
rect 102059 70981 102087 71012
rect 102244 71012 103612 71040
rect 102044 70975 102102 70981
rect 102044 70941 102056 70975
rect 102090 70941 102102 70975
rect 102044 70935 102102 70941
rect 102134 70932 102140 70984
rect 102192 70932 102198 70984
rect 102244 70981 102272 71012
rect 103606 71000 103612 71012
rect 103664 71040 103670 71052
rect 103701 71043 103759 71049
rect 103701 71040 103713 71043
rect 103664 71012 103713 71040
rect 103664 71000 103670 71012
rect 103701 71009 103713 71012
rect 103747 71009 103759 71043
rect 103701 71003 103759 71009
rect 103790 71000 103796 71052
rect 103848 71040 103854 71052
rect 104253 71043 104311 71049
rect 104253 71040 104265 71043
rect 103848 71012 104265 71040
rect 103848 71000 103854 71012
rect 104253 71009 104265 71012
rect 104299 71040 104311 71043
rect 104897 71043 104955 71049
rect 104897 71040 104909 71043
rect 104299 71012 104909 71040
rect 104299 71009 104311 71012
rect 104253 71003 104311 71009
rect 104897 71009 104909 71012
rect 104943 71009 104955 71043
rect 104897 71003 104955 71009
rect 105081 71043 105139 71049
rect 105081 71009 105093 71043
rect 105127 71040 105139 71043
rect 105262 71040 105268 71052
rect 105127 71012 105268 71040
rect 105127 71009 105139 71012
rect 105081 71003 105139 71009
rect 105262 71000 105268 71012
rect 105320 71000 105326 71052
rect 105538 71000 105544 71052
rect 105596 71000 105602 71052
rect 106182 71000 106188 71052
rect 106240 71040 106246 71052
rect 106240 71012 106412 71040
rect 106240 71000 106246 71012
rect 102229 70975 102287 70981
rect 102229 70941 102241 70975
rect 102275 70941 102287 70975
rect 102229 70935 102287 70941
rect 102413 70975 102471 70981
rect 102413 70941 102425 70975
rect 102459 70972 102471 70975
rect 102778 70972 102784 70984
rect 102459 70944 102784 70972
rect 102459 70941 102471 70944
rect 102413 70935 102471 70941
rect 102244 70904 102272 70935
rect 102778 70932 102784 70944
rect 102836 70932 102842 70984
rect 103422 70932 103428 70984
rect 103480 70972 103486 70984
rect 104345 70975 104403 70981
rect 104345 70972 104357 70975
rect 103480 70944 104357 70972
rect 103480 70932 103486 70944
rect 104345 70941 104357 70944
rect 104391 70941 104403 70975
rect 104345 70935 104403 70941
rect 105173 70975 105231 70981
rect 105173 70941 105185 70975
rect 105219 70972 105231 70975
rect 105814 70972 105820 70984
rect 105219 70944 105820 70972
rect 105219 70941 105231 70944
rect 105173 70935 105231 70941
rect 105814 70932 105820 70944
rect 105872 70972 105878 70984
rect 106384 70981 106412 71012
rect 106093 70975 106151 70981
rect 106093 70972 106105 70975
rect 105872 70944 106105 70972
rect 105872 70932 105878 70944
rect 106093 70941 106105 70944
rect 106139 70941 106151 70975
rect 106093 70935 106151 70941
rect 106369 70975 106427 70981
rect 106369 70941 106381 70975
rect 106415 70941 106427 70975
rect 106369 70935 106427 70941
rect 108209 70975 108267 70981
rect 108209 70941 108221 70975
rect 108255 70972 108267 70975
rect 108482 70972 108488 70984
rect 108255 70944 108488 70972
rect 108255 70941 108267 70944
rect 108209 70935 108267 70941
rect 97000 70876 98132 70904
rect 98380 70876 102272 70904
rect 102597 70907 102655 70913
rect 56134 70836 56140 70848
rect 55186 70808 56140 70836
rect 56134 70796 56140 70808
rect 56192 70796 56198 70848
rect 72694 70796 72700 70848
rect 72752 70796 72758 70848
rect 80793 70839 80851 70845
rect 80793 70805 80805 70839
rect 80839 70836 80851 70839
rect 89254 70836 89260 70848
rect 80839 70808 89260 70836
rect 80839 70805 80851 70808
rect 80793 70799 80851 70805
rect 89254 70796 89260 70808
rect 89312 70796 89318 70848
rect 92934 70796 92940 70848
rect 92992 70796 92998 70848
rect 93026 70796 93032 70848
rect 93084 70836 93090 70848
rect 93581 70839 93639 70845
rect 93581 70836 93593 70839
rect 93084 70808 93593 70836
rect 93084 70796 93090 70808
rect 93581 70805 93593 70808
rect 93627 70805 93639 70839
rect 93581 70799 93639 70805
rect 93854 70796 93860 70848
rect 93912 70796 93918 70848
rect 96890 70796 96896 70848
rect 96948 70796 96954 70848
rect 97534 70796 97540 70848
rect 97592 70836 97598 70848
rect 97902 70836 97908 70848
rect 97592 70808 97908 70836
rect 97592 70796 97598 70808
rect 97902 70796 97908 70808
rect 97960 70796 97966 70848
rect 97994 70796 98000 70848
rect 98052 70796 98058 70848
rect 98104 70836 98132 70876
rect 102597 70873 102609 70907
rect 102643 70904 102655 70907
rect 103054 70904 103060 70916
rect 102643 70876 103060 70904
rect 102643 70873 102655 70876
rect 102597 70867 102655 70873
rect 103054 70864 103060 70876
rect 103112 70864 103118 70916
rect 103517 70907 103575 70913
rect 103517 70873 103529 70907
rect 103563 70904 103575 70907
rect 105078 70904 105084 70916
rect 103563 70876 105084 70904
rect 103563 70873 103575 70876
rect 103517 70867 103575 70873
rect 105078 70864 105084 70876
rect 105136 70864 105142 70916
rect 105538 70864 105544 70916
rect 105596 70904 105602 70916
rect 106001 70907 106059 70913
rect 106001 70904 106013 70907
rect 105596 70876 106013 70904
rect 105596 70864 105602 70876
rect 106001 70873 106013 70876
rect 106047 70904 106059 70907
rect 106185 70907 106243 70913
rect 106185 70904 106197 70907
rect 106047 70876 106197 70904
rect 106047 70873 106059 70876
rect 106001 70867 106059 70873
rect 106185 70873 106197 70876
rect 106231 70873 106243 70907
rect 106185 70867 106243 70873
rect 98454 70836 98460 70848
rect 98104 70808 98460 70836
rect 98454 70796 98460 70808
rect 98512 70796 98518 70848
rect 98914 70796 98920 70848
rect 98972 70836 98978 70848
rect 99377 70839 99435 70845
rect 99377 70836 99389 70839
rect 98972 70808 99389 70836
rect 98972 70796 98978 70808
rect 99377 70805 99389 70808
rect 99423 70805 99435 70839
rect 99377 70799 99435 70805
rect 100018 70796 100024 70848
rect 100076 70836 100082 70848
rect 101125 70839 101183 70845
rect 101125 70836 101137 70839
rect 100076 70808 101137 70836
rect 100076 70796 100082 70808
rect 101125 70805 101137 70808
rect 101171 70836 101183 70839
rect 101766 70836 101772 70848
rect 101171 70808 101772 70836
rect 101171 70805 101183 70808
rect 101125 70799 101183 70805
rect 101766 70796 101772 70808
rect 101824 70796 101830 70848
rect 103146 70796 103152 70848
rect 103204 70796 103210 70848
rect 103609 70839 103667 70845
rect 103609 70805 103621 70839
rect 103655 70836 103667 70839
rect 103977 70839 104035 70845
rect 103977 70836 103989 70839
rect 103655 70808 103989 70836
rect 103655 70805 103667 70808
rect 103609 70799 103667 70805
rect 103977 70805 103989 70808
rect 104023 70805 104035 70839
rect 103977 70799 104035 70805
rect 105630 70796 105636 70848
rect 105688 70796 105694 70848
rect 105801 70839 105859 70845
rect 105801 70805 105813 70839
rect 105847 70836 105859 70839
rect 106384 70836 106412 70935
rect 108482 70932 108488 70944
rect 108540 70932 108546 70984
rect 105847 70808 106412 70836
rect 105847 70805 105859 70808
rect 105801 70799 105859 70805
rect 1104 70746 108836 70768
rect 1104 70694 4874 70746
rect 4926 70694 4938 70746
rect 4990 70694 5002 70746
rect 5054 70694 5066 70746
rect 5118 70694 5130 70746
rect 5182 70694 35594 70746
rect 35646 70694 35658 70746
rect 35710 70694 35722 70746
rect 35774 70694 35786 70746
rect 35838 70694 35850 70746
rect 35902 70694 66314 70746
rect 66366 70694 66378 70746
rect 66430 70694 66442 70746
rect 66494 70694 66506 70746
rect 66558 70694 66570 70746
rect 66622 70694 97034 70746
rect 97086 70694 97098 70746
rect 97150 70694 97162 70746
rect 97214 70694 97226 70746
rect 97278 70694 97290 70746
rect 97342 70694 108836 70746
rect 1104 70672 108836 70694
rect 30558 70592 30564 70644
rect 30616 70592 30622 70644
rect 32125 70635 32183 70641
rect 32125 70632 32137 70635
rect 31726 70604 32137 70632
rect 28442 70524 28448 70576
rect 28500 70564 28506 70576
rect 31726 70564 31754 70604
rect 32125 70601 32137 70604
rect 32171 70601 32183 70635
rect 32125 70595 32183 70601
rect 34514 70592 34520 70644
rect 34572 70592 34578 70644
rect 87782 70592 87788 70644
rect 87840 70632 87846 70644
rect 87969 70635 88027 70641
rect 87969 70632 87981 70635
rect 87840 70604 87981 70632
rect 87840 70592 87846 70604
rect 87969 70601 87981 70604
rect 88015 70601 88027 70635
rect 87969 70595 88027 70601
rect 88150 70592 88156 70644
rect 88208 70632 88214 70644
rect 93029 70635 93087 70641
rect 93029 70632 93041 70635
rect 88208 70604 93041 70632
rect 88208 70592 88214 70604
rect 93029 70601 93041 70604
rect 93075 70632 93087 70635
rect 93210 70632 93216 70644
rect 93075 70604 93216 70632
rect 93075 70601 93087 70604
rect 93029 70595 93087 70601
rect 93210 70592 93216 70604
rect 93268 70592 93274 70644
rect 97074 70592 97080 70644
rect 97132 70592 97138 70644
rect 97184 70604 99374 70632
rect 34333 70567 34391 70573
rect 34333 70564 34345 70567
rect 28500 70536 31754 70564
rect 31956 70536 34345 70564
rect 28500 70524 28506 70536
rect 31662 70456 31668 70508
rect 31720 70505 31726 70508
rect 31720 70459 31732 70505
rect 31720 70456 31726 70459
rect 31846 70456 31852 70508
rect 31904 70496 31910 70508
rect 31956 70505 31984 70536
rect 33520 70505 33548 70536
rect 34333 70533 34345 70536
rect 34379 70564 34391 70567
rect 35526 70564 35532 70576
rect 34379 70536 35532 70564
rect 34379 70533 34391 70536
rect 34333 70527 34391 70533
rect 35526 70524 35532 70536
rect 35584 70564 35590 70576
rect 35584 70536 35940 70564
rect 35584 70524 35590 70536
rect 35912 70505 35940 70536
rect 84838 70524 84844 70576
rect 84896 70564 84902 70576
rect 90177 70567 90235 70573
rect 90177 70564 90189 70567
rect 84896 70536 90189 70564
rect 84896 70524 84902 70536
rect 90177 70533 90189 70536
rect 90223 70564 90235 70567
rect 90358 70564 90364 70576
rect 90223 70536 90364 70564
rect 90223 70533 90235 70536
rect 90177 70527 90235 70533
rect 90358 70524 90364 70536
rect 90416 70564 90422 70576
rect 91189 70567 91247 70573
rect 91189 70564 91201 70567
rect 90416 70536 91201 70564
rect 90416 70524 90422 70536
rect 91189 70533 91201 70536
rect 91235 70533 91247 70567
rect 97184 70564 97212 70604
rect 97629 70567 97687 70573
rect 97629 70564 97641 70567
rect 91189 70527 91247 70533
rect 91572 70536 97212 70564
rect 97368 70536 97641 70564
rect 31941 70499 31999 70505
rect 31941 70496 31953 70499
rect 31904 70468 31953 70496
rect 31904 70456 31910 70468
rect 31941 70465 31953 70468
rect 31987 70465 31999 70499
rect 31941 70459 31999 70465
rect 33249 70499 33307 70505
rect 33249 70465 33261 70499
rect 33295 70496 33307 70499
rect 33505 70499 33563 70505
rect 33295 70468 33456 70496
rect 33295 70465 33307 70468
rect 33249 70459 33307 70465
rect 33428 70428 33456 70468
rect 33505 70465 33517 70499
rect 33551 70465 33563 70499
rect 33505 70459 33563 70465
rect 35641 70499 35699 70505
rect 35641 70465 35653 70499
rect 35687 70496 35699 70499
rect 35897 70499 35955 70505
rect 35687 70468 35848 70496
rect 35687 70465 35699 70468
rect 35641 70459 35699 70465
rect 34514 70428 34520 70440
rect 33428 70400 34520 70428
rect 34514 70388 34520 70400
rect 34572 70388 34578 70440
rect 35820 70428 35848 70468
rect 35897 70465 35909 70499
rect 35943 70465 35955 70499
rect 35897 70459 35955 70465
rect 88153 70499 88211 70505
rect 88153 70465 88165 70499
rect 88199 70496 88211 70499
rect 88794 70496 88800 70508
rect 88199 70468 88800 70496
rect 88199 70465 88211 70468
rect 88153 70459 88211 70465
rect 88794 70456 88800 70468
rect 88852 70456 88858 70508
rect 90913 70499 90971 70505
rect 90913 70465 90925 70499
rect 90959 70496 90971 70499
rect 91097 70499 91155 70505
rect 91097 70496 91109 70499
rect 90959 70468 91109 70496
rect 90959 70465 90971 70468
rect 90913 70459 90971 70465
rect 91097 70465 91109 70468
rect 91143 70496 91155 70499
rect 91572 70496 91600 70536
rect 91143 70468 91600 70496
rect 96065 70499 96123 70505
rect 91143 70465 91155 70468
rect 91097 70459 91155 70465
rect 96065 70465 96077 70499
rect 96111 70496 96123 70499
rect 97074 70496 97080 70508
rect 96111 70468 97080 70496
rect 96111 70465 96123 70468
rect 96065 70459 96123 70465
rect 97074 70456 97080 70468
rect 97132 70456 97138 70508
rect 97258 70456 97264 70508
rect 97316 70456 97322 70508
rect 41138 70428 41144 70440
rect 35820 70400 41144 70428
rect 41138 70388 41144 70400
rect 41196 70388 41202 70440
rect 88337 70431 88395 70437
rect 88337 70397 88349 70431
rect 88383 70428 88395 70431
rect 91002 70428 91008 70440
rect 88383 70400 91008 70428
rect 88383 70397 88395 70400
rect 88337 70391 88395 70397
rect 91002 70388 91008 70400
rect 91060 70388 91066 70440
rect 96157 70431 96215 70437
rect 96157 70397 96169 70431
rect 96203 70428 96215 70431
rect 96798 70428 96804 70440
rect 96203 70400 96804 70428
rect 96203 70397 96215 70400
rect 96157 70391 96215 70397
rect 96798 70388 96804 70400
rect 96856 70388 96862 70440
rect 96433 70363 96491 70369
rect 96433 70329 96445 70363
rect 96479 70360 96491 70363
rect 97368 70360 97396 70536
rect 97629 70533 97641 70536
rect 97675 70533 97687 70567
rect 97629 70527 97687 70533
rect 97902 70524 97908 70576
rect 97960 70564 97966 70576
rect 97960 70536 98316 70564
rect 97960 70524 97966 70536
rect 97721 70499 97779 70505
rect 97721 70465 97733 70499
rect 97767 70496 97779 70499
rect 97810 70496 97816 70508
rect 97767 70468 97816 70496
rect 97767 70465 97779 70468
rect 97721 70459 97779 70465
rect 97810 70456 97816 70468
rect 97868 70456 97874 70508
rect 98178 70456 98184 70508
rect 98236 70456 98242 70508
rect 98288 70505 98316 70536
rect 98362 70524 98368 70576
rect 98420 70564 98426 70576
rect 98733 70567 98791 70573
rect 98733 70564 98745 70567
rect 98420 70536 98745 70564
rect 98420 70524 98426 70536
rect 98733 70533 98745 70536
rect 98779 70533 98791 70567
rect 99346 70564 99374 70604
rect 99466 70592 99472 70644
rect 99524 70592 99530 70644
rect 99576 70604 102456 70632
rect 99576 70564 99604 70604
rect 99346 70536 99604 70564
rect 98733 70527 98791 70533
rect 99650 70524 99656 70576
rect 99708 70564 99714 70576
rect 102428 70564 102456 70604
rect 103606 70592 103612 70644
rect 103664 70592 103670 70644
rect 105262 70592 105268 70644
rect 105320 70632 105326 70644
rect 106182 70632 106188 70644
rect 105320 70604 106188 70632
rect 105320 70592 105326 70604
rect 106182 70592 106188 70604
rect 106240 70592 106246 70644
rect 108114 70592 108120 70644
rect 108172 70632 108178 70644
rect 108301 70635 108359 70641
rect 108301 70632 108313 70635
rect 108172 70604 108313 70632
rect 108172 70592 108178 70604
rect 108301 70601 108313 70604
rect 108347 70601 108359 70635
rect 108301 70595 108359 70601
rect 105538 70564 105544 70576
rect 99708 70536 101352 70564
rect 102428 70536 105544 70564
rect 99708 70524 99714 70536
rect 101324 70508 101352 70536
rect 105538 70524 105544 70536
rect 105596 70524 105602 70576
rect 105630 70524 105636 70576
rect 105688 70564 105694 70576
rect 105817 70567 105875 70573
rect 105817 70564 105829 70567
rect 105688 70536 105829 70564
rect 105688 70524 105694 70536
rect 105817 70533 105829 70536
rect 105863 70533 105875 70567
rect 105817 70527 105875 70533
rect 105998 70524 106004 70576
rect 106056 70524 106062 70576
rect 98273 70499 98331 70505
rect 98273 70465 98285 70499
rect 98319 70465 98331 70499
rect 98273 70459 98331 70465
rect 98457 70499 98515 70505
rect 98457 70465 98469 70499
rect 98503 70465 98515 70499
rect 98457 70459 98515 70465
rect 97442 70388 97448 70440
rect 97500 70428 97506 70440
rect 97537 70431 97595 70437
rect 97537 70428 97549 70431
rect 97500 70400 97549 70428
rect 97500 70388 97506 70400
rect 97537 70397 97549 70400
rect 97583 70428 97595 70431
rect 97626 70428 97632 70440
rect 97583 70400 97632 70428
rect 97583 70397 97595 70400
rect 97537 70391 97595 70397
rect 97626 70388 97632 70400
rect 97684 70388 97690 70440
rect 97902 70388 97908 70440
rect 97960 70428 97966 70440
rect 98472 70428 98500 70459
rect 98546 70456 98552 70508
rect 98604 70496 98610 70508
rect 99285 70499 99343 70505
rect 98604 70468 99144 70496
rect 98604 70456 98610 70468
rect 97960 70400 98500 70428
rect 97960 70388 97966 70400
rect 96479 70332 97396 70360
rect 96479 70329 96491 70332
rect 96433 70323 96491 70329
rect 98086 70320 98092 70372
rect 98144 70320 98150 70372
rect 99116 70369 99144 70468
rect 99285 70465 99297 70499
rect 99331 70465 99343 70499
rect 99285 70459 99343 70465
rect 99190 70388 99196 70440
rect 99248 70428 99254 70440
rect 99300 70428 99328 70459
rect 99374 70456 99380 70508
rect 99432 70456 99438 70508
rect 99561 70499 99619 70505
rect 99561 70465 99573 70499
rect 99607 70465 99619 70499
rect 99561 70459 99619 70465
rect 99576 70428 99604 70459
rect 100202 70456 100208 70508
rect 100260 70456 100266 70508
rect 101306 70456 101312 70508
rect 101364 70496 101370 70508
rect 101953 70499 102011 70505
rect 101953 70496 101965 70499
rect 101364 70468 101965 70496
rect 101364 70456 101370 70468
rect 101953 70465 101965 70468
rect 101999 70496 102011 70499
rect 102134 70496 102140 70508
rect 101999 70468 102140 70496
rect 101999 70465 102011 70468
rect 101953 70459 102011 70465
rect 102134 70456 102140 70468
rect 102192 70456 102198 70508
rect 103793 70499 103851 70505
rect 103793 70465 103805 70499
rect 103839 70496 103851 70499
rect 103882 70496 103888 70508
rect 103839 70468 103888 70496
rect 103839 70465 103851 70468
rect 103793 70459 103851 70465
rect 103882 70456 103888 70468
rect 103940 70496 103946 70508
rect 105078 70496 105084 70508
rect 103940 70468 105084 70496
rect 103940 70456 103946 70468
rect 105078 70456 105084 70468
rect 105136 70496 105142 70508
rect 105173 70499 105231 70505
rect 105173 70496 105185 70499
rect 105136 70468 105185 70496
rect 105136 70456 105142 70468
rect 105173 70465 105185 70468
rect 105219 70465 105231 70499
rect 106093 70499 106151 70505
rect 106093 70496 106105 70499
rect 105173 70459 105231 70465
rect 105372 70468 106105 70496
rect 105372 70440 105400 70468
rect 106093 70465 106105 70468
rect 106139 70465 106151 70499
rect 106093 70459 106151 70465
rect 106274 70456 106280 70508
rect 106332 70456 106338 70508
rect 108209 70499 108267 70505
rect 108209 70465 108221 70499
rect 108255 70496 108267 70499
rect 108482 70496 108488 70508
rect 108255 70468 108488 70496
rect 108255 70465 108267 70468
rect 108209 70459 108267 70465
rect 108482 70456 108488 70468
rect 108540 70456 108546 70508
rect 99248 70400 99604 70428
rect 99248 70388 99254 70400
rect 101858 70388 101864 70440
rect 101916 70428 101922 70440
rect 102045 70431 102103 70437
rect 102045 70428 102057 70431
rect 101916 70400 102057 70428
rect 101916 70388 101922 70400
rect 102045 70397 102057 70400
rect 102091 70428 102103 70431
rect 103146 70428 103152 70440
rect 102091 70400 103152 70428
rect 102091 70397 102103 70400
rect 102045 70391 102103 70397
rect 103146 70388 103152 70400
rect 103204 70388 103210 70440
rect 103977 70431 104035 70437
rect 103977 70397 103989 70431
rect 104023 70428 104035 70431
rect 104986 70428 104992 70440
rect 104023 70400 104992 70428
rect 104023 70397 104035 70400
rect 103977 70391 104035 70397
rect 104986 70388 104992 70400
rect 105044 70428 105050 70440
rect 105265 70431 105323 70437
rect 105265 70428 105277 70431
rect 105044 70400 105277 70428
rect 105044 70388 105050 70400
rect 105265 70397 105277 70400
rect 105311 70397 105323 70431
rect 105265 70391 105323 70397
rect 105354 70388 105360 70440
rect 105412 70388 105418 70440
rect 105449 70431 105507 70437
rect 105449 70397 105461 70431
rect 105495 70428 105507 70431
rect 106292 70428 106320 70456
rect 107930 70428 107936 70440
rect 105495 70400 106320 70428
rect 106384 70400 107936 70428
rect 105495 70397 105507 70400
rect 105449 70391 105507 70397
rect 99101 70363 99159 70369
rect 99101 70329 99113 70363
rect 99147 70329 99159 70363
rect 99101 70323 99159 70329
rect 102318 70320 102324 70372
rect 102376 70320 102382 70372
rect 105538 70320 105544 70372
rect 105596 70360 105602 70372
rect 106384 70360 106412 70400
rect 107930 70388 107936 70400
rect 107988 70388 107994 70440
rect 105596 70332 106412 70360
rect 105596 70320 105602 70332
rect 93302 70252 93308 70304
rect 93360 70252 93366 70304
rect 99742 70252 99748 70304
rect 99800 70292 99806 70304
rect 100021 70295 100079 70301
rect 100021 70292 100033 70295
rect 99800 70264 100033 70292
rect 99800 70252 99806 70264
rect 100021 70261 100033 70264
rect 100067 70261 100079 70295
rect 100021 70255 100079 70261
rect 104989 70295 105047 70301
rect 104989 70261 105001 70295
rect 105035 70292 105047 70295
rect 105170 70292 105176 70304
rect 105035 70264 105176 70292
rect 105035 70261 105047 70264
rect 104989 70255 105047 70261
rect 105170 70252 105176 70264
rect 105228 70252 105234 70304
rect 105630 70252 105636 70304
rect 105688 70252 105694 70304
rect 1104 70202 108836 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 34934 70202
rect 34986 70150 34998 70202
rect 35050 70150 35062 70202
rect 35114 70150 35126 70202
rect 35178 70150 35190 70202
rect 35242 70150 65654 70202
rect 65706 70150 65718 70202
rect 65770 70150 65782 70202
rect 65834 70150 65846 70202
rect 65898 70150 65910 70202
rect 65962 70150 96374 70202
rect 96426 70150 96438 70202
rect 96490 70150 96502 70202
rect 96554 70150 96566 70202
rect 96618 70150 96630 70202
rect 96682 70150 108836 70202
rect 1104 70128 108836 70150
rect 31846 70048 31852 70100
rect 31904 70088 31910 70100
rect 32033 70091 32091 70097
rect 32033 70088 32045 70091
rect 31904 70060 32045 70088
rect 31904 70048 31910 70060
rect 32033 70057 32045 70060
rect 32079 70088 32091 70091
rect 32217 70091 32275 70097
rect 32217 70088 32229 70091
rect 32079 70060 32229 70088
rect 32079 70057 32091 70060
rect 32033 70051 32091 70057
rect 32217 70057 32229 70060
rect 32263 70057 32275 70091
rect 32217 70051 32275 70057
rect 35526 70048 35532 70100
rect 35584 70088 35590 70100
rect 35584 70060 37136 70088
rect 35584 70048 35590 70060
rect 32950 69980 32956 70032
rect 33008 70020 33014 70032
rect 35713 70023 35771 70029
rect 35713 70020 35725 70023
rect 33008 69992 35725 70020
rect 33008 69980 33014 69992
rect 35713 69989 35725 69992
rect 35759 69989 35771 70023
rect 35713 69983 35771 69989
rect 37108 69961 37136 70060
rect 72878 70048 72884 70100
rect 72936 70088 72942 70100
rect 73341 70091 73399 70097
rect 73341 70088 73353 70091
rect 72936 70060 73353 70088
rect 72936 70048 72942 70060
rect 73341 70057 73353 70060
rect 73387 70057 73399 70091
rect 73341 70051 73399 70057
rect 75089 70091 75147 70097
rect 75089 70057 75101 70091
rect 75135 70088 75147 70091
rect 75135 70060 80560 70088
rect 75135 70057 75147 70060
rect 75089 70051 75147 70057
rect 37093 69955 37151 69961
rect 37093 69921 37105 69955
rect 37139 69952 37151 69955
rect 38654 69952 38660 69964
rect 37139 69924 38660 69952
rect 37139 69921 37151 69924
rect 37093 69915 37151 69921
rect 38654 69912 38660 69924
rect 38712 69912 38718 69964
rect 73356 69952 73384 70051
rect 73709 69955 73767 69961
rect 73709 69952 73721 69955
rect 73356 69924 73721 69952
rect 73709 69921 73721 69924
rect 73755 69921 73767 69955
rect 73709 69915 73767 69921
rect 79137 69955 79195 69961
rect 79137 69921 79149 69955
rect 79183 69952 79195 69955
rect 79502 69952 79508 69964
rect 79183 69924 79508 69952
rect 79183 69921 79195 69924
rect 79137 69915 79195 69921
rect 77573 69887 77631 69893
rect 77573 69853 77585 69887
rect 77619 69884 77631 69887
rect 79152 69884 79180 69915
rect 79502 69912 79508 69924
rect 79560 69912 79566 69964
rect 80532 69952 80560 70060
rect 81158 70048 81164 70100
rect 81216 70048 81222 70100
rect 89714 70048 89720 70100
rect 89772 70088 89778 70100
rect 90634 70088 90640 70100
rect 89772 70060 90640 70088
rect 89772 70048 89778 70060
rect 90634 70048 90640 70060
rect 90692 70088 90698 70100
rect 91557 70091 91615 70097
rect 91557 70088 91569 70091
rect 90692 70060 91569 70088
rect 90692 70048 90698 70060
rect 91557 70057 91569 70060
rect 91603 70057 91615 70091
rect 91557 70051 91615 70057
rect 97534 70048 97540 70100
rect 97592 70088 97598 70100
rect 97721 70091 97779 70097
rect 97721 70088 97733 70091
rect 97592 70060 97733 70088
rect 97592 70048 97598 70060
rect 97721 70057 97733 70060
rect 97767 70057 97779 70091
rect 97721 70051 97779 70057
rect 98457 70091 98515 70097
rect 98457 70057 98469 70091
rect 98503 70088 98515 70091
rect 99190 70088 99196 70100
rect 98503 70060 99196 70088
rect 98503 70057 98515 70060
rect 98457 70051 98515 70057
rect 99190 70048 99196 70060
rect 99248 70048 99254 70100
rect 99285 70091 99343 70097
rect 99285 70057 99297 70091
rect 99331 70088 99343 70091
rect 99374 70088 99380 70100
rect 99331 70060 99380 70088
rect 99331 70057 99343 70060
rect 99285 70051 99343 70057
rect 99374 70048 99380 70060
rect 99432 70048 99438 70100
rect 99834 70048 99840 70100
rect 99892 70088 99898 70100
rect 99929 70091 99987 70097
rect 99929 70088 99941 70091
rect 99892 70060 99941 70088
rect 99892 70048 99898 70060
rect 99929 70057 99941 70060
rect 99975 70057 99987 70091
rect 99929 70051 99987 70057
rect 100202 70048 100208 70100
rect 100260 70088 100266 70100
rect 100297 70091 100355 70097
rect 100297 70088 100309 70091
rect 100260 70060 100309 70088
rect 100260 70048 100266 70060
rect 100297 70057 100309 70060
rect 100343 70057 100355 70091
rect 101950 70088 101956 70100
rect 100297 70051 100355 70057
rect 100772 70060 101956 70088
rect 80885 70023 80943 70029
rect 80885 69989 80897 70023
rect 80931 70020 80943 70023
rect 88334 70020 88340 70032
rect 80931 69992 88340 70020
rect 80931 69989 80943 69992
rect 80885 69983 80943 69989
rect 88334 69980 88340 69992
rect 88392 69980 88398 70032
rect 90358 69980 90364 70032
rect 90416 70020 90422 70032
rect 91373 70023 91431 70029
rect 91373 70020 91385 70023
rect 90416 69992 91385 70020
rect 90416 69980 90422 69992
rect 91373 69989 91385 69992
rect 91419 69989 91431 70023
rect 91373 69983 91431 69989
rect 95234 69980 95240 70032
rect 95292 70020 95298 70032
rect 96341 70023 96399 70029
rect 96341 70020 96353 70023
rect 95292 69992 96353 70020
rect 95292 69980 95298 69992
rect 96341 69989 96353 69992
rect 96387 69989 96399 70023
rect 96341 69983 96399 69989
rect 97077 70023 97135 70029
rect 97077 69989 97089 70023
rect 97123 70020 97135 70023
rect 97258 70020 97264 70032
rect 97123 69992 97264 70020
rect 97123 69989 97135 69992
rect 97077 69983 97135 69989
rect 97258 69980 97264 69992
rect 97316 70020 97322 70032
rect 97902 70020 97908 70032
rect 97316 69992 97908 70020
rect 97316 69980 97322 69992
rect 97902 69980 97908 69992
rect 97960 69980 97966 70032
rect 98638 69980 98644 70032
rect 98696 69980 98702 70032
rect 100772 70020 100800 70060
rect 101950 70048 101956 70060
rect 102008 70048 102014 70100
rect 105722 70048 105728 70100
rect 105780 70088 105786 70100
rect 108301 70091 108359 70097
rect 108301 70088 108313 70091
rect 105780 70060 108313 70088
rect 105780 70048 105786 70060
rect 108301 70057 108313 70060
rect 108347 70057 108359 70091
rect 108301 70051 108359 70057
rect 99852 69992 100800 70020
rect 100849 70023 100907 70029
rect 83090 69952 83096 69964
rect 80532 69924 83096 69952
rect 83090 69912 83096 69924
rect 83148 69912 83154 69964
rect 85390 69912 85396 69964
rect 85448 69952 85454 69964
rect 89533 69955 89591 69961
rect 89533 69952 89545 69955
rect 85448 69924 89545 69952
rect 85448 69912 85454 69924
rect 89533 69921 89545 69924
rect 89579 69952 89591 69955
rect 90085 69955 90143 69961
rect 90085 69952 90097 69955
rect 89579 69924 90097 69952
rect 89579 69921 89591 69924
rect 89533 69915 89591 69921
rect 90085 69921 90097 69924
rect 90131 69952 90143 69955
rect 90131 69924 90496 69952
rect 90131 69921 90143 69924
rect 90085 69915 90143 69921
rect 77619 69856 79180 69884
rect 77619 69853 77631 69856
rect 77573 69847 77631 69853
rect 79318 69844 79324 69896
rect 79376 69844 79382 69896
rect 86770 69884 86776 69896
rect 79704 69856 86776 69884
rect 36848 69819 36906 69825
rect 36848 69785 36860 69819
rect 36894 69816 36906 69819
rect 45094 69816 45100 69828
rect 36894 69788 45100 69816
rect 36894 69785 36906 69788
rect 36848 69779 36906 69785
rect 45094 69776 45100 69788
rect 45152 69776 45158 69828
rect 77846 69825 77852 69828
rect 73954 69819 74012 69825
rect 73954 69816 73966 69819
rect 73540 69788 73966 69816
rect 30653 69751 30711 69757
rect 30653 69717 30665 69751
rect 30699 69748 30711 69751
rect 31662 69748 31668 69760
rect 30699 69720 31668 69748
rect 30699 69717 30711 69720
rect 30653 69711 30711 69717
rect 31662 69708 31668 69720
rect 31720 69708 31726 69760
rect 66714 69708 66720 69760
rect 66772 69708 66778 69760
rect 72418 69708 72424 69760
rect 72476 69748 72482 69760
rect 73540 69757 73568 69788
rect 73954 69785 73966 69788
rect 74000 69785 74012 69819
rect 73954 69779 74012 69785
rect 77481 69819 77539 69825
rect 77481 69785 77493 69819
rect 77527 69816 77539 69819
rect 77840 69816 77852 69825
rect 77527 69788 77852 69816
rect 77527 69785 77539 69788
rect 77481 69779 77539 69785
rect 77840 69779 77852 69788
rect 77846 69776 77852 69779
rect 77904 69776 77910 69828
rect 79704 69816 79732 69856
rect 86770 69844 86776 69856
rect 86828 69844 86834 69896
rect 90358 69844 90364 69896
rect 90416 69844 90422 69896
rect 90468 69893 90496 69924
rect 90634 69912 90640 69964
rect 90692 69912 90698 69964
rect 95053 69955 95111 69961
rect 95053 69921 95065 69955
rect 95099 69952 95111 69955
rect 95694 69952 95700 69964
rect 95099 69924 95700 69952
rect 95099 69921 95111 69924
rect 95053 69915 95111 69921
rect 95694 69912 95700 69924
rect 95752 69912 95758 69964
rect 96801 69955 96859 69961
rect 96801 69921 96813 69955
rect 96847 69952 96859 69955
rect 97810 69952 97816 69964
rect 96847 69924 97816 69952
rect 96847 69921 96859 69924
rect 96801 69915 96859 69921
rect 97810 69912 97816 69924
rect 97868 69912 97874 69964
rect 98656 69952 98684 69980
rect 99852 69961 99880 69992
rect 100849 69989 100861 70023
rect 100895 69989 100907 70023
rect 100849 69983 100907 69989
rect 97920 69924 98684 69952
rect 99837 69955 99895 69961
rect 90453 69887 90511 69893
rect 90453 69853 90465 69887
rect 90499 69884 90511 69887
rect 91005 69887 91063 69893
rect 91005 69884 91017 69887
rect 90499 69856 91017 69884
rect 90499 69853 90511 69856
rect 90453 69847 90511 69853
rect 91005 69853 91017 69856
rect 91051 69853 91063 69887
rect 91005 69847 91063 69853
rect 94041 69887 94099 69893
rect 94041 69853 94053 69887
rect 94087 69884 94099 69887
rect 94314 69884 94320 69896
rect 94087 69856 94320 69884
rect 94087 69853 94099 69856
rect 94041 69847 94099 69853
rect 94314 69844 94320 69856
rect 94372 69844 94378 69896
rect 94685 69887 94743 69893
rect 94685 69853 94697 69887
rect 94731 69884 94743 69887
rect 94866 69884 94872 69896
rect 94731 69856 94872 69884
rect 94731 69853 94743 69856
rect 94685 69847 94743 69853
rect 94866 69844 94872 69856
rect 94924 69884 94930 69896
rect 95145 69887 95203 69893
rect 95145 69884 95157 69887
rect 94924 69856 95157 69884
rect 94924 69844 94930 69856
rect 95145 69853 95157 69856
rect 95191 69853 95203 69887
rect 95145 69847 95203 69853
rect 96065 69887 96123 69893
rect 96065 69853 96077 69887
rect 96111 69884 96123 69887
rect 96154 69884 96160 69896
rect 96111 69856 96160 69884
rect 96111 69853 96123 69856
rect 96065 69847 96123 69853
rect 96154 69844 96160 69856
rect 96212 69844 96218 69896
rect 96709 69887 96767 69893
rect 96709 69853 96721 69887
rect 96755 69884 96767 69887
rect 97534 69884 97540 69896
rect 96755 69856 97540 69884
rect 96755 69853 96767 69856
rect 96709 69847 96767 69853
rect 97534 69844 97540 69856
rect 97592 69844 97598 69896
rect 97920 69893 97948 69924
rect 99837 69921 99849 69955
rect 99883 69921 99895 69955
rect 100864 69952 100892 69983
rect 99837 69915 99895 69921
rect 100220 69924 100892 69952
rect 97721 69887 97779 69893
rect 97721 69853 97733 69887
rect 97767 69853 97779 69887
rect 97721 69847 97779 69853
rect 97905 69887 97963 69893
rect 97905 69853 97917 69887
rect 97951 69853 97963 69887
rect 97905 69847 97963 69853
rect 98457 69887 98515 69893
rect 98457 69853 98469 69887
rect 98503 69853 98515 69887
rect 98457 69847 98515 69853
rect 98641 69887 98699 69893
rect 98641 69853 98653 69887
rect 98687 69884 98699 69887
rect 99006 69884 99012 69896
rect 98687 69856 99012 69884
rect 98687 69853 98699 69856
rect 98641 69847 98699 69853
rect 78968 69788 79732 69816
rect 79772 69819 79830 69825
rect 78968 69757 78996 69788
rect 79772 69785 79784 69819
rect 79818 69785 79830 69819
rect 79772 69779 79830 69785
rect 73525 69751 73583 69757
rect 73525 69748 73537 69751
rect 72476 69720 73537 69748
rect 72476 69708 72482 69720
rect 73525 69717 73537 69720
rect 73571 69717 73583 69751
rect 73525 69711 73583 69717
rect 78953 69751 79011 69757
rect 78953 69717 78965 69751
rect 78999 69717 79011 69751
rect 78953 69711 79011 69717
rect 79318 69708 79324 69760
rect 79376 69748 79382 69760
rect 79796 69748 79824 69779
rect 92474 69776 92480 69828
rect 92532 69816 92538 69828
rect 93762 69816 93768 69828
rect 92532 69788 93768 69816
rect 92532 69776 92538 69788
rect 93762 69776 93768 69788
rect 93820 69816 93826 69828
rect 94225 69819 94283 69825
rect 94225 69816 94237 69819
rect 93820 69788 94237 69816
rect 93820 69776 93826 69788
rect 94225 69785 94237 69788
rect 94271 69785 94283 69819
rect 94225 69779 94283 69785
rect 94409 69819 94467 69825
rect 94409 69785 94421 69819
rect 94455 69816 94467 69819
rect 96341 69819 96399 69825
rect 94455 69788 96292 69816
rect 94455 69785 94467 69788
rect 94409 69779 94467 69785
rect 79376 69720 79824 69748
rect 79376 69708 79382 69720
rect 94774 69708 94780 69760
rect 94832 69708 94838 69760
rect 96062 69708 96068 69760
rect 96120 69748 96126 69760
rect 96157 69751 96215 69757
rect 96157 69748 96169 69751
rect 96120 69720 96169 69748
rect 96120 69708 96126 69720
rect 96157 69717 96169 69720
rect 96203 69717 96215 69751
rect 96264 69748 96292 69788
rect 96341 69785 96353 69819
rect 96387 69816 96399 69819
rect 97442 69816 97448 69828
rect 96387 69788 97448 69816
rect 96387 69785 96399 69788
rect 96341 69779 96399 69785
rect 97442 69776 97448 69788
rect 97500 69776 97506 69828
rect 97736 69816 97764 69847
rect 98178 69816 98184 69828
rect 97736 69788 98184 69816
rect 98178 69776 98184 69788
rect 98236 69776 98242 69828
rect 98472 69816 98500 69847
rect 99006 69844 99012 69856
rect 99064 69844 99070 69896
rect 99101 69887 99159 69893
rect 99101 69853 99113 69887
rect 99147 69884 99159 69887
rect 99466 69884 99472 69896
rect 99147 69856 99472 69884
rect 99147 69853 99159 69856
rect 99101 69847 99159 69853
rect 99116 69816 99144 69847
rect 99466 69844 99472 69856
rect 99524 69844 99530 69896
rect 99742 69844 99748 69896
rect 99800 69844 99806 69896
rect 100220 69893 100248 69924
rect 101398 69912 101404 69964
rect 101456 69952 101462 69964
rect 101456 69924 101628 69952
rect 101456 69912 101462 69924
rect 100205 69887 100263 69893
rect 100205 69853 100217 69887
rect 100251 69853 100263 69887
rect 100205 69847 100263 69853
rect 100389 69887 100447 69893
rect 100389 69853 100401 69887
rect 100435 69853 100447 69887
rect 100389 69847 100447 69853
rect 98472 69788 99144 69816
rect 100404 69816 100432 69847
rect 100478 69844 100484 69896
rect 100536 69844 100542 69896
rect 100846 69884 100852 69896
rect 100588 69856 100852 69884
rect 100588 69816 100616 69856
rect 100846 69844 100852 69856
rect 100904 69844 100910 69896
rect 100938 69844 100944 69896
rect 100996 69844 101002 69896
rect 101306 69844 101312 69896
rect 101364 69844 101370 69896
rect 101490 69844 101496 69896
rect 101548 69844 101554 69896
rect 101600 69884 101628 69924
rect 101950 69912 101956 69964
rect 102008 69912 102014 69964
rect 103606 69912 103612 69964
rect 103664 69952 103670 69964
rect 104621 69955 104679 69961
rect 104621 69952 104633 69955
rect 103664 69924 104633 69952
rect 103664 69912 103670 69924
rect 104621 69921 104633 69924
rect 104667 69921 104679 69955
rect 104621 69915 104679 69921
rect 104986 69912 104992 69964
rect 105044 69952 105050 69964
rect 105044 69924 105216 69952
rect 105044 69912 105050 69924
rect 101861 69887 101919 69893
rect 101861 69884 101873 69887
rect 101600 69856 101873 69884
rect 101861 69853 101873 69856
rect 101907 69853 101919 69887
rect 101861 69847 101919 69853
rect 104437 69887 104495 69893
rect 104437 69853 104449 69887
rect 104483 69884 104495 69887
rect 104894 69884 104900 69896
rect 104483 69856 104900 69884
rect 104483 69853 104495 69856
rect 104437 69847 104495 69853
rect 104894 69844 104900 69856
rect 104952 69844 104958 69896
rect 105078 69844 105084 69896
rect 105136 69844 105142 69896
rect 105188 69893 105216 69924
rect 105173 69887 105231 69893
rect 105173 69853 105185 69887
rect 105219 69853 105231 69887
rect 105173 69847 105231 69853
rect 105262 69844 105268 69896
rect 105320 69844 105326 69896
rect 108209 69887 108267 69893
rect 108209 69853 108221 69887
rect 108255 69884 108267 69887
rect 108482 69884 108488 69896
rect 108255 69856 108488 69884
rect 108255 69853 108267 69856
rect 108209 69847 108267 69853
rect 108482 69844 108488 69856
rect 108540 69844 108546 69896
rect 100404 69788 100616 69816
rect 100754 69776 100760 69828
rect 100812 69816 100818 69828
rect 101125 69819 101183 69825
rect 101125 69816 101137 69819
rect 100812 69788 101137 69816
rect 100812 69776 100818 69788
rect 101125 69785 101137 69788
rect 101171 69816 101183 69819
rect 101674 69816 101680 69828
rect 101171 69788 101680 69816
rect 101171 69785 101183 69788
rect 101125 69779 101183 69785
rect 101674 69776 101680 69788
rect 101732 69776 101738 69828
rect 104529 69819 104587 69825
rect 104529 69785 104541 69819
rect 104575 69816 104587 69819
rect 105630 69816 105636 69828
rect 104575 69788 105636 69816
rect 104575 69785 104587 69788
rect 104529 69779 104587 69785
rect 105630 69776 105636 69788
rect 105688 69776 105694 69828
rect 96798 69748 96804 69760
rect 96264 69720 96804 69748
rect 96157 69711 96215 69717
rect 96798 69708 96804 69720
rect 96856 69708 96862 69760
rect 99561 69751 99619 69757
rect 99561 69717 99573 69751
rect 99607 69748 99619 69751
rect 99650 69748 99656 69760
rect 99607 69720 99656 69748
rect 99607 69717 99619 69720
rect 99561 69711 99619 69717
rect 99650 69708 99656 69720
rect 99708 69708 99714 69760
rect 100018 69708 100024 69760
rect 100076 69708 100082 69760
rect 100110 69708 100116 69760
rect 100168 69708 100174 69760
rect 100665 69751 100723 69757
rect 100665 69717 100677 69751
rect 100711 69748 100723 69751
rect 100938 69748 100944 69760
rect 100711 69720 100944 69748
rect 100711 69717 100723 69720
rect 100665 69711 100723 69717
rect 100938 69708 100944 69720
rect 100996 69748 101002 69760
rect 101309 69751 101367 69757
rect 101309 69748 101321 69751
rect 100996 69720 101321 69748
rect 100996 69708 101002 69720
rect 101309 69717 101321 69720
rect 101355 69717 101367 69751
rect 101309 69711 101367 69717
rect 102226 69708 102232 69760
rect 102284 69708 102290 69760
rect 103330 69708 103336 69760
rect 103388 69748 103394 69760
rect 104069 69751 104127 69757
rect 104069 69748 104081 69751
rect 103388 69720 104081 69748
rect 103388 69708 103394 69720
rect 104069 69717 104081 69720
rect 104115 69717 104127 69751
rect 104069 69711 104127 69717
rect 104894 69708 104900 69760
rect 104952 69708 104958 69760
rect 1104 69658 108836 69680
rect 1104 69606 4874 69658
rect 4926 69606 4938 69658
rect 4990 69606 5002 69658
rect 5054 69606 5066 69658
rect 5118 69606 5130 69658
rect 5182 69606 35594 69658
rect 35646 69606 35658 69658
rect 35710 69606 35722 69658
rect 35774 69606 35786 69658
rect 35838 69606 35850 69658
rect 35902 69606 66314 69658
rect 66366 69606 66378 69658
rect 66430 69606 66442 69658
rect 66494 69606 66506 69658
rect 66558 69606 66570 69658
rect 66622 69606 97034 69658
rect 97086 69606 97098 69658
rect 97150 69606 97162 69658
rect 97214 69606 97226 69658
rect 97278 69606 97290 69658
rect 97342 69606 108836 69658
rect 1104 69584 108836 69606
rect 42426 69504 42432 69556
rect 42484 69504 42490 69556
rect 62853 69547 62911 69553
rect 62853 69513 62865 69547
rect 62899 69544 62911 69547
rect 62899 69516 67312 69544
rect 62899 69513 62911 69516
rect 62853 69507 62911 69513
rect 63129 69479 63187 69485
rect 63129 69476 63141 69479
rect 61488 69448 63141 69476
rect 43553 69411 43611 69417
rect 43553 69377 43565 69411
rect 43599 69408 43611 69411
rect 43714 69408 43720 69420
rect 43599 69380 43720 69408
rect 43599 69377 43611 69380
rect 43553 69371 43611 69377
rect 43714 69368 43720 69380
rect 43772 69368 43778 69420
rect 61488 69417 61516 69448
rect 63129 69445 63141 69448
rect 63175 69476 63187 69479
rect 67174 69476 67180 69488
rect 63175 69448 67180 69476
rect 63175 69445 63187 69448
rect 63129 69439 63187 69445
rect 66640 69417 66668 69448
rect 67174 69436 67180 69448
rect 67232 69436 67238 69488
rect 61473 69411 61531 69417
rect 61473 69377 61485 69411
rect 61519 69377 61531 69411
rect 61729 69411 61787 69417
rect 61729 69408 61741 69411
rect 61473 69371 61531 69377
rect 61580 69380 61741 69408
rect 43809 69343 43867 69349
rect 43809 69309 43821 69343
rect 43855 69309 43867 69343
rect 61580 69340 61608 69380
rect 61729 69377 61741 69380
rect 61775 69377 61787 69411
rect 61729 69371 61787 69377
rect 66625 69411 66683 69417
rect 66625 69377 66637 69411
rect 66671 69377 66683 69411
rect 66625 69371 66683 69377
rect 66714 69368 66720 69420
rect 66772 69408 66778 69420
rect 66881 69411 66939 69417
rect 66881 69408 66893 69411
rect 66772 69380 66893 69408
rect 66772 69368 66778 69380
rect 66881 69377 66893 69380
rect 66927 69377 66939 69411
rect 67284 69408 67312 69516
rect 67358 69504 67364 69556
rect 67416 69544 67422 69556
rect 68281 69547 68339 69553
rect 68281 69544 68293 69547
rect 67416 69516 68293 69544
rect 67416 69504 67422 69516
rect 68281 69513 68293 69516
rect 68327 69544 68339 69547
rect 69106 69544 69112 69556
rect 68327 69516 69112 69544
rect 68327 69513 68339 69516
rect 68281 69507 68339 69513
rect 69106 69504 69112 69516
rect 69164 69504 69170 69556
rect 79318 69504 79324 69556
rect 79376 69544 79382 69556
rect 79505 69547 79563 69553
rect 79505 69544 79517 69547
rect 79376 69516 79517 69544
rect 79376 69504 79382 69516
rect 79505 69513 79517 69516
rect 79551 69513 79563 69547
rect 79505 69507 79563 69513
rect 88794 69504 88800 69556
rect 88852 69504 88858 69556
rect 92093 69547 92151 69553
rect 89180 69516 92060 69544
rect 69014 69408 69020 69420
rect 67284 69380 69020 69408
rect 66881 69371 66939 69377
rect 69014 69368 69020 69380
rect 69072 69368 69078 69420
rect 86310 69368 86316 69420
rect 86368 69408 86374 69420
rect 89180 69417 89208 69516
rect 89533 69479 89591 69485
rect 89533 69445 89545 69479
rect 89579 69476 89591 69479
rect 89579 69448 90390 69476
rect 89579 69445 89591 69448
rect 89533 69439 89591 69445
rect 91554 69436 91560 69488
rect 91612 69436 91618 69488
rect 89165 69411 89223 69417
rect 89165 69408 89177 69411
rect 86368 69380 89177 69408
rect 86368 69368 86374 69380
rect 89165 69377 89177 69380
rect 89211 69377 89223 69411
rect 89165 69371 89223 69377
rect 89441 69411 89499 69417
rect 89441 69377 89453 69411
rect 89487 69408 89499 69411
rect 89714 69408 89720 69420
rect 89487 69380 89720 69408
rect 89487 69377 89499 69380
rect 89441 69371 89499 69377
rect 89714 69368 89720 69380
rect 89772 69368 89778 69420
rect 91830 69368 91836 69420
rect 91888 69368 91894 69420
rect 92032 69408 92060 69516
rect 92093 69513 92105 69547
rect 92139 69544 92151 69547
rect 92934 69544 92940 69556
rect 92139 69516 92940 69544
rect 92139 69513 92151 69516
rect 92093 69507 92151 69513
rect 92934 69504 92940 69516
rect 92992 69504 92998 69556
rect 97810 69504 97816 69556
rect 97868 69504 97874 69556
rect 97997 69547 98055 69553
rect 97997 69513 98009 69547
rect 98043 69544 98055 69547
rect 99466 69544 99472 69556
rect 98043 69516 99472 69544
rect 98043 69513 98055 69516
rect 97997 69507 98055 69513
rect 99466 69504 99472 69516
rect 99524 69504 99530 69556
rect 100297 69547 100355 69553
rect 100297 69513 100309 69547
rect 100343 69544 100355 69547
rect 100938 69544 100944 69556
rect 100343 69516 100944 69544
rect 100343 69513 100355 69516
rect 100297 69507 100355 69513
rect 100938 69504 100944 69516
rect 100996 69504 101002 69556
rect 102597 69547 102655 69553
rect 102597 69513 102609 69547
rect 102643 69513 102655 69547
rect 102597 69507 102655 69513
rect 92290 69436 92296 69488
rect 92348 69436 92354 69488
rect 99558 69476 99564 69488
rect 99268 69448 99564 69476
rect 92474 69408 92480 69420
rect 92032 69380 92480 69408
rect 92474 69368 92480 69380
rect 92532 69368 92538 69420
rect 92569 69411 92627 69417
rect 92569 69377 92581 69411
rect 92615 69408 92627 69411
rect 93026 69408 93032 69420
rect 92615 69380 93032 69408
rect 92615 69377 92627 69380
rect 92569 69371 92627 69377
rect 93026 69368 93032 69380
rect 93084 69368 93090 69420
rect 97994 69411 98052 69417
rect 97994 69377 98006 69411
rect 98040 69408 98052 69411
rect 98270 69408 98276 69420
rect 98040 69380 98276 69408
rect 98040 69377 98052 69380
rect 97994 69371 98052 69377
rect 98270 69368 98276 69380
rect 98328 69368 98334 69420
rect 98365 69411 98423 69417
rect 98365 69377 98377 69411
rect 98411 69408 98423 69411
rect 98730 69408 98736 69420
rect 98411 69380 98736 69408
rect 98411 69377 98423 69380
rect 98365 69371 98423 69377
rect 98730 69368 98736 69380
rect 98788 69368 98794 69420
rect 98824 69411 98882 69417
rect 98824 69377 98836 69411
rect 98870 69377 98882 69411
rect 98824 69371 98882 69377
rect 43809 69303 43867 69309
rect 61488 69312 61608 69340
rect 42168 69244 42932 69272
rect 42168 69216 42196 69244
rect 42150 69164 42156 69216
rect 42208 69164 42214 69216
rect 42904 69204 42932 69244
rect 43824 69216 43852 69303
rect 61488 69216 61516 69312
rect 66438 69300 66444 69352
rect 66496 69340 66502 69352
rect 66732 69340 66760 69368
rect 66496 69312 66760 69340
rect 66496 69300 66502 69312
rect 89070 69300 89076 69352
rect 89128 69300 89134 69352
rect 89809 69343 89867 69349
rect 89809 69309 89821 69343
rect 89855 69340 89867 69343
rect 91848 69340 91876 69368
rect 92845 69343 92903 69349
rect 92845 69340 92857 69343
rect 89855 69312 91784 69340
rect 91848 69312 92857 69340
rect 89855 69309 89867 69312
rect 89809 69303 89867 69309
rect 91756 69272 91784 69312
rect 92845 69309 92857 69312
rect 92891 69309 92903 69343
rect 92845 69303 92903 69309
rect 94958 69300 94964 69352
rect 95016 69340 95022 69352
rect 95878 69340 95884 69352
rect 95016 69312 95884 69340
rect 95016 69300 95022 69312
rect 95878 69300 95884 69312
rect 95936 69300 95942 69352
rect 98457 69343 98515 69349
rect 98457 69309 98469 69343
rect 98503 69340 98515 69343
rect 98549 69343 98607 69349
rect 98549 69340 98561 69343
rect 98503 69312 98561 69340
rect 98503 69309 98515 69312
rect 98457 69303 98515 69309
rect 98549 69309 98561 69312
rect 98595 69309 98607 69343
rect 98840 69340 98868 69371
rect 98914 69368 98920 69420
rect 98972 69368 98978 69420
rect 99098 69368 99104 69420
rect 99156 69368 99162 69420
rect 99268 69417 99296 69448
rect 99558 69436 99564 69448
rect 99616 69436 99622 69488
rect 100481 69479 100539 69485
rect 100481 69445 100493 69479
rect 100527 69476 100539 69479
rect 100846 69476 100852 69488
rect 100527 69448 100852 69476
rect 100527 69445 100539 69448
rect 100481 69439 100539 69445
rect 100846 69436 100852 69448
rect 100904 69476 100910 69488
rect 102612 69476 102640 69507
rect 100904 69448 102640 69476
rect 100904 69436 100910 69448
rect 99268 69411 99343 69417
rect 99268 69380 99297 69411
rect 99285 69377 99297 69380
rect 99331 69377 99343 69411
rect 99285 69371 99343 69377
rect 99374 69368 99380 69420
rect 99432 69408 99438 69420
rect 99469 69411 99527 69417
rect 99469 69408 99481 69411
rect 99432 69380 99481 69408
rect 99432 69368 99438 69380
rect 99469 69377 99481 69380
rect 99515 69377 99527 69411
rect 99469 69371 99527 69377
rect 99484 69340 99512 69371
rect 99650 69368 99656 69420
rect 99708 69368 99714 69420
rect 99742 69368 99748 69420
rect 99800 69408 99806 69420
rect 99929 69411 99987 69417
rect 99929 69408 99941 69411
rect 99800 69380 99941 69408
rect 99800 69368 99806 69380
rect 99929 69377 99941 69380
rect 99975 69377 99987 69411
rect 99929 69371 99987 69377
rect 100205 69411 100263 69417
rect 100205 69377 100217 69411
rect 100251 69408 100263 69411
rect 100754 69408 100760 69420
rect 100251 69380 100760 69408
rect 100251 69377 100263 69380
rect 100205 69371 100263 69377
rect 100754 69368 100760 69380
rect 100812 69368 100818 69420
rect 101490 69368 101496 69420
rect 101548 69408 101554 69420
rect 101876 69417 101904 69448
rect 101677 69411 101735 69417
rect 101677 69408 101689 69411
rect 101548 69380 101689 69408
rect 101548 69368 101554 69380
rect 101677 69377 101689 69380
rect 101723 69377 101735 69411
rect 101677 69371 101735 69377
rect 101861 69411 101919 69417
rect 101861 69377 101873 69411
rect 101907 69377 101919 69411
rect 101861 69371 101919 69377
rect 100846 69340 100852 69352
rect 98840 69312 99374 69340
rect 99484 69312 100852 69340
rect 98549 69303 98607 69309
rect 99346 69272 99374 69312
rect 100846 69300 100852 69312
rect 100904 69300 100910 69352
rect 101692 69340 101720 69371
rect 102318 69368 102324 69420
rect 102376 69408 102382 69420
rect 102597 69411 102655 69417
rect 102597 69408 102609 69411
rect 102376 69380 102609 69408
rect 102376 69368 102382 69380
rect 102597 69377 102609 69380
rect 102643 69408 102655 69411
rect 103238 69408 103244 69420
rect 102643 69380 103244 69408
rect 102643 69377 102655 69380
rect 102597 69371 102655 69377
rect 103238 69368 103244 69380
rect 103296 69368 103302 69420
rect 103330 69368 103336 69420
rect 103388 69368 103394 69420
rect 103514 69368 103520 69420
rect 103572 69408 103578 69420
rect 103793 69411 103851 69417
rect 103793 69408 103805 69411
rect 103572 69380 103805 69408
rect 103572 69368 103578 69380
rect 103793 69377 103805 69380
rect 103839 69377 103851 69411
rect 103793 69371 103851 69377
rect 103977 69411 104035 69417
rect 103977 69377 103989 69411
rect 104023 69377 104035 69411
rect 103977 69371 104035 69377
rect 102042 69340 102048 69352
rect 101692 69312 102048 69340
rect 102042 69300 102048 69312
rect 102100 69300 102106 69352
rect 102410 69300 102416 69352
rect 102468 69300 102474 69352
rect 102962 69300 102968 69352
rect 103020 69300 103026 69352
rect 103348 69340 103376 69368
rect 103992 69340 104020 69371
rect 104618 69368 104624 69420
rect 104676 69408 104682 69420
rect 104805 69411 104863 69417
rect 104805 69408 104817 69411
rect 104676 69380 104817 69408
rect 104676 69368 104682 69380
rect 104805 69377 104817 69380
rect 104851 69377 104863 69411
rect 104805 69371 104863 69377
rect 104986 69368 104992 69420
rect 105044 69368 105050 69420
rect 103348 69312 104020 69340
rect 99561 69275 99619 69281
rect 99561 69272 99573 69275
rect 91756 69244 92796 69272
rect 99346 69244 99573 69272
rect 92768 69216 92796 69244
rect 99561 69241 99573 69244
rect 99607 69241 99619 69275
rect 99561 69235 99619 69241
rect 43806 69204 43812 69216
rect 42904 69176 43812 69204
rect 43806 69164 43812 69176
rect 43864 69164 43870 69216
rect 61381 69207 61439 69213
rect 61381 69173 61393 69207
rect 61427 69204 61439 69207
rect 61470 69204 61476 69216
rect 61427 69176 61476 69204
rect 61427 69173 61439 69176
rect 61381 69167 61439 69173
rect 61470 69164 61476 69176
rect 61528 69164 61534 69216
rect 68005 69207 68063 69213
rect 68005 69173 68017 69207
rect 68051 69204 68063 69207
rect 74534 69204 74540 69216
rect 68051 69176 74540 69204
rect 68051 69173 68063 69176
rect 68005 69167 68063 69173
rect 74534 69164 74540 69176
rect 74592 69164 74598 69216
rect 91738 69164 91744 69216
rect 91796 69204 91802 69216
rect 91925 69207 91983 69213
rect 91925 69204 91937 69207
rect 91796 69176 91937 69204
rect 91796 69164 91802 69176
rect 91925 69173 91937 69176
rect 91971 69173 91983 69207
rect 91925 69167 91983 69173
rect 92109 69207 92167 69213
rect 92109 69173 92121 69207
rect 92155 69204 92167 69207
rect 92477 69207 92535 69213
rect 92477 69204 92489 69207
rect 92155 69176 92489 69204
rect 92155 69173 92167 69176
rect 92109 69167 92167 69173
rect 92477 69173 92489 69176
rect 92523 69173 92535 69207
rect 92477 69167 92535 69173
rect 92750 69164 92756 69216
rect 92808 69164 92814 69216
rect 98914 69164 98920 69216
rect 98972 69204 98978 69216
rect 99285 69207 99343 69213
rect 99285 69204 99297 69207
rect 98972 69176 99297 69204
rect 98972 69164 98978 69176
rect 99285 69173 99297 69176
rect 99331 69173 99343 69207
rect 99285 69167 99343 69173
rect 99650 69164 99656 69216
rect 99708 69204 99714 69216
rect 99745 69207 99803 69213
rect 99745 69204 99757 69207
rect 99708 69176 99757 69204
rect 99708 69164 99714 69176
rect 99745 69173 99757 69176
rect 99791 69173 99803 69207
rect 99745 69167 99803 69173
rect 100478 69164 100484 69216
rect 100536 69204 100542 69216
rect 101122 69204 101128 69216
rect 100536 69176 101128 69204
rect 100536 69164 100542 69176
rect 101122 69164 101128 69176
rect 101180 69164 101186 69216
rect 101766 69164 101772 69216
rect 101824 69164 101830 69216
rect 103149 69207 103207 69213
rect 103149 69173 103161 69207
rect 103195 69204 103207 69207
rect 103422 69204 103428 69216
rect 103195 69176 103428 69204
rect 103195 69173 103207 69176
rect 103149 69167 103207 69173
rect 103422 69164 103428 69176
rect 103480 69164 103486 69216
rect 103606 69164 103612 69216
rect 103664 69164 103670 69216
rect 104526 69164 104532 69216
rect 104584 69204 104590 69216
rect 104621 69207 104679 69213
rect 104621 69204 104633 69207
rect 104584 69176 104633 69204
rect 104584 69164 104590 69176
rect 104621 69173 104633 69176
rect 104667 69173 104679 69207
rect 104621 69167 104679 69173
rect 1104 69114 108836 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 96374 69114
rect 96426 69062 96438 69114
rect 96490 69062 96502 69114
rect 96554 69062 96566 69114
rect 96618 69062 96630 69114
rect 96682 69062 108836 69114
rect 1104 69040 108836 69062
rect 43806 68960 43812 69012
rect 43864 69000 43870 69012
rect 44729 69003 44787 69009
rect 44729 69000 44741 69003
rect 43864 68972 44741 69000
rect 43864 68960 43870 68972
rect 44729 68969 44741 68972
rect 44775 69000 44787 69003
rect 44775 68972 46428 69000
rect 44775 68969 44787 68972
rect 44729 68963 44787 68969
rect 42702 68892 42708 68944
rect 42760 68932 42766 68944
rect 45005 68935 45063 68941
rect 45005 68932 45017 68935
rect 42760 68904 45017 68932
rect 42760 68892 42766 68904
rect 45005 68901 45017 68904
rect 45051 68901 45063 68935
rect 45005 68895 45063 68901
rect 46400 68873 46428 68972
rect 58618 68960 58624 69012
rect 58676 68960 58682 69012
rect 60277 69003 60335 69009
rect 60277 68969 60289 69003
rect 60323 69000 60335 69003
rect 67358 69000 67364 69012
rect 60323 68972 64874 69000
rect 60323 68969 60335 68972
rect 60277 68963 60335 68969
rect 46385 68867 46443 68873
rect 46385 68833 46397 68867
rect 46431 68833 46443 68867
rect 58636 68864 58664 68960
rect 58897 68867 58955 68873
rect 58897 68864 58909 68867
rect 58636 68836 58909 68864
rect 46385 68827 46443 68833
rect 58897 68833 58909 68836
rect 58943 68833 58955 68867
rect 58897 68827 58955 68833
rect 64846 68796 64874 68972
rect 65628 68972 67364 69000
rect 65628 68873 65656 68972
rect 67358 68960 67364 68972
rect 67416 68960 67422 69012
rect 87049 69003 87107 69009
rect 87049 69000 87061 69003
rect 86926 68972 87061 69000
rect 66993 68935 67051 68941
rect 66993 68901 67005 68935
rect 67039 68932 67051 68935
rect 70394 68932 70400 68944
rect 67039 68904 70400 68932
rect 67039 68901 67051 68904
rect 66993 68895 67051 68901
rect 70394 68892 70400 68904
rect 70452 68892 70458 68944
rect 65613 68867 65671 68873
rect 65613 68833 65625 68867
rect 65659 68833 65671 68867
rect 65613 68827 65671 68833
rect 86926 68808 86954 68972
rect 87049 68969 87061 68972
rect 87095 69000 87107 69003
rect 89714 69000 89720 69012
rect 87095 68972 89720 69000
rect 87095 68969 87107 68972
rect 87049 68963 87107 68969
rect 89714 68960 89720 68972
rect 89772 69000 89778 69012
rect 90085 69003 90143 69009
rect 90085 69000 90097 69003
rect 89772 68972 90097 69000
rect 89772 68960 89778 68972
rect 68554 68796 68560 68808
rect 64846 68768 68560 68796
rect 68554 68756 68560 68768
rect 68612 68756 68618 68808
rect 86681 68799 86739 68805
rect 86681 68765 86693 68799
rect 86727 68796 86739 68799
rect 86862 68796 86868 68808
rect 86727 68768 86868 68796
rect 86727 68765 86739 68768
rect 86681 68759 86739 68765
rect 86862 68756 86868 68768
rect 86920 68768 86954 68808
rect 89824 68805 89852 68972
rect 90085 68969 90097 68972
rect 90131 68969 90143 69003
rect 90085 68963 90143 68969
rect 93302 68960 93308 69012
rect 93360 69000 93366 69012
rect 93581 69003 93639 69009
rect 93581 69000 93593 69003
rect 93360 68972 93593 69000
rect 93360 68960 93366 68972
rect 93581 68969 93593 68972
rect 93627 69000 93639 69003
rect 95970 69000 95976 69012
rect 93627 68972 95976 69000
rect 93627 68969 93639 68972
rect 93581 68963 93639 68969
rect 91649 68867 91707 68873
rect 91649 68833 91661 68867
rect 91695 68864 91707 68867
rect 91738 68864 91744 68876
rect 91695 68836 91744 68864
rect 91695 68833 91707 68836
rect 91649 68827 91707 68833
rect 91738 68824 91744 68836
rect 91796 68824 91802 68876
rect 89809 68799 89867 68805
rect 86920 68756 86926 68768
rect 89809 68765 89821 68799
rect 89855 68765 89867 68799
rect 91373 68799 91431 68805
rect 91373 68796 91385 68799
rect 89809 68759 89867 68765
rect 91112 68768 91385 68796
rect 42521 68731 42579 68737
rect 42521 68697 42533 68731
rect 42567 68728 42579 68731
rect 43714 68728 43720 68740
rect 42567 68700 43720 68728
rect 42567 68697 42579 68700
rect 42521 68691 42579 68697
rect 43714 68688 43720 68700
rect 43772 68688 43778 68740
rect 46140 68731 46198 68737
rect 46140 68697 46152 68731
rect 46186 68728 46198 68731
rect 46186 68700 46520 68728
rect 46186 68697 46198 68700
rect 46140 68691 46198 68697
rect 46492 68672 46520 68700
rect 58710 68688 58716 68740
rect 58768 68728 58774 68740
rect 59142 68731 59200 68737
rect 59142 68728 59154 68731
rect 58768 68700 59154 68728
rect 58768 68688 58774 68700
rect 59142 68697 59154 68700
rect 59188 68697 59200 68731
rect 59142 68691 59200 68697
rect 65880 68731 65938 68737
rect 65880 68697 65892 68731
rect 65926 68728 65938 68731
rect 66070 68728 66076 68740
rect 65926 68700 66076 68728
rect 65926 68697 65938 68700
rect 65880 68691 65938 68697
rect 66070 68688 66076 68700
rect 66128 68728 66134 68740
rect 91112 68737 91140 68768
rect 91373 68765 91385 68768
rect 91419 68765 91431 68799
rect 91373 68759 91431 68765
rect 93397 68799 93455 68805
rect 93397 68765 93409 68799
rect 93443 68796 93455 68799
rect 93596 68796 93624 68963
rect 95970 68960 95976 68972
rect 96028 69000 96034 69012
rect 96028 68972 96614 69000
rect 96028 68960 96034 68972
rect 96586 68932 96614 68972
rect 98270 68960 98276 69012
rect 98328 68960 98334 69012
rect 100573 69003 100631 69009
rect 100573 68969 100585 69003
rect 100619 69000 100631 69003
rect 100846 69000 100852 69012
rect 100619 68972 100852 69000
rect 100619 68969 100631 68972
rect 100573 68963 100631 68969
rect 100846 68960 100852 68972
rect 100904 68960 100910 69012
rect 102962 68960 102968 69012
rect 103020 69000 103026 69012
rect 103241 69003 103299 69009
rect 103241 69000 103253 69003
rect 103020 68972 103253 69000
rect 103020 68960 103026 68972
rect 103241 68969 103253 68972
rect 103287 68969 103299 69003
rect 103241 68963 103299 68969
rect 104802 68960 104808 69012
rect 104860 69000 104866 69012
rect 104986 69000 104992 69012
rect 104860 68972 104992 69000
rect 104860 68960 104866 68972
rect 104986 68960 104992 68972
rect 105044 69000 105050 69012
rect 105081 69003 105139 69009
rect 105081 69000 105093 69003
rect 105044 68972 105093 69000
rect 105044 68960 105050 68972
rect 105081 68969 105093 68972
rect 105127 68969 105139 69003
rect 105081 68963 105139 68969
rect 105262 68960 105268 69012
rect 105320 68960 105326 69012
rect 100294 68932 100300 68944
rect 96586 68904 100300 68932
rect 100294 68892 100300 68904
rect 100352 68892 100358 68944
rect 100757 68935 100815 68941
rect 100757 68901 100769 68935
rect 100803 68901 100815 68935
rect 100757 68895 100815 68901
rect 94869 68867 94927 68873
rect 94869 68833 94881 68867
rect 94915 68864 94927 68867
rect 95234 68864 95240 68876
rect 94915 68836 95240 68864
rect 94915 68833 94927 68836
rect 94869 68827 94927 68833
rect 95234 68824 95240 68836
rect 95292 68824 95298 68876
rect 95510 68824 95516 68876
rect 95568 68824 95574 68876
rect 95973 68867 96031 68873
rect 95973 68833 95985 68867
rect 96019 68864 96031 68867
rect 96154 68864 96160 68876
rect 96019 68836 96160 68864
rect 96019 68833 96031 68836
rect 95973 68827 96031 68833
rect 96154 68824 96160 68836
rect 96212 68864 96218 68876
rect 99929 68867 99987 68873
rect 99929 68864 99941 68867
rect 96212 68836 97120 68864
rect 96212 68824 96218 68836
rect 94777 68799 94835 68805
rect 94777 68796 94789 68799
rect 93443 68768 93624 68796
rect 94516 68768 94789 68796
rect 93443 68765 93455 68768
rect 93397 68759 93455 68765
rect 67085 68731 67143 68737
rect 67085 68728 67097 68731
rect 66128 68700 67097 68728
rect 66128 68688 66134 68700
rect 67085 68697 67097 68700
rect 67131 68697 67143 68731
rect 91097 68731 91155 68737
rect 91097 68728 91109 68731
rect 67085 68691 67143 68697
rect 89686 68700 91109 68728
rect 46474 68620 46480 68672
rect 46532 68620 46538 68672
rect 61470 68620 61476 68672
rect 61528 68620 61534 68672
rect 86770 68620 86776 68672
rect 86828 68620 86834 68672
rect 89254 68620 89260 68672
rect 89312 68660 89318 68672
rect 89686 68660 89714 68700
rect 91097 68697 91109 68700
rect 91143 68697 91155 68731
rect 91097 68691 91155 68697
rect 91204 68700 92138 68728
rect 89312 68632 89714 68660
rect 89901 68663 89959 68669
rect 89312 68620 89318 68632
rect 89901 68629 89913 68663
rect 89947 68660 89959 68663
rect 91204 68660 91232 68700
rect 94516 68672 94544 68768
rect 94777 68765 94789 68768
rect 94823 68796 94835 68799
rect 94958 68796 94964 68808
rect 94823 68768 94964 68796
rect 94823 68765 94835 68768
rect 94777 68759 94835 68765
rect 94958 68756 94964 68768
rect 95016 68756 95022 68808
rect 95881 68799 95939 68805
rect 95881 68765 95893 68799
rect 95927 68796 95939 68799
rect 96062 68796 96068 68808
rect 95927 68768 96068 68796
rect 95927 68765 95939 68768
rect 95881 68759 95939 68765
rect 96062 68756 96068 68768
rect 96120 68756 96126 68808
rect 97092 68805 97120 68836
rect 99346 68836 99941 68864
rect 97077 68799 97135 68805
rect 97077 68765 97089 68799
rect 97123 68765 97135 68799
rect 97077 68759 97135 68765
rect 97442 68756 97448 68808
rect 97500 68796 97506 68808
rect 98365 68799 98423 68805
rect 98365 68796 98377 68799
rect 97500 68768 98377 68796
rect 97500 68756 97506 68768
rect 98365 68765 98377 68768
rect 98411 68796 98423 68799
rect 99346 68796 99374 68836
rect 99929 68833 99941 68836
rect 99975 68864 99987 68867
rect 100772 68864 100800 68895
rect 101398 68864 101404 68876
rect 99975 68836 100708 68864
rect 100772 68836 101404 68864
rect 99975 68833 99987 68836
rect 99929 68827 99987 68833
rect 98411 68768 99374 68796
rect 99558 68799 99616 68805
rect 98411 68765 98423 68768
rect 98365 68759 98423 68765
rect 99558 68765 99570 68799
rect 99604 68796 99616 68799
rect 99742 68796 99748 68808
rect 99604 68768 99748 68796
rect 99604 68765 99616 68768
rect 99558 68759 99616 68765
rect 99742 68756 99748 68768
rect 99800 68756 99806 68808
rect 100021 68799 100079 68805
rect 100021 68765 100033 68799
rect 100067 68796 100079 68799
rect 100294 68796 100300 68808
rect 100067 68768 100300 68796
rect 100067 68765 100079 68768
rect 100021 68759 100079 68765
rect 100294 68756 100300 68768
rect 100352 68756 100358 68808
rect 100680 68796 100708 68836
rect 101398 68824 101404 68836
rect 101456 68824 101462 68876
rect 101766 68824 101772 68876
rect 101824 68864 101830 68876
rect 102137 68867 102195 68873
rect 102137 68864 102149 68867
rect 101824 68836 102149 68864
rect 101824 68824 101830 68836
rect 102137 68833 102149 68836
rect 102183 68833 102195 68867
rect 102137 68827 102195 68833
rect 102226 68824 102232 68876
rect 102284 68824 102290 68876
rect 102965 68867 103023 68873
rect 102965 68833 102977 68867
rect 103011 68864 103023 68867
rect 103146 68864 103152 68876
rect 103011 68836 103152 68864
rect 103011 68833 103023 68836
rect 102965 68827 103023 68833
rect 103146 68824 103152 68836
rect 103204 68824 103210 68876
rect 105354 68864 105360 68876
rect 103532 68836 105360 68864
rect 100849 68799 100907 68805
rect 100849 68796 100861 68799
rect 100680 68768 100861 68796
rect 100849 68765 100861 68768
rect 100895 68765 100907 68799
rect 100849 68759 100907 68765
rect 101033 68799 101091 68805
rect 101033 68765 101045 68799
rect 101079 68796 101091 68799
rect 101122 68796 101128 68808
rect 101079 68768 101128 68796
rect 101079 68765 101091 68768
rect 101033 68759 101091 68765
rect 101122 68756 101128 68768
rect 101180 68756 101186 68808
rect 101214 68756 101220 68808
rect 101272 68756 101278 68808
rect 103054 68756 103060 68808
rect 103112 68756 103118 68808
rect 103238 68756 103244 68808
rect 103296 68796 103302 68808
rect 103333 68799 103391 68805
rect 103333 68796 103345 68799
rect 103296 68768 103345 68796
rect 103296 68756 103302 68768
rect 103333 68765 103345 68768
rect 103379 68765 103391 68799
rect 103333 68759 103391 68765
rect 103422 68756 103428 68808
rect 103480 68756 103486 68808
rect 96080 68728 96108 68756
rect 97169 68731 97227 68737
rect 97169 68728 97181 68731
rect 96080 68700 97181 68728
rect 97169 68697 97181 68700
rect 97215 68697 97227 68731
rect 97169 68691 97227 68697
rect 97261 68731 97319 68737
rect 97261 68697 97273 68731
rect 97307 68728 97319 68731
rect 97994 68728 98000 68740
rect 97307 68700 98000 68728
rect 97307 68697 97319 68700
rect 97261 68691 97319 68697
rect 97994 68688 98000 68700
rect 98052 68728 98058 68740
rect 98730 68728 98736 68740
rect 98052 68700 98736 68728
rect 98052 68688 98058 68700
rect 98730 68688 98736 68700
rect 98788 68728 98794 68740
rect 99190 68728 99196 68740
rect 98788 68700 99196 68728
rect 98788 68688 98794 68700
rect 99190 68688 99196 68700
rect 99248 68688 99254 68740
rect 100389 68731 100447 68737
rect 100389 68697 100401 68731
rect 100435 68697 100447 68731
rect 100389 68691 100447 68697
rect 100605 68731 100663 68737
rect 100605 68697 100617 68731
rect 100651 68728 100663 68731
rect 100938 68728 100944 68740
rect 100651 68700 100944 68728
rect 100651 68697 100663 68700
rect 100605 68691 100663 68697
rect 89947 68632 91232 68660
rect 89947 68629 89959 68632
rect 89901 68623 89959 68629
rect 94498 68620 94504 68672
rect 94556 68620 94562 68672
rect 95142 68620 95148 68672
rect 95200 68620 95206 68672
rect 96890 68620 96896 68672
rect 96948 68620 96954 68672
rect 97902 68620 97908 68672
rect 97960 68660 97966 68672
rect 99377 68663 99435 68669
rect 99377 68660 99389 68663
rect 97960 68632 99389 68660
rect 97960 68620 97966 68632
rect 99377 68629 99389 68632
rect 99423 68629 99435 68663
rect 99377 68623 99435 68629
rect 99561 68663 99619 68669
rect 99561 68629 99573 68663
rect 99607 68660 99619 68663
rect 99650 68660 99656 68672
rect 99607 68632 99656 68660
rect 99607 68629 99619 68632
rect 99561 68623 99619 68629
rect 99650 68620 99656 68632
rect 99708 68620 99714 68672
rect 100404 68660 100432 68691
rect 100938 68688 100944 68700
rect 100996 68688 101002 68740
rect 101232 68728 101260 68756
rect 103532 68728 103560 68836
rect 103606 68756 103612 68808
rect 103664 68756 103670 68808
rect 103698 68756 103704 68808
rect 103756 68796 103762 68808
rect 104529 68799 104587 68805
rect 103756 68768 104388 68796
rect 103756 68756 103762 68768
rect 101140 68700 103560 68728
rect 101140 68672 101168 68700
rect 101122 68660 101128 68672
rect 100404 68632 101128 68660
rect 101122 68620 101128 68632
rect 101180 68620 101186 68672
rect 101214 68620 101220 68672
rect 101272 68660 101278 68672
rect 101677 68663 101735 68669
rect 101677 68660 101689 68663
rect 101272 68632 101689 68660
rect 101272 68620 101278 68632
rect 101677 68629 101689 68632
rect 101723 68629 101735 68663
rect 101677 68623 101735 68629
rect 102042 68620 102048 68672
rect 102100 68620 102106 68672
rect 102597 68663 102655 68669
rect 102597 68629 102609 68663
rect 102643 68660 102655 68663
rect 102870 68660 102876 68672
rect 102643 68632 102876 68660
rect 102643 68629 102655 68632
rect 102597 68623 102655 68629
rect 102870 68620 102876 68632
rect 102928 68660 102934 68672
rect 104360 68669 104388 68768
rect 104529 68765 104541 68799
rect 104575 68796 104587 68799
rect 104618 68796 104624 68808
rect 104575 68768 104624 68796
rect 104575 68765 104587 68768
rect 104529 68759 104587 68765
rect 104618 68756 104624 68768
rect 104676 68756 104682 68808
rect 104802 68756 104808 68808
rect 104860 68756 104866 68808
rect 105004 68805 105032 68836
rect 105354 68824 105360 68836
rect 105412 68824 105418 68876
rect 104989 68799 105047 68805
rect 104989 68765 105001 68799
rect 105035 68765 105047 68799
rect 104989 68759 105047 68765
rect 104894 68688 104900 68740
rect 104952 68728 104958 68740
rect 105170 68728 105176 68740
rect 104952 68700 105176 68728
rect 104952 68688 104958 68700
rect 105170 68688 105176 68700
rect 105228 68737 105234 68740
rect 105228 68731 105291 68737
rect 105228 68697 105245 68731
rect 105279 68697 105291 68731
rect 105228 68691 105291 68697
rect 105228 68688 105234 68691
rect 105446 68688 105452 68740
rect 105504 68688 105510 68740
rect 103885 68663 103943 68669
rect 103885 68660 103897 68663
rect 102928 68632 103897 68660
rect 102928 68620 102934 68632
rect 103885 68629 103897 68632
rect 103931 68629 103943 68663
rect 103885 68623 103943 68629
rect 104345 68663 104403 68669
rect 104345 68629 104357 68663
rect 104391 68660 104403 68663
rect 104434 68660 104440 68672
rect 104391 68632 104440 68660
rect 104391 68629 104403 68632
rect 104345 68623 104403 68629
rect 104434 68620 104440 68632
rect 104492 68620 104498 68672
rect 1104 68570 108836 68592
rect 1104 68518 4874 68570
rect 4926 68518 4938 68570
rect 4990 68518 5002 68570
rect 5054 68518 5066 68570
rect 5118 68518 5130 68570
rect 5182 68518 35594 68570
rect 35646 68518 35658 68570
rect 35710 68518 35722 68570
rect 35774 68518 35786 68570
rect 35838 68518 35850 68570
rect 35902 68518 66314 68570
rect 66366 68518 66378 68570
rect 66430 68518 66442 68570
rect 66494 68518 66506 68570
rect 66558 68518 66570 68570
rect 66622 68518 97034 68570
rect 97086 68518 97098 68570
rect 97150 68518 97162 68570
rect 97214 68518 97226 68570
rect 97278 68518 97290 68570
rect 97342 68518 108836 68570
rect 1104 68496 108836 68518
rect 38654 68416 38660 68468
rect 38712 68416 38718 68468
rect 38838 68416 38844 68468
rect 38896 68416 38902 68468
rect 91554 68416 91560 68468
rect 91612 68416 91618 68468
rect 91725 68459 91783 68465
rect 91725 68425 91737 68459
rect 91771 68456 91783 68459
rect 92934 68456 92940 68468
rect 91771 68428 92940 68456
rect 91771 68425 91783 68428
rect 91725 68419 91783 68425
rect 92934 68416 92940 68428
rect 92992 68416 92998 68468
rect 96062 68416 96068 68468
rect 96120 68456 96126 68468
rect 96249 68459 96307 68465
rect 96249 68456 96261 68459
rect 96120 68428 96261 68456
rect 96120 68416 96126 68428
rect 96249 68425 96261 68428
rect 96295 68425 96307 68459
rect 96249 68419 96307 68425
rect 96341 68459 96399 68465
rect 96341 68425 96353 68459
rect 96387 68425 96399 68459
rect 96341 68419 96399 68425
rect 38672 68388 38700 68416
rect 42150 68388 42156 68400
rect 38672 68360 42156 68388
rect 39942 68280 39948 68332
rect 40000 68329 40006 68332
rect 40236 68329 40264 68360
rect 42150 68348 42156 68360
rect 42208 68348 42214 68400
rect 91002 68348 91008 68400
rect 91060 68388 91066 68400
rect 91922 68388 91928 68400
rect 91060 68360 91928 68388
rect 91060 68348 91066 68360
rect 91922 68348 91928 68360
rect 91980 68388 91986 68400
rect 92290 68388 92296 68400
rect 91980 68360 92296 68388
rect 91980 68348 91986 68360
rect 92290 68348 92296 68360
rect 92348 68348 92354 68400
rect 94774 68348 94780 68400
rect 94832 68388 94838 68400
rect 94961 68391 95019 68397
rect 94961 68388 94973 68391
rect 94832 68360 94973 68388
rect 94832 68348 94838 68360
rect 94961 68357 94973 68360
rect 95007 68357 95019 68391
rect 96080 68388 96108 68416
rect 94961 68351 95019 68357
rect 95804 68360 96108 68388
rect 96356 68388 96384 68419
rect 98178 68416 98184 68468
rect 98236 68416 98242 68468
rect 100110 68416 100116 68468
rect 100168 68456 100174 68468
rect 100205 68459 100263 68465
rect 100205 68456 100217 68459
rect 100168 68428 100217 68456
rect 100168 68416 100174 68428
rect 100205 68425 100217 68428
rect 100251 68425 100263 68459
rect 100205 68419 100263 68425
rect 100294 68416 100300 68468
rect 100352 68456 100358 68468
rect 101769 68459 101827 68465
rect 101769 68456 101781 68459
rect 100352 68428 100708 68456
rect 100352 68416 100358 68428
rect 97994 68388 98000 68400
rect 96356 68360 98000 68388
rect 40000 68283 40012 68329
rect 40221 68323 40279 68329
rect 40221 68289 40233 68323
rect 40267 68289 40279 68323
rect 40221 68283 40279 68289
rect 40000 68280 40006 68283
rect 95234 68280 95240 68332
rect 95292 68280 95298 68332
rect 95804 68329 95832 68360
rect 95789 68323 95847 68329
rect 95789 68289 95801 68323
rect 95835 68289 95847 68323
rect 95789 68283 95847 68289
rect 95973 68323 96031 68329
rect 95973 68289 95985 68323
rect 96019 68320 96031 68323
rect 96154 68320 96160 68332
rect 96019 68292 96160 68320
rect 96019 68289 96031 68292
rect 95973 68283 96031 68289
rect 96154 68280 96160 68292
rect 96212 68280 96218 68332
rect 96246 68280 96252 68332
rect 96304 68320 96310 68332
rect 96356 68320 96384 68360
rect 96304 68292 96384 68320
rect 96525 68323 96583 68329
rect 96304 68280 96310 68292
rect 96525 68289 96537 68323
rect 96571 68320 96583 68323
rect 97077 68323 97135 68329
rect 97077 68320 97089 68323
rect 96571 68292 97089 68320
rect 96571 68289 96583 68292
rect 96525 68283 96583 68289
rect 97077 68289 97089 68292
rect 97123 68320 97135 68323
rect 97442 68320 97448 68332
rect 97123 68292 97448 68320
rect 97123 68289 97135 68292
rect 97077 68283 97135 68289
rect 97442 68280 97448 68292
rect 97500 68280 97506 68332
rect 95050 68212 95056 68264
rect 95108 68212 95114 68264
rect 96172 68252 96200 68280
rect 97552 68261 97580 68360
rect 97994 68348 98000 68360
rect 98052 68348 98058 68400
rect 99926 68348 99932 68400
rect 99984 68388 99990 68400
rect 100573 68391 100631 68397
rect 100573 68388 100585 68391
rect 99984 68360 100585 68388
rect 99984 68348 99990 68360
rect 100573 68357 100585 68360
rect 100619 68357 100631 68391
rect 100680 68388 100708 68428
rect 100956 68428 101781 68456
rect 100956 68388 100984 68428
rect 101769 68425 101781 68428
rect 101815 68425 101827 68459
rect 101769 68419 101827 68425
rect 101858 68416 101864 68468
rect 101916 68456 101922 68468
rect 101953 68459 102011 68465
rect 101953 68456 101965 68459
rect 101916 68428 101965 68456
rect 101916 68416 101922 68428
rect 101953 68425 101965 68428
rect 101999 68456 102011 68459
rect 102318 68456 102324 68468
rect 101999 68428 102324 68456
rect 101999 68425 102011 68428
rect 101953 68419 102011 68425
rect 102318 68416 102324 68428
rect 102376 68416 102382 68468
rect 102410 68416 102416 68468
rect 102468 68456 102474 68468
rect 102965 68459 103023 68465
rect 102965 68456 102977 68459
rect 102468 68428 102977 68456
rect 102468 68416 102474 68428
rect 102965 68425 102977 68428
rect 103011 68425 103023 68459
rect 102965 68419 103023 68425
rect 103333 68459 103391 68465
rect 103333 68425 103345 68459
rect 103379 68456 103391 68459
rect 103606 68456 103612 68468
rect 103379 68428 103612 68456
rect 103379 68425 103391 68428
rect 103333 68419 103391 68425
rect 103606 68416 103612 68428
rect 103664 68416 103670 68468
rect 105081 68459 105139 68465
rect 105081 68456 105093 68459
rect 103900 68428 105093 68456
rect 101214 68388 101220 68400
rect 100680 68360 100984 68388
rect 101048 68360 101220 68388
rect 100573 68351 100631 68357
rect 97626 68280 97632 68332
rect 97684 68320 97690 68332
rect 97813 68323 97871 68329
rect 97813 68320 97825 68323
rect 97684 68292 97825 68320
rect 97684 68280 97690 68292
rect 97813 68289 97825 68292
rect 97859 68289 97871 68323
rect 97813 68283 97871 68289
rect 98546 68280 98552 68332
rect 98604 68320 98610 68332
rect 99101 68323 99159 68329
rect 99101 68320 99113 68323
rect 98604 68292 99113 68320
rect 98604 68280 98610 68292
rect 99101 68289 99113 68292
rect 99147 68289 99159 68323
rect 99101 68283 99159 68289
rect 99282 68280 99288 68332
rect 99340 68280 99346 68332
rect 99558 68280 99564 68332
rect 99616 68280 99622 68332
rect 99834 68280 99840 68332
rect 99892 68280 99898 68332
rect 100202 68280 100208 68332
rect 100260 68320 100266 68332
rect 100389 68323 100447 68329
rect 100389 68320 100401 68323
rect 100260 68292 100401 68320
rect 100260 68280 100266 68292
rect 100389 68289 100401 68292
rect 100435 68289 100447 68323
rect 100389 68283 100447 68289
rect 96801 68255 96859 68261
rect 96801 68252 96813 68255
rect 96172 68224 96813 68252
rect 96801 68221 96813 68224
rect 96847 68221 96859 68255
rect 96801 68215 96859 68221
rect 96893 68255 96951 68261
rect 96893 68221 96905 68255
rect 96939 68221 96951 68255
rect 96893 68215 96951 68221
rect 96985 68255 97043 68261
rect 96985 68221 96997 68255
rect 97031 68252 97043 68255
rect 97537 68255 97595 68261
rect 97537 68252 97549 68255
rect 97031 68224 97549 68252
rect 97031 68221 97043 68224
rect 96985 68215 97043 68221
rect 97537 68221 97549 68224
rect 97583 68221 97595 68255
rect 97537 68215 97595 68221
rect 97721 68255 97779 68261
rect 97721 68221 97733 68255
rect 97767 68252 97779 68255
rect 97902 68252 97908 68264
rect 97767 68224 97908 68252
rect 97767 68221 97779 68224
rect 97721 68215 97779 68221
rect 95786 68144 95792 68196
rect 95844 68184 95850 68196
rect 96249 68187 96307 68193
rect 96249 68184 96261 68187
rect 95844 68156 96261 68184
rect 95844 68144 95850 68156
rect 96249 68153 96261 68156
rect 96295 68153 96307 68187
rect 96908 68184 96936 68215
rect 97902 68212 97908 68224
rect 97960 68212 97966 68264
rect 99466 68212 99472 68264
rect 99524 68252 99530 68264
rect 99929 68255 99987 68261
rect 99929 68252 99941 68255
rect 99524 68224 99941 68252
rect 99524 68212 99530 68224
rect 99929 68221 99941 68224
rect 99975 68221 99987 68255
rect 99929 68215 99987 68221
rect 100113 68255 100171 68261
rect 100113 68221 100125 68255
rect 100159 68252 100171 68255
rect 100404 68252 100432 68283
rect 100662 68280 100668 68332
rect 100720 68280 100726 68332
rect 100757 68323 100815 68329
rect 100757 68289 100769 68323
rect 100803 68320 100815 68323
rect 100846 68320 100852 68332
rect 100803 68292 100852 68320
rect 100803 68289 100815 68292
rect 100757 68283 100815 68289
rect 100846 68280 100852 68292
rect 100904 68280 100910 68332
rect 101048 68320 101076 68360
rect 101214 68348 101220 68360
rect 101272 68348 101278 68400
rect 101398 68348 101404 68400
rect 101456 68348 101462 68400
rect 100956 68292 101076 68320
rect 100956 68252 100984 68292
rect 101122 68280 101128 68332
rect 101180 68280 101186 68332
rect 101585 68323 101643 68329
rect 101585 68289 101597 68323
rect 101631 68320 101643 68323
rect 101861 68323 101919 68329
rect 101861 68320 101873 68323
rect 101631 68292 101873 68320
rect 101631 68289 101643 68292
rect 101585 68283 101643 68289
rect 101861 68289 101873 68292
rect 101907 68289 101919 68323
rect 101861 68283 101919 68289
rect 102137 68323 102195 68329
rect 102137 68289 102149 68323
rect 102183 68320 102195 68323
rect 102226 68320 102232 68332
rect 102183 68292 102232 68320
rect 102183 68289 102195 68292
rect 102137 68283 102195 68289
rect 100159 68224 100248 68252
rect 100404 68224 100984 68252
rect 100159 68221 100171 68224
rect 100113 68215 100171 68221
rect 96249 68147 96307 68153
rect 96540 68156 96936 68184
rect 91741 68119 91799 68125
rect 91741 68085 91753 68119
rect 91787 68116 91799 68119
rect 93394 68116 93400 68128
rect 91787 68088 93400 68116
rect 91787 68085 91799 68088
rect 91741 68079 91799 68085
rect 93394 68076 93400 68088
rect 93452 68076 93458 68128
rect 95142 68076 95148 68128
rect 95200 68076 95206 68128
rect 95326 68076 95332 68128
rect 95384 68116 95390 68128
rect 95421 68119 95479 68125
rect 95421 68116 95433 68119
rect 95384 68088 95433 68116
rect 95384 68076 95390 68088
rect 95421 68085 95433 68088
rect 95467 68085 95479 68119
rect 95421 68079 95479 68085
rect 95878 68076 95884 68128
rect 95936 68076 95942 68128
rect 96062 68076 96068 68128
rect 96120 68116 96126 68128
rect 96540 68116 96568 68156
rect 96120 68088 96568 68116
rect 96617 68119 96675 68125
rect 96120 68076 96126 68088
rect 96617 68085 96629 68119
rect 96663 68116 96675 68119
rect 96706 68116 96712 68128
rect 96663 68088 96712 68116
rect 96663 68085 96675 68088
rect 96617 68079 96675 68085
rect 96706 68076 96712 68088
rect 96764 68076 96770 68128
rect 100220 68116 100248 68224
rect 101030 68212 101036 68264
rect 101088 68252 101094 68264
rect 101309 68255 101367 68261
rect 101309 68252 101321 68255
rect 101088 68224 101321 68252
rect 101088 68212 101094 68224
rect 101309 68221 101321 68224
rect 101355 68221 101367 68255
rect 101309 68215 101367 68221
rect 100294 68144 100300 68196
rect 100352 68184 100358 68196
rect 100849 68187 100907 68193
rect 100849 68184 100861 68187
rect 100352 68156 100861 68184
rect 100352 68144 100358 68156
rect 100849 68153 100861 68156
rect 100895 68184 100907 68187
rect 101600 68184 101628 68283
rect 102226 68280 102232 68292
rect 102284 68280 102290 68332
rect 103149 68323 103207 68329
rect 103149 68289 103161 68323
rect 103195 68320 103207 68323
rect 103330 68320 103336 68332
rect 103195 68292 103336 68320
rect 103195 68289 103207 68292
rect 103149 68283 103207 68289
rect 103330 68280 103336 68292
rect 103388 68280 103394 68332
rect 103425 68323 103483 68329
rect 103425 68289 103437 68323
rect 103471 68320 103483 68323
rect 103698 68320 103704 68332
rect 103471 68292 103704 68320
rect 103471 68289 103483 68292
rect 103425 68283 103483 68289
rect 103698 68280 103704 68292
rect 103756 68280 103762 68332
rect 103900 68329 103928 68428
rect 105081 68425 105093 68428
rect 105127 68456 105139 68459
rect 105262 68456 105268 68468
rect 105127 68428 105268 68456
rect 105127 68425 105139 68428
rect 105081 68419 105139 68425
rect 105262 68416 105268 68428
rect 105320 68416 105326 68468
rect 104084 68360 105216 68388
rect 104084 68329 104112 68360
rect 105188 68332 105216 68360
rect 103885 68323 103943 68329
rect 103885 68289 103897 68323
rect 103931 68289 103943 68323
rect 103885 68283 103943 68289
rect 104069 68323 104127 68329
rect 104069 68289 104081 68323
rect 104115 68289 104127 68323
rect 104621 68323 104679 68329
rect 104621 68320 104633 68323
rect 104069 68283 104127 68289
rect 104176 68292 104633 68320
rect 104176 68252 104204 68292
rect 104621 68289 104633 68292
rect 104667 68289 104679 68323
rect 104621 68283 104679 68289
rect 104894 68280 104900 68332
rect 104952 68280 104958 68332
rect 105170 68280 105176 68332
rect 105228 68280 105234 68332
rect 100895 68156 101628 68184
rect 101692 68224 104204 68252
rect 100895 68153 100907 68156
rect 100849 68147 100907 68153
rect 100570 68116 100576 68128
rect 100220 68088 100576 68116
rect 100570 68076 100576 68088
rect 100628 68116 100634 68128
rect 101692 68116 101720 68224
rect 104526 68212 104532 68264
rect 104584 68212 104590 68264
rect 104912 68252 104940 68280
rect 105446 68252 105452 68264
rect 104912 68224 105452 68252
rect 105446 68212 105452 68224
rect 105504 68212 105510 68264
rect 101950 68144 101956 68196
rect 102008 68184 102014 68196
rect 102137 68187 102195 68193
rect 102137 68184 102149 68187
rect 102008 68156 102149 68184
rect 102008 68144 102014 68156
rect 102137 68153 102149 68156
rect 102183 68153 102195 68187
rect 102137 68147 102195 68153
rect 102502 68144 102508 68196
rect 102560 68184 102566 68196
rect 104253 68187 104311 68193
rect 104253 68184 104265 68187
rect 102560 68156 104265 68184
rect 102560 68144 102566 68156
rect 104253 68153 104265 68156
rect 104299 68153 104311 68187
rect 104253 68147 104311 68153
rect 104618 68144 104624 68196
rect 104676 68184 104682 68196
rect 104897 68187 104955 68193
rect 104897 68184 104909 68187
rect 104676 68156 104909 68184
rect 104676 68144 104682 68156
rect 104897 68153 104909 68156
rect 104943 68153 104955 68187
rect 104897 68147 104955 68153
rect 100628 68088 101720 68116
rect 100628 68076 100634 68088
rect 103974 68076 103980 68128
rect 104032 68076 104038 68128
rect 1104 68026 108836 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 96374 68026
rect 96426 67974 96438 68026
rect 96490 67974 96502 68026
rect 96554 67974 96566 68026
rect 96618 67974 96630 68026
rect 96682 67974 108836 68026
rect 1104 67952 108836 67974
rect 89070 67872 89076 67924
rect 89128 67912 89134 67924
rect 89257 67915 89315 67921
rect 89257 67912 89269 67915
rect 89128 67884 89269 67912
rect 89128 67872 89134 67884
rect 89257 67881 89269 67884
rect 89303 67912 89315 67915
rect 89438 67912 89444 67924
rect 89303 67884 89444 67912
rect 89303 67881 89315 67884
rect 89257 67875 89315 67881
rect 89438 67872 89444 67884
rect 89496 67872 89502 67924
rect 89717 67915 89775 67921
rect 89717 67881 89729 67915
rect 89763 67912 89775 67915
rect 90818 67912 90824 67924
rect 89763 67884 90824 67912
rect 89763 67881 89775 67884
rect 89717 67875 89775 67881
rect 90818 67872 90824 67884
rect 90876 67872 90882 67924
rect 91922 67872 91928 67924
rect 91980 67912 91986 67924
rect 94685 67915 94743 67921
rect 94685 67912 94697 67915
rect 91980 67884 94697 67912
rect 91980 67872 91986 67884
rect 94685 67881 94697 67884
rect 94731 67881 94743 67915
rect 94685 67875 94743 67881
rect 98730 67872 98736 67924
rect 98788 67912 98794 67924
rect 98917 67915 98975 67921
rect 98917 67912 98929 67915
rect 98788 67884 98929 67912
rect 98788 67872 98794 67884
rect 98917 67881 98929 67884
rect 98963 67912 98975 67915
rect 99282 67912 99288 67924
rect 98963 67884 99288 67912
rect 98963 67881 98975 67884
rect 98917 67875 98975 67881
rect 99282 67872 99288 67884
rect 99340 67872 99346 67924
rect 100018 67872 100024 67924
rect 100076 67912 100082 67924
rect 100297 67915 100355 67921
rect 100297 67912 100309 67915
rect 100076 67884 100309 67912
rect 100076 67872 100082 67884
rect 100297 67881 100309 67884
rect 100343 67881 100355 67915
rect 100297 67875 100355 67881
rect 101674 67872 101680 67924
rect 101732 67872 101738 67924
rect 101766 67872 101772 67924
rect 101824 67912 101830 67924
rect 102686 67912 102692 67924
rect 101824 67884 102692 67912
rect 101824 67872 101830 67884
rect 102686 67872 102692 67884
rect 102744 67872 102750 67924
rect 107930 67872 107936 67924
rect 107988 67912 107994 67924
rect 108301 67915 108359 67921
rect 108301 67912 108313 67915
rect 107988 67884 108313 67912
rect 107988 67872 107994 67884
rect 108301 67881 108313 67884
rect 108347 67881 108359 67915
rect 108301 67875 108359 67881
rect 89533 67847 89591 67853
rect 89533 67813 89545 67847
rect 89579 67813 89591 67847
rect 89533 67807 89591 67813
rect 86770 67736 86776 67788
rect 86828 67776 86834 67788
rect 88705 67779 88763 67785
rect 86828 67748 87644 67776
rect 86828 67736 86834 67748
rect 84749 67711 84807 67717
rect 84749 67677 84761 67711
rect 84795 67708 84807 67711
rect 84933 67711 84991 67717
rect 84933 67708 84945 67711
rect 84795 67680 84945 67708
rect 84795 67677 84807 67680
rect 84749 67671 84807 67677
rect 84933 67677 84945 67680
rect 84979 67708 84991 67711
rect 86034 67708 86040 67720
rect 84979 67680 86040 67708
rect 84979 67677 84991 67680
rect 84933 67671 84991 67677
rect 86034 67668 86040 67680
rect 86092 67708 86098 67720
rect 86865 67711 86923 67717
rect 86865 67708 86877 67711
rect 86092 67680 86877 67708
rect 86092 67668 86098 67680
rect 86865 67677 86877 67680
rect 86911 67708 86923 67711
rect 87138 67708 87144 67720
rect 86911 67680 87144 67708
rect 86911 67677 86923 67680
rect 86865 67671 86923 67677
rect 87138 67668 87144 67680
rect 87196 67668 87202 67720
rect 87616 67694 87644 67748
rect 88705 67745 88717 67779
rect 88751 67776 88763 67779
rect 89548 67776 89576 67807
rect 94406 67804 94412 67856
rect 94464 67844 94470 67856
rect 95053 67847 95111 67853
rect 95053 67844 95065 67847
rect 94464 67816 95065 67844
rect 94464 67804 94470 67816
rect 95053 67813 95065 67816
rect 95099 67813 95111 67847
rect 98822 67844 98828 67856
rect 95053 67807 95111 67813
rect 97828 67816 98828 67844
rect 88751 67748 89576 67776
rect 88751 67745 88763 67748
rect 88705 67739 88763 67745
rect 94958 67736 94964 67788
rect 95016 67736 95022 67788
rect 95182 67779 95240 67785
rect 95182 67745 95194 67779
rect 95228 67776 95240 67779
rect 95694 67776 95700 67788
rect 95228 67748 95700 67776
rect 95228 67745 95240 67748
rect 95182 67739 95240 67745
rect 95694 67736 95700 67748
rect 95752 67736 95758 67788
rect 95878 67736 95884 67788
rect 95936 67736 95942 67788
rect 88981 67711 89039 67717
rect 88981 67677 88993 67711
rect 89027 67708 89039 67711
rect 89254 67708 89260 67720
rect 89027 67680 89260 67708
rect 89027 67677 89039 67680
rect 88981 67671 89039 67677
rect 89254 67668 89260 67680
rect 89312 67668 89318 67720
rect 89456 67680 89944 67708
rect 70210 67600 70216 67652
rect 70268 67640 70274 67652
rect 74350 67640 74356 67652
rect 70268 67612 74356 67640
rect 70268 67600 70274 67612
rect 74350 67600 74356 67612
rect 74408 67640 74414 67652
rect 89456 67649 89484 67680
rect 89714 67649 89720 67652
rect 82817 67643 82875 67649
rect 82817 67640 82829 67643
rect 74408 67612 82829 67640
rect 74408 67600 74414 67612
rect 82817 67609 82829 67612
rect 82863 67640 82875 67643
rect 83001 67643 83059 67649
rect 83001 67640 83013 67643
rect 82863 67612 83013 67640
rect 82863 67609 82875 67612
rect 82817 67603 82875 67609
rect 83001 67609 83013 67612
rect 83047 67609 83059 67643
rect 83001 67603 83059 67609
rect 86957 67643 87015 67649
rect 86957 67609 86969 67643
rect 87003 67640 87015 67643
rect 89441 67643 89499 67649
rect 87003 67612 87460 67640
rect 87003 67609 87015 67612
rect 86957 67603 87015 67609
rect 87432 67584 87460 67612
rect 89441 67609 89453 67643
rect 89487 67609 89499 67643
rect 89441 67603 89499 67609
rect 89701 67643 89720 67649
rect 89701 67609 89713 67643
rect 89701 67603 89720 67609
rect 89714 67600 89720 67603
rect 89772 67600 89778 67652
rect 89916 67649 89944 67680
rect 95326 67668 95332 67720
rect 95384 67668 95390 67720
rect 95789 67711 95847 67717
rect 95789 67677 95801 67711
rect 95835 67708 95847 67711
rect 96246 67708 96252 67720
rect 95835 67680 96252 67708
rect 95835 67677 95847 67680
rect 95789 67671 95847 67677
rect 96246 67668 96252 67680
rect 96304 67668 96310 67720
rect 97828 67708 97856 67816
rect 98822 67804 98828 67816
rect 98880 67844 98886 67856
rect 98880 67816 99052 67844
rect 98880 67804 98886 67816
rect 97902 67736 97908 67788
rect 97960 67776 97966 67788
rect 97960 67748 98224 67776
rect 97960 67736 97966 67748
rect 98196 67717 98224 67748
rect 98546 67736 98552 67788
rect 98604 67736 98610 67788
rect 98656 67748 98868 67776
rect 97997 67711 98055 67717
rect 97997 67708 98009 67711
rect 97828 67680 98009 67708
rect 97997 67677 98009 67680
rect 98043 67677 98055 67711
rect 97997 67671 98055 67677
rect 98181 67711 98239 67717
rect 98181 67677 98193 67711
rect 98227 67708 98239 67711
rect 98656 67708 98684 67748
rect 98840 67717 98868 67748
rect 99024 67717 99052 67816
rect 99190 67804 99196 67856
rect 99248 67844 99254 67856
rect 99248 67816 99374 67844
rect 99248 67804 99254 67816
rect 99346 67776 99374 67816
rect 99742 67804 99748 67856
rect 99800 67844 99806 67856
rect 100754 67844 100760 67856
rect 99800 67816 100760 67844
rect 99800 67804 99806 67816
rect 100754 67804 100760 67816
rect 100812 67804 100818 67856
rect 102870 67844 102876 67856
rect 101324 67816 102876 67844
rect 99466 67776 99472 67788
rect 99346 67748 99472 67776
rect 99466 67736 99472 67748
rect 99524 67776 99530 67788
rect 101324 67785 101352 67816
rect 102870 67804 102876 67816
rect 102928 67804 102934 67856
rect 102962 67804 102968 67856
rect 103020 67804 103026 67856
rect 99653 67779 99711 67785
rect 99653 67776 99665 67779
rect 99524 67748 99665 67776
rect 99524 67736 99530 67748
rect 99653 67745 99665 67748
rect 99699 67745 99711 67779
rect 99653 67739 99711 67745
rect 101309 67779 101367 67785
rect 101309 67745 101321 67779
rect 101355 67745 101367 67779
rect 101309 67739 101367 67745
rect 102318 67736 102324 67788
rect 102376 67736 102382 67788
rect 98227 67680 98684 67708
rect 98733 67711 98791 67717
rect 98227 67677 98239 67680
rect 98181 67671 98239 67677
rect 98733 67677 98745 67711
rect 98779 67677 98791 67711
rect 98733 67671 98791 67677
rect 98825 67711 98883 67717
rect 98825 67677 98837 67711
rect 98871 67677 98883 67711
rect 98825 67671 98883 67677
rect 99009 67711 99067 67717
rect 99009 67677 99021 67711
rect 99055 67677 99067 67711
rect 99009 67671 99067 67677
rect 89901 67643 89959 67649
rect 89901 67609 89913 67643
rect 89947 67640 89959 67643
rect 89990 67640 89996 67652
rect 89947 67612 89996 67640
rect 89947 67609 89959 67612
rect 89901 67603 89959 67609
rect 89990 67600 89996 67612
rect 90048 67640 90054 67652
rect 91002 67640 91008 67652
rect 90048 67612 91008 67640
rect 90048 67600 90054 67612
rect 91002 67600 91008 67612
rect 91060 67600 91066 67652
rect 98270 67600 98276 67652
rect 98328 67640 98334 67652
rect 98748 67640 98776 67671
rect 99098 67668 99104 67720
rect 99156 67708 99162 67720
rect 100941 67711 100999 67717
rect 100941 67708 100953 67711
rect 99156 67680 100953 67708
rect 99156 67668 99162 67680
rect 100941 67677 100953 67680
rect 100987 67708 100999 67711
rect 101030 67708 101036 67720
rect 100987 67680 101036 67708
rect 100987 67677 100999 67680
rect 100941 67671 100999 67677
rect 101030 67668 101036 67680
rect 101088 67668 101094 67720
rect 101125 67711 101183 67717
rect 101125 67677 101137 67711
rect 101171 67708 101183 67711
rect 101674 67708 101680 67720
rect 101171 67680 101680 67708
rect 101171 67677 101183 67680
rect 101125 67671 101183 67677
rect 101674 67668 101680 67680
rect 101732 67668 101738 67720
rect 101861 67711 101919 67717
rect 101861 67677 101873 67711
rect 101907 67677 101919 67711
rect 101861 67671 101919 67677
rect 98914 67640 98920 67652
rect 98328 67612 98920 67640
rect 98328 67600 98334 67612
rect 98914 67600 98920 67612
rect 98972 67600 98978 67652
rect 99742 67600 99748 67652
rect 99800 67640 99806 67652
rect 99929 67643 99987 67649
rect 99929 67640 99941 67643
rect 99800 67612 99941 67640
rect 99800 67600 99806 67612
rect 99929 67609 99941 67612
rect 99975 67609 99987 67643
rect 99929 67603 99987 67609
rect 100294 67600 100300 67652
rect 100352 67640 100358 67652
rect 101876 67640 101904 67671
rect 101950 67668 101956 67720
rect 102008 67668 102014 67720
rect 102134 67668 102140 67720
rect 102192 67668 102198 67720
rect 102226 67668 102232 67720
rect 102284 67702 102290 67720
rect 102284 67674 102323 67702
rect 102284 67668 102290 67674
rect 102502 67668 102508 67720
rect 102560 67668 102566 67720
rect 102597 67711 102655 67717
rect 102597 67677 102609 67711
rect 102643 67708 102655 67711
rect 102686 67708 102692 67720
rect 102643 67680 102692 67708
rect 102643 67677 102655 67680
rect 102597 67671 102655 67677
rect 102686 67668 102692 67680
rect 102744 67668 102750 67720
rect 102778 67668 102784 67720
rect 102836 67668 102842 67720
rect 102873 67711 102931 67717
rect 102873 67677 102885 67711
rect 102919 67708 102931 67711
rect 103241 67711 103299 67717
rect 102919 67680 103100 67708
rect 102919 67677 102931 67680
rect 102873 67671 102931 67677
rect 102229 67665 102287 67668
rect 100352 67612 101904 67640
rect 100352 67600 100358 67612
rect 102410 67600 102416 67652
rect 102468 67640 102474 67652
rect 102965 67643 103023 67649
rect 102965 67640 102977 67643
rect 102468 67612 102977 67640
rect 102468 67600 102474 67612
rect 102965 67609 102977 67612
rect 103011 67609 103023 67643
rect 102965 67603 103023 67609
rect 103072 67640 103100 67680
rect 103241 67677 103253 67711
rect 103287 67708 103299 67711
rect 103698 67708 103704 67720
rect 103287 67680 103704 67708
rect 103287 67677 103299 67680
rect 103241 67671 103299 67677
rect 103698 67668 103704 67680
rect 103756 67668 103762 67720
rect 108209 67711 108267 67717
rect 108209 67677 108221 67711
rect 108255 67708 108267 67711
rect 108482 67708 108488 67720
rect 108255 67680 108488 67708
rect 108255 67677 108267 67680
rect 108209 67671 108267 67677
rect 108482 67668 108488 67680
rect 108540 67668 108546 67720
rect 103330 67640 103336 67652
rect 103072 67612 103336 67640
rect 87414 67532 87420 67584
rect 87472 67532 87478 67584
rect 89070 67532 89076 67584
rect 89128 67532 89134 67584
rect 89241 67575 89299 67581
rect 89241 67541 89253 67575
rect 89287 67572 89299 67575
rect 89346 67572 89352 67584
rect 89287 67544 89352 67572
rect 89287 67541 89299 67544
rect 89241 67535 89299 67541
rect 89346 67532 89352 67544
rect 89404 67532 89410 67584
rect 95326 67532 95332 67584
rect 95384 67572 95390 67584
rect 95421 67575 95479 67581
rect 95421 67572 95433 67575
rect 95384 67544 95433 67572
rect 95384 67532 95390 67544
rect 95421 67541 95433 67544
rect 95467 67541 95479 67575
rect 95421 67535 95479 67541
rect 99650 67532 99656 67584
rect 99708 67572 99714 67584
rect 99837 67575 99895 67581
rect 99837 67572 99849 67575
rect 99708 67544 99849 67572
rect 99708 67532 99714 67544
rect 99837 67541 99849 67544
rect 99883 67541 99895 67575
rect 99837 67535 99895 67541
rect 100846 67532 100852 67584
rect 100904 67572 100910 67584
rect 103072 67572 103100 67612
rect 103330 67600 103336 67612
rect 103388 67600 103394 67652
rect 100904 67544 103100 67572
rect 100904 67532 100910 67544
rect 103146 67532 103152 67584
rect 103204 67532 103210 67584
rect 1104 67482 108836 67504
rect 1104 67430 4874 67482
rect 4926 67430 4938 67482
rect 4990 67430 5002 67482
rect 5054 67430 5066 67482
rect 5118 67430 5130 67482
rect 5182 67430 35594 67482
rect 35646 67430 35658 67482
rect 35710 67430 35722 67482
rect 35774 67430 35786 67482
rect 35838 67430 35850 67482
rect 35902 67430 66314 67482
rect 66366 67430 66378 67482
rect 66430 67430 66442 67482
rect 66494 67430 66506 67482
rect 66558 67430 66570 67482
rect 66622 67430 97034 67482
rect 97086 67430 97098 67482
rect 97150 67430 97162 67482
rect 97214 67430 97226 67482
rect 97278 67430 97290 67482
rect 97342 67430 108836 67482
rect 1104 67408 108836 67430
rect 86862 67328 86868 67380
rect 86920 67368 86926 67380
rect 86957 67371 87015 67377
rect 86957 67368 86969 67371
rect 86920 67340 86969 67368
rect 86920 67328 86926 67340
rect 86957 67337 86969 67340
rect 87003 67337 87015 67371
rect 86957 67331 87015 67337
rect 87414 67328 87420 67380
rect 87472 67368 87478 67380
rect 89073 67371 89131 67377
rect 89073 67368 89085 67371
rect 87472 67340 89085 67368
rect 87472 67328 87478 67340
rect 89073 67337 89085 67340
rect 89119 67337 89131 67371
rect 89073 67331 89131 67337
rect 86681 67235 86739 67241
rect 86681 67201 86693 67235
rect 86727 67232 86739 67235
rect 86880 67232 86908 67328
rect 89088 67300 89116 67331
rect 89346 67328 89352 67380
rect 89404 67368 89410 67380
rect 89533 67371 89591 67377
rect 89533 67368 89545 67371
rect 89404 67340 89545 67368
rect 89404 67328 89410 67340
rect 89533 67337 89545 67340
rect 89579 67337 89591 67371
rect 90174 67368 90180 67380
rect 89533 67331 89591 67337
rect 89824 67340 90180 67368
rect 89824 67300 89852 67340
rect 90174 67328 90180 67340
rect 90232 67368 90238 67380
rect 90821 67371 90879 67377
rect 90821 67368 90833 67371
rect 90232 67340 90833 67368
rect 90232 67328 90238 67340
rect 90821 67337 90833 67340
rect 90867 67368 90879 67371
rect 90867 67340 91232 67368
rect 90867 67337 90879 67340
rect 90821 67331 90879 67337
rect 89088 67272 89852 67300
rect 89898 67260 89904 67312
rect 89956 67300 89962 67312
rect 91005 67303 91063 67309
rect 91005 67300 91017 67303
rect 89956 67272 91017 67300
rect 89956 67260 89962 67272
rect 91005 67269 91017 67272
rect 91051 67269 91063 67303
rect 91204 67300 91232 67340
rect 92934 67328 92940 67380
rect 92992 67328 92998 67380
rect 93394 67328 93400 67380
rect 93452 67328 93458 67380
rect 95234 67328 95240 67380
rect 95292 67368 95298 67380
rect 96798 67377 96804 67380
rect 95421 67371 95479 67377
rect 95421 67368 95433 67371
rect 95292 67340 95433 67368
rect 95292 67328 95298 67340
rect 95421 67337 95433 67340
rect 95467 67337 95479 67371
rect 95421 67331 95479 67337
rect 96785 67371 96804 67377
rect 96785 67337 96797 67371
rect 96785 67331 96804 67337
rect 96798 67328 96804 67331
rect 96856 67328 96862 67380
rect 97261 67371 97319 67377
rect 97261 67368 97273 67371
rect 97000 67340 97273 67368
rect 91462 67300 91468 67312
rect 91204 67272 91468 67300
rect 91005 67263 91063 67269
rect 86727 67204 86908 67232
rect 86727 67201 86739 67204
rect 86681 67195 86739 67201
rect 89346 67192 89352 67244
rect 89404 67232 89410 67244
rect 89441 67235 89499 67241
rect 89441 67232 89453 67235
rect 89404 67204 89453 67232
rect 89404 67192 89410 67204
rect 89441 67201 89453 67204
rect 89487 67232 89499 67235
rect 89717 67235 89775 67241
rect 89717 67232 89729 67235
rect 89487 67204 89729 67232
rect 89487 67201 89499 67204
rect 89441 67195 89499 67201
rect 89717 67201 89729 67204
rect 89763 67201 89775 67235
rect 89717 67195 89775 67201
rect 90453 67235 90511 67241
rect 90453 67201 90465 67235
rect 90499 67232 90511 67235
rect 91186 67232 91192 67244
rect 90499 67204 91192 67232
rect 90499 67201 90511 67204
rect 90453 67195 90511 67201
rect 89732 67096 89760 67195
rect 91186 67192 91192 67204
rect 91244 67192 91250 67244
rect 91296 67241 91324 67272
rect 91462 67260 91468 67272
rect 91520 67260 91526 67312
rect 92566 67260 92572 67312
rect 92624 67300 92630 67312
rect 93026 67300 93032 67312
rect 92624 67272 93032 67300
rect 92624 67260 92630 67272
rect 93026 67260 93032 67272
rect 93084 67300 93090 67312
rect 93305 67303 93363 67309
rect 93305 67300 93317 67303
rect 93084 67272 93317 67300
rect 93084 67260 93090 67272
rect 93305 67269 93317 67272
rect 93351 67300 93363 67303
rect 93351 67272 93624 67300
rect 93351 67269 93363 67272
rect 93305 67263 93363 67269
rect 91281 67235 91339 67241
rect 91281 67201 91293 67235
rect 91327 67201 91339 67235
rect 91281 67195 91339 67201
rect 92750 67192 92756 67244
rect 92808 67232 92814 67244
rect 93596 67241 93624 67272
rect 92845 67235 92903 67241
rect 92845 67232 92857 67235
rect 92808 67204 92857 67232
rect 92808 67192 92814 67204
rect 92845 67201 92857 67204
rect 92891 67232 92903 67235
rect 93121 67235 93179 67241
rect 93121 67232 93133 67235
rect 92891 67204 93133 67232
rect 92891 67201 92903 67204
rect 92845 67195 92903 67201
rect 93121 67201 93133 67204
rect 93167 67232 93179 67235
rect 93397 67235 93455 67241
rect 93397 67232 93409 67235
rect 93167 67204 93409 67232
rect 93167 67201 93179 67204
rect 93121 67195 93179 67201
rect 93397 67201 93409 67204
rect 93443 67201 93455 67235
rect 93397 67195 93455 67201
rect 93581 67235 93639 67241
rect 93581 67201 93593 67235
rect 93627 67201 93639 67235
rect 93581 67195 93639 67201
rect 95329 67235 95387 67241
rect 95329 67201 95341 67235
rect 95375 67232 95387 67235
rect 95789 67235 95847 67241
rect 95789 67232 95801 67235
rect 95375 67204 95801 67232
rect 95375 67201 95387 67204
rect 95329 67195 95387 67201
rect 95789 67201 95801 67204
rect 95835 67232 95847 67235
rect 95970 67232 95976 67244
rect 95835 67204 95976 67232
rect 95835 67201 95847 67204
rect 95789 67195 95847 67201
rect 93412 67164 93440 67195
rect 95970 67192 95976 67204
rect 96028 67192 96034 67244
rect 96816 67232 96844 67328
rect 97000 67309 97028 67340
rect 97261 67337 97273 67340
rect 97307 67368 97319 67371
rect 99098 67368 99104 67380
rect 97307 67340 99104 67368
rect 97307 67337 97319 67340
rect 97261 67331 97319 67337
rect 99098 67328 99104 67340
rect 99156 67328 99162 67380
rect 99558 67328 99564 67380
rect 99616 67368 99622 67380
rect 102410 67368 102416 67380
rect 99616 67340 100156 67368
rect 99616 67328 99622 67340
rect 96985 67303 97043 67309
rect 96985 67269 96997 67303
rect 97031 67269 97043 67303
rect 96985 67263 97043 67269
rect 99484 67272 99788 67300
rect 99484 67241 99512 67272
rect 97077 67235 97135 67241
rect 97077 67232 97089 67235
rect 96816 67204 97089 67232
rect 97077 67201 97089 67204
rect 97123 67201 97135 67235
rect 97077 67195 97135 67201
rect 97353 67235 97411 67241
rect 97353 67201 97365 67235
rect 97399 67201 97411 67235
rect 97353 67195 97411 67201
rect 99469 67235 99527 67241
rect 99469 67201 99481 67235
rect 99515 67201 99527 67235
rect 99469 67195 99527 67201
rect 93765 67167 93823 67173
rect 93765 67164 93777 67167
rect 93412 67136 93777 67164
rect 93765 67133 93777 67136
rect 93811 67164 93823 67167
rect 94498 67164 94504 67176
rect 93811 67136 94504 67164
rect 93811 67133 93823 67136
rect 93765 67127 93823 67133
rect 94498 67124 94504 67136
rect 94556 67164 94562 67176
rect 94556 67136 94912 67164
rect 94556 67124 94562 67136
rect 92198 67096 92204 67108
rect 89732 67068 92204 67096
rect 92198 67056 92204 67068
rect 92256 67096 92262 67108
rect 94774 67096 94780 67108
rect 92256 67068 94780 67096
rect 92256 67056 92262 67068
rect 94774 67056 94780 67068
rect 94832 67056 94838 67108
rect 94884 67096 94912 67136
rect 95510 67124 95516 67176
rect 95568 67164 95574 67176
rect 95697 67167 95755 67173
rect 95697 67164 95709 67167
rect 95568 67136 95709 67164
rect 95568 67124 95574 67136
rect 95697 67133 95709 67136
rect 95743 67133 95755 67167
rect 95697 67127 95755 67133
rect 96890 67124 96896 67176
rect 96948 67164 96954 67176
rect 97368 67164 97396 67195
rect 99650 67192 99656 67244
rect 99708 67192 99714 67244
rect 99760 67232 99788 67272
rect 99834 67260 99840 67312
rect 99892 67300 99898 67312
rect 99929 67303 99987 67309
rect 99929 67300 99941 67303
rect 99892 67272 99941 67300
rect 99892 67260 99898 67272
rect 99929 67269 99941 67272
rect 99975 67269 99987 67303
rect 99929 67263 99987 67269
rect 100018 67260 100024 67312
rect 100076 67260 100082 67312
rect 100128 67309 100156 67340
rect 101324 67340 102416 67368
rect 101324 67312 101352 67340
rect 102410 67328 102416 67340
rect 102468 67328 102474 67380
rect 102778 67328 102784 67380
rect 102836 67368 102842 67380
rect 103057 67371 103115 67377
rect 103057 67368 103069 67371
rect 102836 67340 103069 67368
rect 102836 67328 102842 67340
rect 103057 67337 103069 67340
rect 103103 67337 103115 67371
rect 103057 67331 103115 67337
rect 100113 67303 100171 67309
rect 100113 67269 100125 67303
rect 100159 67269 100171 67303
rect 100757 67303 100815 67309
rect 100757 67300 100769 67303
rect 100113 67263 100171 67269
rect 100312 67272 100769 67300
rect 100312 67241 100340 67272
rect 100757 67269 100769 67272
rect 100803 67300 100815 67303
rect 101306 67300 101312 67312
rect 100803 67272 101312 67300
rect 100803 67269 100815 67272
rect 100757 67263 100815 67269
rect 101306 67260 101312 67272
rect 101364 67260 101370 67312
rect 101950 67300 101956 67312
rect 101692 67272 101956 67300
rect 100297 67235 100355 67241
rect 100297 67232 100309 67235
rect 99760 67204 100309 67232
rect 100297 67201 100309 67204
rect 100343 67201 100355 67235
rect 100297 67195 100355 67201
rect 100389 67235 100447 67241
rect 100389 67201 100401 67235
rect 100435 67232 100447 67235
rect 100573 67235 100631 67241
rect 100573 67232 100585 67235
rect 100435 67204 100585 67232
rect 100435 67201 100447 67204
rect 100389 67195 100447 67201
rect 100573 67201 100585 67204
rect 100619 67201 100631 67235
rect 100573 67195 100631 67201
rect 96948 67136 97396 67164
rect 99668 67164 99696 67192
rect 100110 67164 100116 67176
rect 99668 67136 100116 67164
rect 96948 67124 96954 67136
rect 100110 67124 100116 67136
rect 100168 67164 100174 67176
rect 100404 67164 100432 67195
rect 100846 67192 100852 67244
rect 100904 67232 100910 67244
rect 101692 67241 101720 67272
rect 101950 67260 101956 67272
rect 102008 67300 102014 67312
rect 102505 67303 102563 67309
rect 102505 67300 102517 67303
rect 102008 67272 102517 67300
rect 102008 67260 102014 67272
rect 102505 67269 102517 67272
rect 102551 67269 102563 67303
rect 102505 67263 102563 67269
rect 102870 67260 102876 67312
rect 102928 67260 102934 67312
rect 103209 67303 103267 67309
rect 103209 67300 103221 67303
rect 102980 67272 103221 67300
rect 102980 67244 103008 67272
rect 103209 67269 103221 67272
rect 103255 67269 103267 67303
rect 103209 67263 103267 67269
rect 103425 67303 103483 67309
rect 103425 67269 103437 67303
rect 103471 67300 103483 67303
rect 103514 67300 103520 67312
rect 103471 67272 103520 67300
rect 103471 67269 103483 67272
rect 103425 67263 103483 67269
rect 101493 67235 101551 67241
rect 101493 67232 101505 67235
rect 100904 67204 101505 67232
rect 100904 67192 100910 67204
rect 101493 67201 101505 67204
rect 101539 67201 101551 67235
rect 101493 67195 101551 67201
rect 101677 67235 101735 67241
rect 101677 67201 101689 67235
rect 101723 67201 101735 67235
rect 101677 67195 101735 67201
rect 101766 67192 101772 67244
rect 101824 67192 101830 67244
rect 101861 67235 101919 67241
rect 101861 67201 101873 67235
rect 101907 67201 101919 67235
rect 102226 67232 102232 67244
rect 101861 67195 101919 67201
rect 102152 67204 102232 67232
rect 100168 67136 100432 67164
rect 100168 67124 100174 67136
rect 100938 67124 100944 67176
rect 100996 67164 101002 67176
rect 101784 67164 101812 67192
rect 100996 67136 101812 67164
rect 100996 67124 101002 67136
rect 100570 67096 100576 67108
rect 94884 67068 100576 67096
rect 100570 67056 100576 67068
rect 100628 67056 100634 67108
rect 101876 67096 101904 67195
rect 102152 67173 102180 67204
rect 102226 67192 102232 67204
rect 102284 67192 102290 67244
rect 102594 67192 102600 67244
rect 102652 67232 102658 67244
rect 102689 67235 102747 67241
rect 102689 67232 102701 67235
rect 102652 67204 102701 67232
rect 102652 67192 102658 67204
rect 102689 67201 102701 67204
rect 102735 67201 102747 67235
rect 102689 67195 102747 67201
rect 102962 67192 102968 67244
rect 103020 67192 103026 67244
rect 103440 67232 103468 67263
rect 103514 67260 103520 67272
rect 103572 67300 103578 67312
rect 103974 67300 103980 67312
rect 103572 67272 103980 67300
rect 103572 67260 103578 67272
rect 103974 67260 103980 67272
rect 104032 67260 104038 67312
rect 103072 67204 103468 67232
rect 102137 67167 102195 67173
rect 102137 67133 102149 67167
rect 102183 67133 102195 67167
rect 103072 67164 103100 67204
rect 103698 67192 103704 67244
rect 103756 67192 103762 67244
rect 102137 67127 102195 67133
rect 102244 67136 103100 67164
rect 102244 67096 102272 67136
rect 103146 67124 103152 67176
rect 103204 67164 103210 67176
rect 103885 67167 103943 67173
rect 103885 67164 103897 67167
rect 103204 67136 103897 67164
rect 103204 67124 103210 67136
rect 103885 67133 103897 67136
rect 103931 67133 103943 67167
rect 103885 67127 103943 67133
rect 103517 67099 103575 67105
rect 103517 67096 103529 67099
rect 101876 67068 102272 67096
rect 102336 67068 103529 67096
rect 86770 66988 86776 67040
rect 86828 66988 86834 67040
rect 89806 66988 89812 67040
rect 89864 67028 89870 67040
rect 90361 67031 90419 67037
rect 90361 67028 90373 67031
rect 89864 67000 90373 67028
rect 89864 66988 89870 67000
rect 90361 66997 90373 67000
rect 90407 66997 90419 67031
rect 90361 66991 90419 66997
rect 96154 66988 96160 67040
rect 96212 67028 96218 67040
rect 96617 67031 96675 67037
rect 96617 67028 96629 67031
rect 96212 67000 96629 67028
rect 96212 66988 96218 67000
rect 96617 66997 96629 67000
rect 96663 66997 96675 67031
rect 96617 66991 96675 66997
rect 96801 67031 96859 67037
rect 96801 66997 96813 67031
rect 96847 67028 96859 67031
rect 96890 67028 96896 67040
rect 96847 67000 96896 67028
rect 96847 66997 96859 67000
rect 96801 66991 96859 66997
rect 96890 66988 96896 67000
rect 96948 66988 96954 67040
rect 97074 66988 97080 67040
rect 97132 66988 97138 67040
rect 100662 66988 100668 67040
rect 100720 67028 100726 67040
rect 100941 67031 100999 67037
rect 100941 67028 100953 67031
rect 100720 67000 100953 67028
rect 100720 66988 100726 67000
rect 100941 66997 100953 67000
rect 100987 66997 100999 67031
rect 100941 66991 100999 66997
rect 102042 66988 102048 67040
rect 102100 67028 102106 67040
rect 102336 67028 102364 67068
rect 103517 67065 103529 67068
rect 103563 67065 103575 67099
rect 103517 67059 103575 67065
rect 102100 67000 102364 67028
rect 102100 66988 102106 67000
rect 102870 66988 102876 67040
rect 102928 67028 102934 67040
rect 103241 67031 103299 67037
rect 103241 67028 103253 67031
rect 102928 67000 103253 67028
rect 102928 66988 102934 67000
rect 103241 66997 103253 67000
rect 103287 66997 103299 67031
rect 103241 66991 103299 66997
rect 1104 66938 108836 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 96374 66938
rect 96426 66886 96438 66938
rect 96490 66886 96502 66938
rect 96554 66886 96566 66938
rect 96618 66886 96630 66938
rect 96682 66886 108836 66938
rect 1104 66864 108836 66886
rect 89438 66784 89444 66836
rect 89496 66784 89502 66836
rect 89806 66784 89812 66836
rect 89864 66784 89870 66836
rect 90634 66784 90640 66836
rect 90692 66824 90698 66836
rect 91186 66824 91192 66836
rect 90692 66796 91192 66824
rect 90692 66784 90698 66796
rect 91186 66784 91192 66796
rect 91244 66824 91250 66836
rect 92385 66827 92443 66833
rect 92385 66824 92397 66827
rect 91244 66796 92397 66824
rect 91244 66784 91250 66796
rect 92385 66793 92397 66796
rect 92431 66793 92443 66827
rect 92385 66787 92443 66793
rect 92474 66784 92480 66836
rect 92532 66824 92538 66836
rect 92569 66827 92627 66833
rect 92569 66824 92581 66827
rect 92532 66796 92581 66824
rect 92532 66784 92538 66796
rect 92569 66793 92581 66796
rect 92615 66793 92627 66827
rect 92569 66787 92627 66793
rect 95694 66784 95700 66836
rect 95752 66824 95758 66836
rect 95789 66827 95847 66833
rect 95789 66824 95801 66827
rect 95752 66796 95801 66824
rect 95752 66784 95758 66796
rect 95789 66793 95801 66796
rect 95835 66793 95847 66827
rect 95789 66787 95847 66793
rect 95970 66784 95976 66836
rect 96028 66784 96034 66836
rect 99745 66827 99803 66833
rect 99745 66793 99757 66827
rect 99791 66824 99803 66827
rect 99926 66824 99932 66836
rect 99791 66796 99932 66824
rect 99791 66793 99803 66796
rect 99745 66787 99803 66793
rect 99926 66784 99932 66796
rect 99984 66784 99990 66836
rect 100110 66784 100116 66836
rect 100168 66824 100174 66836
rect 100205 66827 100263 66833
rect 100205 66824 100217 66827
rect 100168 66796 100217 66824
rect 100168 66784 100174 66796
rect 100205 66793 100217 66796
rect 100251 66793 100263 66827
rect 100205 66787 100263 66793
rect 100570 66784 100576 66836
rect 100628 66824 100634 66836
rect 102134 66824 102140 66836
rect 100628 66796 102140 66824
rect 100628 66784 100634 66796
rect 102134 66784 102140 66796
rect 102192 66784 102198 66836
rect 102597 66827 102655 66833
rect 102597 66793 102609 66827
rect 102643 66824 102655 66827
rect 103146 66824 103152 66836
rect 102643 66796 103152 66824
rect 102643 66793 102655 66796
rect 102597 66787 102655 66793
rect 103146 66784 103152 66796
rect 103204 66784 103210 66836
rect 103698 66784 103704 66836
rect 103756 66824 103762 66836
rect 103793 66827 103851 66833
rect 103793 66824 103805 66827
rect 103756 66796 103805 66824
rect 103756 66784 103762 66796
rect 103793 66793 103805 66796
rect 103839 66793 103851 66827
rect 103793 66787 103851 66793
rect 90177 66759 90235 66765
rect 90177 66756 90189 66759
rect 89686 66728 90189 66756
rect 87233 66691 87291 66697
rect 87233 66657 87245 66691
rect 87279 66688 87291 66691
rect 89686 66688 89714 66728
rect 90177 66725 90189 66728
rect 90223 66756 90235 66759
rect 92014 66756 92020 66768
rect 90223 66728 92020 66756
rect 90223 66725 90235 66728
rect 90177 66719 90235 66725
rect 92014 66716 92020 66728
rect 92072 66756 92078 66768
rect 92109 66759 92167 66765
rect 92109 66756 92121 66759
rect 92072 66728 92121 66756
rect 92072 66716 92078 66728
rect 92109 66725 92121 66728
rect 92155 66756 92167 66759
rect 92492 66756 92520 66784
rect 92155 66728 92520 66756
rect 92155 66725 92167 66728
rect 92109 66719 92167 66725
rect 97626 66716 97632 66768
rect 97684 66716 97690 66768
rect 99834 66756 99840 66768
rect 99392 66728 99840 66756
rect 87279 66660 89714 66688
rect 87279 66657 87291 66660
rect 87233 66651 87291 66657
rect 91462 66648 91468 66700
rect 91520 66688 91526 66700
rect 95053 66691 95111 66697
rect 95053 66688 95065 66691
rect 91520 66660 95065 66688
rect 91520 66648 91526 66660
rect 95053 66657 95065 66660
rect 95099 66688 95111 66691
rect 95234 66688 95240 66700
rect 95099 66660 95240 66688
rect 95099 66657 95111 66660
rect 95053 66651 95111 66657
rect 95234 66648 95240 66660
rect 95292 66688 95298 66700
rect 96062 66688 96068 66700
rect 95292 66660 96068 66688
rect 95292 66648 95298 66660
rect 96062 66648 96068 66660
rect 96120 66648 96126 66700
rect 96154 66648 96160 66700
rect 96212 66648 96218 66700
rect 97353 66691 97411 66697
rect 97353 66657 97365 66691
rect 97399 66688 97411 66691
rect 97442 66688 97448 66700
rect 97399 66660 97448 66688
rect 97399 66657 97411 66660
rect 97353 66651 97411 66657
rect 97442 66648 97448 66660
rect 97500 66648 97506 66700
rect 98546 66688 98552 66700
rect 98380 66660 98552 66688
rect 84933 66623 84991 66629
rect 84933 66589 84945 66623
rect 84979 66620 84991 66623
rect 85209 66623 85267 66629
rect 85209 66620 85221 66623
rect 84979 66592 85221 66620
rect 84979 66589 84991 66592
rect 84933 66583 84991 66589
rect 85209 66589 85221 66592
rect 85255 66620 85267 66623
rect 85390 66620 85396 66632
rect 85255 66592 85396 66620
rect 85255 66589 85267 66592
rect 85209 66583 85267 66589
rect 85390 66580 85396 66592
rect 85448 66580 85454 66632
rect 86770 66580 86776 66632
rect 86828 66620 86834 66632
rect 86828 66592 87906 66620
rect 86828 66580 86834 66592
rect 89254 66580 89260 66632
rect 89312 66580 89318 66632
rect 89346 66580 89352 66632
rect 89404 66580 89410 66632
rect 89533 66623 89591 66629
rect 89533 66589 89545 66623
rect 89579 66620 89591 66623
rect 89898 66620 89904 66632
rect 89579 66592 89904 66620
rect 89579 66589 89591 66592
rect 89533 66583 89591 66589
rect 89898 66580 89904 66592
rect 89956 66580 89962 66632
rect 95602 66580 95608 66632
rect 95660 66620 95666 66632
rect 95973 66623 96031 66629
rect 95973 66620 95985 66623
rect 95660 66592 95985 66620
rect 95660 66580 95666 66592
rect 95973 66589 95985 66592
rect 96019 66589 96031 66623
rect 95973 66583 96031 66589
rect 96249 66623 96307 66629
rect 96249 66589 96261 66623
rect 96295 66620 96307 66623
rect 97074 66620 97080 66632
rect 96295 66592 97080 66620
rect 96295 66589 96307 66592
rect 96249 66583 96307 66589
rect 97074 66580 97080 66592
rect 97132 66580 97138 66632
rect 97261 66623 97319 66629
rect 97261 66589 97273 66623
rect 97307 66620 97319 66623
rect 98270 66620 98276 66632
rect 97307 66592 98276 66620
rect 97307 66589 97319 66592
rect 97261 66583 97319 66589
rect 98270 66580 98276 66592
rect 98328 66580 98334 66632
rect 98380 66629 98408 66660
rect 98546 66648 98552 66660
rect 98604 66648 98610 66700
rect 99392 66697 99420 66728
rect 99834 66716 99840 66728
rect 99892 66716 99898 66768
rect 101858 66716 101864 66768
rect 101916 66716 101922 66768
rect 102778 66716 102784 66768
rect 102836 66756 102842 66768
rect 102836 66728 104112 66756
rect 102836 66716 102842 66728
rect 99377 66691 99435 66697
rect 99377 66657 99389 66691
rect 99423 66657 99435 66691
rect 99377 66651 99435 66657
rect 99466 66648 99472 66700
rect 99524 66648 99530 66700
rect 99558 66648 99564 66700
rect 99616 66688 99622 66700
rect 99616 66660 99880 66688
rect 99616 66648 99622 66660
rect 98365 66623 98423 66629
rect 98365 66589 98377 66623
rect 98411 66589 98423 66623
rect 98365 66583 98423 66589
rect 98730 66580 98736 66632
rect 98788 66580 98794 66632
rect 99101 66623 99159 66629
rect 99101 66589 99113 66623
rect 99147 66620 99159 66623
rect 99576 66620 99604 66648
rect 99147 66592 99604 66620
rect 99147 66589 99159 66592
rect 99101 66583 99159 66589
rect 99650 66580 99656 66632
rect 99708 66580 99714 66632
rect 99852 66629 99880 66660
rect 100478 66648 100484 66700
rect 100536 66688 100542 66700
rect 100757 66691 100815 66697
rect 100757 66688 100769 66691
rect 100536 66660 100769 66688
rect 100536 66648 100542 66660
rect 100757 66657 100769 66660
rect 100803 66657 100815 66691
rect 100757 66651 100815 66657
rect 100846 66648 100852 66700
rect 100904 66688 100910 66700
rect 101677 66691 101735 66697
rect 101677 66688 101689 66691
rect 100904 66660 101689 66688
rect 100904 66648 100910 66660
rect 101677 66657 101689 66660
rect 101723 66657 101735 66691
rect 101677 66651 101735 66657
rect 102137 66691 102195 66697
rect 102137 66657 102149 66691
rect 102183 66688 102195 66691
rect 102226 66688 102232 66700
rect 102183 66660 102232 66688
rect 102183 66657 102195 66660
rect 102137 66651 102195 66657
rect 102226 66648 102232 66660
rect 102284 66648 102290 66700
rect 103238 66648 103244 66700
rect 103296 66648 103302 66700
rect 99837 66623 99895 66629
rect 99837 66589 99849 66623
rect 99883 66620 99895 66623
rect 99929 66623 99987 66629
rect 99929 66620 99941 66623
rect 99883 66592 99941 66620
rect 99883 66589 99895 66592
rect 99837 66583 99895 66589
rect 99929 66589 99941 66592
rect 99975 66589 99987 66623
rect 99929 66583 99987 66589
rect 100113 66623 100171 66629
rect 100113 66589 100125 66623
rect 100159 66620 100171 66623
rect 100662 66620 100668 66632
rect 100159 66592 100668 66620
rect 100159 66589 100171 66592
rect 100113 66583 100171 66589
rect 100662 66580 100668 66592
rect 100720 66580 100726 66632
rect 102778 66580 102784 66632
rect 102836 66580 102842 66632
rect 102870 66580 102876 66632
rect 102928 66580 102934 66632
rect 102965 66623 103023 66629
rect 102965 66589 102977 66623
rect 103011 66620 103023 66623
rect 103256 66620 103284 66648
rect 103011 66592 103284 66620
rect 103011 66589 103023 66592
rect 102965 66583 103023 66589
rect 103330 66580 103336 66632
rect 103388 66580 103394 66632
rect 104084 66629 104112 66728
rect 103977 66623 104035 66629
rect 103977 66620 103989 66623
rect 103440 66592 103989 66620
rect 85025 66555 85083 66561
rect 85025 66521 85037 66555
rect 85071 66552 85083 66555
rect 86862 66552 86868 66564
rect 85071 66524 86868 66552
rect 85071 66521 85083 66524
rect 85025 66515 85083 66521
rect 86862 66512 86868 66524
rect 86920 66512 86926 66564
rect 88981 66555 89039 66561
rect 88981 66521 88993 66555
rect 89027 66552 89039 66555
rect 89027 66524 89668 66552
rect 89027 66521 89039 66524
rect 88981 66515 89039 66521
rect 87138 66444 87144 66496
rect 87196 66484 87202 66496
rect 88242 66484 88248 66496
rect 87196 66456 88248 66484
rect 87196 66444 87202 66456
rect 88242 66444 88248 66456
rect 88300 66444 88306 66496
rect 89640 66493 89668 66524
rect 89990 66512 89996 66564
rect 90048 66512 90054 66564
rect 92290 66512 92296 66564
rect 92348 66552 92354 66564
rect 92750 66552 92756 66564
rect 92348 66524 92756 66552
rect 92348 66512 92354 66524
rect 92750 66512 92756 66524
rect 92808 66512 92814 66564
rect 94501 66555 94559 66561
rect 94501 66521 94513 66555
rect 94547 66552 94559 66555
rect 94774 66552 94780 66564
rect 94547 66524 94780 66552
rect 94547 66521 94559 66524
rect 94501 66515 94559 66521
rect 94774 66512 94780 66524
rect 94832 66552 94838 66564
rect 97626 66552 97632 66564
rect 94832 66524 97632 66552
rect 94832 66512 94838 66524
rect 97626 66512 97632 66524
rect 97684 66512 97690 66564
rect 101674 66512 101680 66564
rect 101732 66552 101738 66564
rect 102888 66552 102916 66580
rect 103440 66552 103468 66592
rect 103977 66589 103989 66592
rect 104023 66589 104035 66623
rect 103977 66583 104035 66589
rect 104069 66623 104127 66629
rect 104069 66589 104081 66623
rect 104115 66589 104127 66623
rect 104069 66583 104127 66589
rect 104345 66623 104403 66629
rect 104345 66589 104357 66623
rect 104391 66620 104403 66623
rect 104805 66623 104863 66629
rect 104805 66620 104817 66623
rect 104391 66592 104817 66620
rect 104391 66589 104403 66592
rect 104345 66583 104403 66589
rect 104805 66589 104817 66592
rect 104851 66589 104863 66623
rect 104805 66583 104863 66589
rect 101732 66524 103468 66552
rect 103716 66524 104020 66552
rect 101732 66512 101738 66524
rect 103716 66496 103744 66524
rect 89625 66487 89683 66493
rect 89625 66453 89637 66487
rect 89671 66453 89683 66487
rect 89625 66447 89683 66453
rect 89793 66487 89851 66493
rect 89793 66453 89805 66487
rect 89839 66484 89851 66487
rect 89898 66484 89904 66496
rect 89839 66456 89904 66484
rect 89839 66453 89851 66456
rect 89793 66447 89851 66453
rect 89898 66444 89904 66456
rect 89956 66444 89962 66496
rect 92566 66493 92572 66496
rect 92553 66487 92572 66493
rect 92553 66453 92565 66487
rect 92553 66447 92572 66453
rect 92566 66444 92572 66447
rect 92624 66444 92630 66496
rect 95418 66444 95424 66496
rect 95476 66484 95482 66496
rect 95878 66484 95884 66496
rect 95476 66456 95884 66484
rect 95476 66444 95482 66456
rect 95878 66444 95884 66456
rect 95936 66444 95942 66496
rect 99926 66444 99932 66496
rect 99984 66444 99990 66496
rect 100570 66444 100576 66496
rect 100628 66444 100634 66496
rect 100665 66487 100723 66493
rect 100665 66453 100677 66487
rect 100711 66484 100723 66487
rect 101306 66484 101312 66496
rect 100711 66456 101312 66484
rect 100711 66453 100723 66456
rect 100665 66447 100723 66453
rect 101306 66444 101312 66456
rect 101364 66444 101370 66496
rect 103698 66444 103704 66496
rect 103756 66444 103762 66496
rect 103992 66484 104020 66524
rect 104158 66512 104164 66564
rect 104216 66512 104222 66564
rect 104437 66555 104495 66561
rect 104437 66521 104449 66555
rect 104483 66521 104495 66555
rect 104437 66515 104495 66521
rect 104452 66484 104480 66515
rect 104618 66512 104624 66564
rect 104676 66512 104682 66564
rect 103992 66456 104480 66484
rect 1104 66394 108836 66416
rect 1104 66342 4874 66394
rect 4926 66342 4938 66394
rect 4990 66342 5002 66394
rect 5054 66342 5066 66394
rect 5118 66342 5130 66394
rect 5182 66342 35594 66394
rect 35646 66342 35658 66394
rect 35710 66342 35722 66394
rect 35774 66342 35786 66394
rect 35838 66342 35850 66394
rect 35902 66342 66314 66394
rect 66366 66342 66378 66394
rect 66430 66342 66442 66394
rect 66494 66342 66506 66394
rect 66558 66342 66570 66394
rect 66622 66342 97034 66394
rect 97086 66342 97098 66394
rect 97150 66342 97162 66394
rect 97214 66342 97226 66394
rect 97278 66342 97290 66394
rect 97342 66342 106658 66394
rect 106710 66342 106722 66394
rect 106774 66342 106786 66394
rect 106838 66342 106850 66394
rect 106902 66342 106914 66394
rect 106966 66342 108836 66394
rect 1104 66320 108836 66342
rect 87138 66280 87144 66292
rect 86696 66252 87144 66280
rect 9490 66172 9496 66224
rect 9548 66212 9554 66224
rect 13814 66212 13820 66224
rect 9548 66184 13820 66212
rect 9548 66172 9554 66184
rect 13814 66172 13820 66184
rect 13872 66172 13878 66224
rect 68646 66172 68652 66224
rect 68704 66172 68710 66224
rect 73154 66172 73160 66224
rect 73212 66212 73218 66224
rect 73341 66215 73399 66221
rect 73341 66212 73353 66215
rect 73212 66184 73353 66212
rect 73212 66172 73218 66184
rect 73341 66181 73353 66184
rect 73387 66181 73399 66215
rect 73341 66175 73399 66181
rect 74169 66215 74227 66221
rect 74169 66181 74181 66215
rect 74215 66212 74227 66215
rect 74350 66212 74356 66224
rect 74215 66184 74356 66212
rect 74215 66181 74227 66184
rect 74169 66175 74227 66181
rect 74350 66172 74356 66184
rect 74408 66172 74414 66224
rect 86037 66215 86095 66221
rect 86037 66181 86049 66215
rect 86083 66212 86095 66215
rect 86696 66212 86724 66252
rect 87138 66240 87144 66252
rect 87196 66240 87202 66292
rect 88610 66240 88616 66292
rect 88668 66280 88674 66292
rect 89257 66283 89315 66289
rect 89257 66280 89269 66283
rect 88668 66252 89269 66280
rect 88668 66240 88674 66252
rect 89257 66249 89269 66252
rect 89303 66280 89315 66283
rect 89346 66280 89352 66292
rect 89303 66252 89352 66280
rect 89303 66249 89315 66252
rect 89257 66243 89315 66249
rect 89346 66240 89352 66252
rect 89404 66240 89410 66292
rect 89898 66240 89904 66292
rect 89956 66280 89962 66292
rect 92017 66283 92075 66289
rect 89956 66252 91692 66280
rect 89956 66240 89962 66252
rect 86083 66184 86724 66212
rect 87969 66215 88027 66221
rect 86083 66181 86095 66184
rect 86037 66175 86095 66181
rect 87969 66181 87981 66215
rect 88015 66212 88027 66215
rect 89070 66212 89076 66224
rect 88015 66184 89076 66212
rect 88015 66181 88027 66184
rect 87969 66175 88027 66181
rect 89070 66172 89076 66184
rect 89128 66172 89134 66224
rect 89714 66172 89720 66224
rect 89772 66212 89778 66224
rect 90269 66215 90327 66221
rect 90269 66212 90281 66215
rect 89772 66184 90281 66212
rect 89772 66172 89778 66184
rect 90269 66181 90281 66184
rect 90315 66181 90327 66215
rect 90269 66175 90327 66181
rect 90634 66172 90640 66224
rect 90692 66212 90698 66224
rect 91664 66221 91692 66252
rect 92017 66249 92029 66283
rect 92063 66280 92075 66283
rect 92290 66280 92296 66292
rect 92063 66252 92296 66280
rect 92063 66249 92075 66252
rect 92017 66243 92075 66249
rect 92290 66240 92296 66252
rect 92348 66240 92354 66292
rect 95418 66240 95424 66292
rect 95476 66289 95482 66292
rect 95476 66283 95495 66289
rect 95483 66249 95495 66283
rect 95476 66243 95495 66249
rect 95476 66240 95482 66243
rect 95602 66240 95608 66292
rect 95660 66240 95666 66292
rect 95786 66240 95792 66292
rect 95844 66240 95850 66292
rect 97169 66283 97227 66289
rect 97169 66249 97181 66283
rect 97215 66280 97227 66283
rect 97442 66280 97448 66292
rect 97215 66252 97448 66280
rect 97215 66249 97227 66252
rect 97169 66243 97227 66249
rect 97442 66240 97448 66252
rect 97500 66240 97506 66292
rect 97626 66240 97632 66292
rect 97684 66280 97690 66292
rect 103974 66280 103980 66292
rect 97684 66252 103980 66280
rect 97684 66240 97690 66252
rect 103974 66240 103980 66252
rect 104032 66240 104038 66292
rect 104069 66283 104127 66289
rect 104069 66249 104081 66283
rect 104115 66280 104127 66283
rect 104158 66280 104164 66292
rect 104115 66252 104164 66280
rect 104115 66249 104127 66252
rect 104069 66243 104127 66249
rect 104158 66240 104164 66252
rect 104216 66240 104222 66292
rect 91649 66215 91707 66221
rect 90692 66184 90864 66212
rect 90692 66172 90698 66184
rect 86862 66104 86868 66156
rect 86920 66104 86926 66156
rect 88242 66104 88248 66156
rect 88300 66144 88306 66156
rect 89254 66144 89260 66156
rect 88300 66116 89260 66144
rect 88300 66104 88306 66116
rect 89254 66104 89260 66116
rect 89312 66104 89318 66156
rect 90174 66104 90180 66156
rect 90232 66144 90238 66156
rect 90453 66147 90511 66153
rect 90453 66144 90465 66147
rect 90232 66116 90465 66144
rect 90232 66104 90238 66116
rect 90453 66113 90465 66116
rect 90499 66144 90511 66147
rect 90726 66144 90732 66156
rect 90499 66116 90732 66144
rect 90499 66113 90511 66116
rect 90453 66107 90511 66113
rect 90726 66104 90732 66116
rect 90784 66104 90790 66156
rect 90836 66150 90864 66184
rect 91649 66181 91661 66215
rect 91695 66181 91707 66215
rect 91649 66175 91707 66181
rect 94240 66184 94912 66212
rect 90913 66150 90971 66153
rect 90836 66147 90971 66150
rect 90836 66122 90925 66147
rect 90913 66113 90925 66122
rect 90959 66113 90971 66147
rect 90913 66107 90971 66113
rect 91833 66147 91891 66153
rect 91833 66113 91845 66147
rect 91879 66113 91891 66147
rect 91833 66107 91891 66113
rect 92109 66147 92167 66153
rect 92109 66113 92121 66147
rect 92155 66144 92167 66147
rect 92566 66144 92572 66156
rect 92155 66116 92572 66144
rect 92155 66113 92167 66116
rect 92109 66107 92167 66113
rect 86221 66079 86279 66085
rect 86221 66045 86233 66079
rect 86267 66076 86279 66079
rect 88610 66076 88616 66088
rect 86267 66048 88616 66076
rect 86267 66045 86279 66048
rect 86221 66039 86279 66045
rect 88610 66036 88616 66048
rect 88668 66036 88674 66088
rect 90818 66036 90824 66088
rect 90876 66036 90882 66088
rect 91465 66079 91523 66085
rect 91465 66045 91477 66079
rect 91511 66076 91523 66079
rect 91848 66076 91876 66107
rect 92566 66104 92572 66116
rect 92624 66104 92630 66156
rect 93765 66147 93823 66153
rect 93765 66113 93777 66147
rect 93811 66144 93823 66147
rect 94130 66144 94136 66156
rect 93811 66116 94136 66144
rect 93811 66113 93823 66116
rect 93765 66107 93823 66113
rect 92382 66076 92388 66088
rect 91511 66048 92388 66076
rect 91511 66045 91523 66048
rect 91465 66039 91523 66045
rect 92382 66036 92388 66048
rect 92440 66076 92446 66088
rect 93780 66076 93808 66107
rect 94130 66104 94136 66116
rect 94188 66104 94194 66156
rect 94240 66085 94268 66184
rect 94774 66104 94780 66156
rect 94832 66104 94838 66156
rect 94884 66144 94912 66184
rect 95234 66172 95240 66224
rect 95292 66172 95298 66224
rect 95878 66212 95884 66224
rect 95804 66184 95884 66212
rect 95326 66144 95332 66156
rect 94884 66116 95332 66144
rect 95326 66104 95332 66116
rect 95384 66104 95390 66156
rect 95697 66147 95755 66153
rect 95697 66113 95709 66147
rect 95743 66144 95755 66147
rect 95804 66144 95832 66184
rect 95878 66172 95884 66184
rect 95936 66212 95942 66224
rect 96706 66212 96712 66224
rect 95936 66184 96712 66212
rect 95936 66172 95942 66184
rect 96706 66172 96712 66184
rect 96764 66172 96770 66224
rect 100754 66212 100760 66224
rect 96908 66184 100760 66212
rect 95743 66116 95832 66144
rect 95973 66147 96031 66153
rect 95743 66113 95755 66116
rect 95697 66107 95755 66113
rect 95973 66113 95985 66147
rect 96019 66144 96031 66147
rect 96062 66144 96068 66156
rect 96019 66116 96068 66144
rect 96019 66113 96031 66116
rect 95973 66107 96031 66113
rect 96062 66104 96068 66116
rect 96120 66144 96126 66156
rect 96908 66153 96936 66184
rect 100754 66172 100760 66184
rect 100812 66212 100818 66224
rect 100812 66184 101260 66212
rect 100812 66172 100818 66184
rect 96893 66147 96951 66153
rect 96120 66116 96660 66144
rect 96120 66104 96126 66116
rect 92440 66048 93808 66076
rect 94225 66079 94283 66085
rect 92440 66036 92446 66048
rect 94225 66045 94237 66079
rect 94271 66045 94283 66079
rect 94225 66039 94283 66045
rect 94869 66079 94927 66085
rect 94869 66045 94881 66079
rect 94915 66076 94927 66079
rect 94915 66048 96568 66076
rect 94915 66045 94927 66048
rect 94869 66039 94927 66045
rect 89254 65968 89260 66020
rect 89312 66008 89318 66020
rect 95878 66008 95884 66020
rect 89312 65980 95884 66008
rect 89312 65968 89318 65980
rect 95878 65968 95884 65980
rect 95936 66008 95942 66020
rect 96540 66017 96568 66048
rect 96249 66011 96307 66017
rect 96249 66008 96261 66011
rect 95936 65980 96261 66008
rect 95936 65968 95942 65980
rect 96249 65977 96261 65980
rect 96295 65977 96307 66011
rect 96249 65971 96307 65977
rect 96525 66011 96583 66017
rect 96525 65977 96537 66011
rect 96571 65977 96583 66011
rect 96525 65971 96583 65977
rect 88242 65900 88248 65952
rect 88300 65940 88306 65952
rect 88337 65943 88395 65949
rect 88337 65940 88349 65943
rect 88300 65912 88349 65940
rect 88300 65900 88306 65912
rect 88337 65909 88349 65912
rect 88383 65909 88395 65943
rect 88337 65903 88395 65909
rect 90726 65900 90732 65952
rect 90784 65940 90790 65952
rect 91005 65943 91063 65949
rect 91005 65940 91017 65943
rect 90784 65912 91017 65940
rect 90784 65900 90790 65912
rect 91005 65909 91017 65912
rect 91051 65909 91063 65943
rect 91005 65903 91063 65909
rect 94406 65900 94412 65952
rect 94464 65900 94470 65952
rect 94958 65900 94964 65952
rect 95016 65940 95022 65952
rect 95053 65943 95111 65949
rect 95053 65940 95065 65943
rect 95016 65912 95065 65940
rect 95016 65900 95022 65912
rect 95053 65909 95065 65912
rect 95099 65909 95111 65943
rect 95053 65903 95111 65909
rect 95421 65943 95479 65949
rect 95421 65909 95433 65943
rect 95467 65940 95479 65943
rect 95786 65940 95792 65952
rect 95467 65912 95792 65940
rect 95467 65909 95479 65912
rect 95421 65903 95479 65909
rect 95786 65900 95792 65912
rect 95844 65900 95850 65952
rect 95970 65900 95976 65952
rect 96028 65900 96034 65952
rect 96157 65943 96215 65949
rect 96157 65909 96169 65943
rect 96203 65940 96215 65943
rect 96632 65940 96660 66116
rect 96893 66113 96905 66147
rect 96939 66113 96951 66147
rect 96893 66107 96951 66113
rect 97534 66104 97540 66156
rect 97592 66104 97598 66156
rect 98546 66104 98552 66156
rect 98604 66104 98610 66156
rect 98730 66104 98736 66156
rect 98788 66104 98794 66156
rect 99285 66147 99343 66153
rect 99285 66113 99297 66147
rect 99331 66144 99343 66147
rect 99374 66144 99380 66156
rect 99331 66116 99380 66144
rect 99331 66113 99343 66116
rect 99285 66107 99343 66113
rect 99374 66104 99380 66116
rect 99432 66144 99438 66156
rect 99650 66144 99656 66156
rect 99432 66116 99656 66144
rect 99432 66104 99438 66116
rect 99650 66104 99656 66116
rect 99708 66104 99714 66156
rect 100389 66147 100447 66153
rect 100389 66113 100401 66147
rect 100435 66144 100447 66147
rect 100846 66144 100852 66156
rect 100435 66116 100852 66144
rect 100435 66113 100447 66116
rect 100389 66107 100447 66113
rect 100846 66104 100852 66116
rect 100904 66104 100910 66156
rect 96985 66079 97043 66085
rect 96985 66076 96997 66079
rect 96908 66048 96997 66076
rect 96908 66020 96936 66048
rect 96985 66045 96997 66048
rect 97031 66045 97043 66079
rect 96985 66039 97043 66045
rect 97629 66079 97687 66085
rect 97629 66045 97641 66079
rect 97675 66076 97687 66079
rect 97902 66076 97908 66088
rect 97675 66048 97908 66076
rect 97675 66045 97687 66048
rect 97629 66039 97687 66045
rect 97902 66036 97908 66048
rect 97960 66036 97966 66088
rect 98365 66079 98423 66085
rect 98365 66045 98377 66079
rect 98411 66076 98423 66079
rect 98748 66076 98776 66104
rect 98411 66048 98776 66076
rect 99193 66079 99251 66085
rect 98411 66045 98423 66048
rect 98365 66039 98423 66045
rect 99193 66045 99205 66079
rect 99239 66076 99251 66079
rect 99926 66076 99932 66088
rect 99239 66048 99932 66076
rect 99239 66045 99251 66048
rect 99193 66039 99251 66045
rect 99926 66036 99932 66048
rect 99984 66036 99990 66088
rect 100294 66036 100300 66088
rect 100352 66036 100358 66088
rect 101232 66076 101260 66184
rect 101306 66172 101312 66224
rect 101364 66172 101370 66224
rect 102778 66212 102784 66224
rect 102428 66184 102784 66212
rect 101401 66147 101459 66153
rect 101401 66113 101413 66147
rect 101447 66144 101459 66147
rect 101677 66147 101735 66153
rect 101677 66144 101689 66147
rect 101447 66116 101689 66144
rect 101447 66113 101459 66116
rect 101401 66107 101459 66113
rect 101677 66113 101689 66116
rect 101723 66113 101735 66147
rect 101677 66107 101735 66113
rect 101861 66147 101919 66153
rect 101861 66113 101873 66147
rect 101907 66144 101919 66147
rect 101950 66144 101956 66156
rect 101907 66116 101956 66144
rect 101907 66113 101919 66116
rect 101861 66107 101919 66113
rect 101950 66104 101956 66116
rect 102008 66104 102014 66156
rect 102428 66153 102456 66184
rect 102778 66172 102784 66184
rect 102836 66172 102842 66224
rect 102229 66147 102287 66153
rect 102229 66144 102241 66147
rect 102060 66116 102241 66144
rect 102060 66085 102088 66116
rect 102229 66113 102241 66116
rect 102275 66113 102287 66147
rect 102229 66107 102287 66113
rect 102413 66147 102471 66153
rect 102413 66113 102425 66147
rect 102459 66113 102471 66147
rect 102413 66107 102471 66113
rect 102597 66147 102655 66153
rect 102597 66113 102609 66147
rect 102643 66144 102655 66147
rect 102870 66144 102876 66156
rect 102643 66116 102876 66144
rect 102643 66113 102655 66116
rect 102597 66107 102655 66113
rect 102870 66104 102876 66116
rect 102928 66104 102934 66156
rect 103698 66104 103704 66156
rect 103756 66144 103762 66156
rect 103885 66147 103943 66153
rect 103885 66144 103897 66147
rect 103756 66116 103897 66144
rect 103756 66104 103762 66116
rect 103885 66113 103897 66116
rect 103931 66113 103943 66147
rect 103885 66107 103943 66113
rect 104069 66147 104127 66153
rect 104069 66113 104081 66147
rect 104115 66144 104127 66147
rect 104618 66144 104624 66156
rect 104115 66116 104624 66144
rect 104115 66113 104127 66116
rect 104069 66107 104127 66113
rect 104618 66104 104624 66116
rect 104676 66104 104682 66156
rect 102045 66079 102103 66085
rect 102045 66076 102057 66079
rect 101232 66048 102057 66076
rect 102045 66045 102057 66048
rect 102091 66045 102103 66079
rect 102045 66039 102103 66045
rect 102137 66079 102195 66085
rect 102137 66045 102149 66079
rect 102183 66076 102195 66079
rect 103514 66076 103520 66088
rect 102183 66048 103520 66076
rect 102183 66045 102195 66048
rect 102137 66039 102195 66045
rect 103514 66036 103520 66048
rect 103572 66036 103578 66088
rect 96890 65968 96896 66020
rect 96948 65968 96954 66020
rect 98733 66011 98791 66017
rect 98733 65977 98745 66011
rect 98779 66008 98791 66011
rect 99374 66008 99380 66020
rect 98779 65980 99380 66008
rect 98779 65977 98791 65980
rect 98733 65971 98791 65977
rect 99374 65968 99380 65980
rect 99432 65968 99438 66020
rect 99653 66011 99711 66017
rect 99653 65977 99665 66011
rect 99699 66008 99711 66011
rect 99742 66008 99748 66020
rect 99699 65980 99748 66008
rect 99699 65977 99711 65980
rect 99653 65971 99711 65977
rect 99742 65968 99748 65980
rect 99800 65968 99806 66020
rect 103698 66008 103704 66020
rect 100496 65980 103704 66008
rect 100496 65940 100524 65980
rect 103698 65968 103704 65980
rect 103756 65968 103762 66020
rect 96203 65912 100524 65940
rect 96203 65909 96215 65912
rect 96157 65903 96215 65909
rect 100570 65900 100576 65952
rect 100628 65940 100634 65952
rect 100665 65943 100723 65949
rect 100665 65940 100677 65943
rect 100628 65912 100677 65940
rect 100628 65900 100634 65912
rect 100665 65909 100677 65912
rect 100711 65909 100723 65943
rect 100665 65903 100723 65909
rect 1104 65850 108836 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 96374 65850
rect 96426 65798 96438 65850
rect 96490 65798 96502 65850
rect 96554 65798 96566 65850
rect 96618 65798 96630 65850
rect 96682 65798 105922 65850
rect 105974 65798 105986 65850
rect 106038 65798 106050 65850
rect 106102 65798 106114 65850
rect 106166 65798 106178 65850
rect 106230 65798 108836 65850
rect 1104 65776 108836 65798
rect 94130 65696 94136 65748
rect 94188 65736 94194 65748
rect 103606 65736 103612 65748
rect 94188 65708 103612 65736
rect 94188 65696 94194 65708
rect 103606 65696 103612 65708
rect 103664 65696 103670 65748
rect 94866 65628 94872 65680
rect 94924 65668 94930 65680
rect 102226 65668 102232 65680
rect 94924 65640 102232 65668
rect 94924 65628 94930 65640
rect 102226 65628 102232 65640
rect 102284 65628 102290 65680
rect 1104 65306 7912 65328
rect 1104 65254 4874 65306
rect 4926 65254 4938 65306
rect 4990 65254 5002 65306
rect 5054 65254 5066 65306
rect 5118 65254 5130 65306
rect 5182 65254 7912 65306
rect 1104 65232 7912 65254
rect 104052 65306 108836 65328
rect 104052 65254 106658 65306
rect 106710 65254 106722 65306
rect 106774 65254 106786 65306
rect 106838 65254 106850 65306
rect 106902 65254 106914 65306
rect 106966 65254 108836 65306
rect 104052 65232 108836 65254
rect 1104 64762 7912 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 7912 64762
rect 1104 64688 7912 64710
rect 104052 64762 108836 64784
rect 104052 64710 105922 64762
rect 105974 64710 105986 64762
rect 106038 64710 106050 64762
rect 106102 64710 106114 64762
rect 106166 64710 106178 64762
rect 106230 64710 108836 64762
rect 104052 64688 108836 64710
rect 1104 64218 7912 64240
rect 1104 64166 4874 64218
rect 4926 64166 4938 64218
rect 4990 64166 5002 64218
rect 5054 64166 5066 64218
rect 5118 64166 5130 64218
rect 5182 64166 7912 64218
rect 1104 64144 7912 64166
rect 104052 64218 108836 64240
rect 104052 64166 106658 64218
rect 106710 64166 106722 64218
rect 106774 64166 106786 64218
rect 106838 64166 106850 64218
rect 106902 64166 106914 64218
rect 106966 64166 108836 64218
rect 104052 64144 108836 64166
rect 1104 63674 7912 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 7912 63674
rect 1104 63600 7912 63622
rect 104052 63674 108836 63696
rect 104052 63622 105922 63674
rect 105974 63622 105986 63674
rect 106038 63622 106050 63674
rect 106102 63622 106114 63674
rect 106166 63622 106178 63674
rect 106230 63622 108836 63674
rect 104052 63600 108836 63622
rect 1104 63130 7912 63152
rect 1104 63078 4874 63130
rect 4926 63078 4938 63130
rect 4990 63078 5002 63130
rect 5054 63078 5066 63130
rect 5118 63078 5130 63130
rect 5182 63078 7912 63130
rect 1104 63056 7912 63078
rect 104052 63130 108836 63152
rect 104052 63078 106658 63130
rect 106710 63078 106722 63130
rect 106774 63078 106786 63130
rect 106838 63078 106850 63130
rect 106902 63078 106914 63130
rect 106966 63078 108836 63130
rect 104052 63056 108836 63078
rect 1104 62586 7912 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 7912 62586
rect 1104 62512 7912 62534
rect 104052 62586 108836 62608
rect 104052 62534 105922 62586
rect 105974 62534 105986 62586
rect 106038 62534 106050 62586
rect 106102 62534 106114 62586
rect 106166 62534 106178 62586
rect 106230 62534 108836 62586
rect 104052 62512 108836 62534
rect 1104 62042 7912 62064
rect 1104 61990 4874 62042
rect 4926 61990 4938 62042
rect 4990 61990 5002 62042
rect 5054 61990 5066 62042
rect 5118 61990 5130 62042
rect 5182 61990 7912 62042
rect 1104 61968 7912 61990
rect 104052 62042 108836 62064
rect 104052 61990 106658 62042
rect 106710 61990 106722 62042
rect 106774 61990 106786 62042
rect 106838 61990 106850 62042
rect 106902 61990 106914 62042
rect 106966 61990 108836 62042
rect 104052 61968 108836 61990
rect 1104 61498 7912 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 7912 61498
rect 1104 61424 7912 61446
rect 104052 61498 108836 61520
rect 104052 61446 105922 61498
rect 105974 61446 105986 61498
rect 106038 61446 106050 61498
rect 106102 61446 106114 61498
rect 106166 61446 106178 61498
rect 106230 61446 108836 61498
rect 104052 61424 108836 61446
rect 1104 60954 7912 60976
rect 1104 60902 4874 60954
rect 4926 60902 4938 60954
rect 4990 60902 5002 60954
rect 5054 60902 5066 60954
rect 5118 60902 5130 60954
rect 5182 60902 7912 60954
rect 1104 60880 7912 60902
rect 104052 60954 108836 60976
rect 104052 60902 106658 60954
rect 106710 60902 106722 60954
rect 106774 60902 106786 60954
rect 106838 60902 106850 60954
rect 106902 60902 106914 60954
rect 106966 60902 108836 60954
rect 104052 60880 108836 60902
rect 1104 60410 7912 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 7912 60410
rect 1104 60336 7912 60358
rect 104052 60410 108836 60432
rect 104052 60358 105922 60410
rect 105974 60358 105986 60410
rect 106038 60358 106050 60410
rect 106102 60358 106114 60410
rect 106166 60358 106178 60410
rect 106230 60358 108836 60410
rect 104052 60336 108836 60358
rect 104342 60052 104348 60104
rect 104400 60052 104406 60104
rect 1104 59866 7912 59888
rect 1104 59814 4874 59866
rect 4926 59814 4938 59866
rect 4990 59814 5002 59866
rect 5054 59814 5066 59866
rect 5118 59814 5130 59866
rect 5182 59814 7912 59866
rect 1104 59792 7912 59814
rect 104052 59866 108836 59888
rect 104052 59814 106658 59866
rect 106710 59814 106722 59866
rect 106774 59814 106786 59866
rect 106838 59814 106850 59866
rect 106902 59814 106914 59866
rect 106966 59814 108836 59866
rect 104052 59792 108836 59814
rect 1104 59322 7912 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 7912 59322
rect 1104 59248 7912 59270
rect 104052 59322 108836 59344
rect 104052 59270 105922 59322
rect 105974 59270 105986 59322
rect 106038 59270 106050 59322
rect 106102 59270 106114 59322
rect 106166 59270 106178 59322
rect 106230 59270 108836 59322
rect 104052 59248 108836 59270
rect 1104 58778 7912 58800
rect 1104 58726 4874 58778
rect 4926 58726 4938 58778
rect 4990 58726 5002 58778
rect 5054 58726 5066 58778
rect 5118 58726 5130 58778
rect 5182 58726 7912 58778
rect 1104 58704 7912 58726
rect 104052 58778 108836 58800
rect 104052 58726 106658 58778
rect 106710 58726 106722 58778
rect 106774 58726 106786 58778
rect 106838 58726 106850 58778
rect 106902 58726 106914 58778
rect 106966 58726 108836 58778
rect 104052 58704 108836 58726
rect 1104 58234 7912 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 7912 58234
rect 1104 58160 7912 58182
rect 104052 58234 108836 58256
rect 104052 58182 105922 58234
rect 105974 58182 105986 58234
rect 106038 58182 106050 58234
rect 106102 58182 106114 58234
rect 106166 58182 106178 58234
rect 106230 58182 108836 58234
rect 104052 58160 108836 58182
rect 1104 57690 7912 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 7912 57690
rect 1104 57616 7912 57638
rect 104052 57690 108836 57712
rect 104052 57638 106658 57690
rect 106710 57638 106722 57690
rect 106774 57638 106786 57690
rect 106838 57638 106850 57690
rect 106902 57638 106914 57690
rect 106966 57638 108836 57690
rect 104052 57616 108836 57638
rect 1104 57146 7912 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 7912 57146
rect 1104 57072 7912 57094
rect 104052 57146 108836 57168
rect 104052 57094 105922 57146
rect 105974 57094 105986 57146
rect 106038 57094 106050 57146
rect 106102 57094 106114 57146
rect 106166 57094 106178 57146
rect 106230 57094 108836 57146
rect 104052 57072 108836 57094
rect 1104 56602 7912 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 7912 56602
rect 1104 56528 7912 56550
rect 104052 56602 108836 56624
rect 104052 56550 106658 56602
rect 106710 56550 106722 56602
rect 106774 56550 106786 56602
rect 106838 56550 106850 56602
rect 106902 56550 106914 56602
rect 106966 56550 108836 56602
rect 104052 56528 108836 56550
rect 1104 56058 7912 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 7912 56058
rect 1104 55984 7912 56006
rect 104052 56058 108836 56080
rect 104052 56006 105922 56058
rect 105974 56006 105986 56058
rect 106038 56006 106050 56058
rect 106102 56006 106114 56058
rect 106166 56006 106178 56058
rect 106230 56006 108836 56058
rect 104052 55984 108836 56006
rect 1104 55514 7912 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 7912 55514
rect 1104 55440 7912 55462
rect 104052 55514 108836 55536
rect 104052 55462 106658 55514
rect 106710 55462 106722 55514
rect 106774 55462 106786 55514
rect 106838 55462 106850 55514
rect 106902 55462 106914 55514
rect 106966 55462 108836 55514
rect 104052 55440 108836 55462
rect 1104 54970 7912 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 7912 54970
rect 1104 54896 7912 54918
rect 104052 54970 108836 54992
rect 104052 54918 105922 54970
rect 105974 54918 105986 54970
rect 106038 54918 106050 54970
rect 106102 54918 106114 54970
rect 106166 54918 106178 54970
rect 106230 54918 108836 54970
rect 104052 54896 108836 54918
rect 1104 54426 7912 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 7912 54426
rect 1104 54352 7912 54374
rect 104052 54426 108836 54448
rect 104052 54374 106658 54426
rect 106710 54374 106722 54426
rect 106774 54374 106786 54426
rect 106838 54374 106850 54426
rect 106902 54374 106914 54426
rect 106966 54374 108836 54426
rect 104052 54352 108836 54374
rect 1104 53882 7912 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 7912 53882
rect 1104 53808 7912 53830
rect 104052 53882 108836 53904
rect 104052 53830 105922 53882
rect 105974 53830 105986 53882
rect 106038 53830 106050 53882
rect 106102 53830 106114 53882
rect 106166 53830 106178 53882
rect 106230 53830 108836 53882
rect 104052 53808 108836 53830
rect 1104 53338 7912 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 7912 53338
rect 1104 53264 7912 53286
rect 104052 53338 108836 53360
rect 104052 53286 106658 53338
rect 106710 53286 106722 53338
rect 106774 53286 106786 53338
rect 106838 53286 106850 53338
rect 106902 53286 106914 53338
rect 106966 53286 108836 53338
rect 104052 53264 108836 53286
rect 1104 52794 7912 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 7912 52794
rect 1104 52720 7912 52742
rect 104052 52794 108836 52816
rect 104052 52742 105922 52794
rect 105974 52742 105986 52794
rect 106038 52742 106050 52794
rect 106102 52742 106114 52794
rect 106166 52742 106178 52794
rect 106230 52742 108836 52794
rect 104052 52720 108836 52742
rect 1104 52250 7912 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 7912 52250
rect 1104 52176 7912 52198
rect 104052 52250 108836 52272
rect 104052 52198 106658 52250
rect 106710 52198 106722 52250
rect 106774 52198 106786 52250
rect 106838 52198 106850 52250
rect 106902 52198 106914 52250
rect 106966 52198 108836 52250
rect 104052 52176 108836 52198
rect 1104 51706 7912 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 7912 51706
rect 1104 51632 7912 51654
rect 104052 51706 108836 51728
rect 104052 51654 105922 51706
rect 105974 51654 105986 51706
rect 106038 51654 106050 51706
rect 106102 51654 106114 51706
rect 106166 51654 106178 51706
rect 106230 51654 108836 51706
rect 104052 51632 108836 51654
rect 1104 51162 7912 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 7912 51162
rect 1104 51088 7912 51110
rect 104052 51162 108836 51184
rect 104052 51110 106658 51162
rect 106710 51110 106722 51162
rect 106774 51110 106786 51162
rect 106838 51110 106850 51162
rect 106902 51110 106914 51162
rect 106966 51110 108836 51162
rect 104052 51088 108836 51110
rect 1104 50618 7912 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 7912 50618
rect 1104 50544 7912 50566
rect 104052 50618 108836 50640
rect 104052 50566 105922 50618
rect 105974 50566 105986 50618
rect 106038 50566 106050 50618
rect 106102 50566 106114 50618
rect 106166 50566 106178 50618
rect 106230 50566 108836 50618
rect 104052 50544 108836 50566
rect 1104 50074 7912 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 7912 50074
rect 1104 50000 7912 50022
rect 104052 50074 108836 50096
rect 104052 50022 106658 50074
rect 106710 50022 106722 50074
rect 106774 50022 106786 50074
rect 106838 50022 106850 50074
rect 106902 50022 106914 50074
rect 106966 50022 108836 50074
rect 104052 50000 108836 50022
rect 1104 49530 7912 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 7912 49530
rect 1104 49456 7912 49478
rect 104052 49530 108836 49552
rect 104052 49478 105922 49530
rect 105974 49478 105986 49530
rect 106038 49478 106050 49530
rect 106102 49478 106114 49530
rect 106166 49478 106178 49530
rect 106230 49478 108836 49530
rect 104052 49456 108836 49478
rect 1104 48986 7912 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 7912 48986
rect 1104 48912 7912 48934
rect 104052 48986 108836 49008
rect 104052 48934 106658 48986
rect 106710 48934 106722 48986
rect 106774 48934 106786 48986
rect 106838 48934 106850 48986
rect 106902 48934 106914 48986
rect 106966 48934 108836 48986
rect 104052 48912 108836 48934
rect 1104 48442 7912 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 7912 48442
rect 1104 48368 7912 48390
rect 104052 48442 108836 48464
rect 104052 48390 105922 48442
rect 105974 48390 105986 48442
rect 106038 48390 106050 48442
rect 106102 48390 106114 48442
rect 106166 48390 106178 48442
rect 106230 48390 108836 48442
rect 104052 48368 108836 48390
rect 1104 47898 7912 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 7912 47898
rect 1104 47824 7912 47846
rect 104052 47898 108836 47920
rect 104052 47846 106658 47898
rect 106710 47846 106722 47898
rect 106774 47846 106786 47898
rect 106838 47846 106850 47898
rect 106902 47846 106914 47898
rect 106966 47846 108836 47898
rect 104052 47824 108836 47846
rect 1104 47354 7912 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 7912 47354
rect 1104 47280 7912 47302
rect 104052 47354 108836 47376
rect 104052 47302 105922 47354
rect 105974 47302 105986 47354
rect 106038 47302 106050 47354
rect 106102 47302 106114 47354
rect 106166 47302 106178 47354
rect 106230 47302 108836 47354
rect 104052 47280 108836 47302
rect 1104 46810 7912 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 7912 46810
rect 1104 46736 7912 46758
rect 104052 46810 108836 46832
rect 104052 46758 106658 46810
rect 106710 46758 106722 46810
rect 106774 46758 106786 46810
rect 106838 46758 106850 46810
rect 106902 46758 106914 46810
rect 106966 46758 108836 46810
rect 104052 46736 108836 46758
rect 1104 46266 7912 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 7912 46266
rect 1104 46192 7912 46214
rect 104052 46266 108836 46288
rect 104052 46214 105922 46266
rect 105974 46214 105986 46266
rect 106038 46214 106050 46266
rect 106102 46214 106114 46266
rect 106166 46214 106178 46266
rect 106230 46214 108836 46266
rect 104052 46192 108836 46214
rect 1104 45722 7912 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 7912 45722
rect 1104 45648 7912 45670
rect 104052 45722 108836 45744
rect 104052 45670 106658 45722
rect 106710 45670 106722 45722
rect 106774 45670 106786 45722
rect 106838 45670 106850 45722
rect 106902 45670 106914 45722
rect 106966 45670 108836 45722
rect 104052 45648 108836 45670
rect 1104 45178 7912 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 7912 45178
rect 1104 45104 7912 45126
rect 104052 45178 108836 45200
rect 104052 45126 105922 45178
rect 105974 45126 105986 45178
rect 106038 45126 106050 45178
rect 106102 45126 106114 45178
rect 106166 45126 106178 45178
rect 106230 45126 108836 45178
rect 104052 45104 108836 45126
rect 1104 44634 7912 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 7912 44634
rect 1104 44560 7912 44582
rect 104052 44634 108836 44656
rect 104052 44582 106658 44634
rect 106710 44582 106722 44634
rect 106774 44582 106786 44634
rect 106838 44582 106850 44634
rect 106902 44582 106914 44634
rect 106966 44582 108836 44634
rect 104052 44560 108836 44582
rect 1104 44090 7912 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 7912 44090
rect 1104 44016 7912 44038
rect 104052 44090 108836 44112
rect 104052 44038 105922 44090
rect 105974 44038 105986 44090
rect 106038 44038 106050 44090
rect 106102 44038 106114 44090
rect 106166 44038 106178 44090
rect 106230 44038 108836 44090
rect 104052 44016 108836 44038
rect 1104 43546 7912 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 7912 43546
rect 1104 43472 7912 43494
rect 104052 43546 108836 43568
rect 104052 43494 106658 43546
rect 106710 43494 106722 43546
rect 106774 43494 106786 43546
rect 106838 43494 106850 43546
rect 106902 43494 106914 43546
rect 106966 43494 108836 43546
rect 104052 43472 108836 43494
rect 1104 43002 7912 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 7912 43002
rect 1104 42928 7912 42950
rect 104052 43002 108836 43024
rect 104052 42950 105922 43002
rect 105974 42950 105986 43002
rect 106038 42950 106050 43002
rect 106102 42950 106114 43002
rect 106166 42950 106178 43002
rect 106230 42950 108836 43002
rect 104052 42928 108836 42950
rect 1104 42458 7912 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 7912 42458
rect 1104 42384 7912 42406
rect 104052 42458 108836 42480
rect 104052 42406 106658 42458
rect 106710 42406 106722 42458
rect 106774 42406 106786 42458
rect 106838 42406 106850 42458
rect 106902 42406 106914 42458
rect 106966 42406 108836 42458
rect 104052 42384 108836 42406
rect 1104 41914 7912 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 7912 41914
rect 1104 41840 7912 41862
rect 104052 41914 108836 41936
rect 104052 41862 105922 41914
rect 105974 41862 105986 41914
rect 106038 41862 106050 41914
rect 106102 41862 106114 41914
rect 106166 41862 106178 41914
rect 106230 41862 108836 41914
rect 104052 41840 108836 41862
rect 7558 41420 7564 41472
rect 7616 41420 7622 41472
rect 1104 41370 7912 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 7912 41370
rect 1104 41296 7912 41318
rect 104052 41370 108836 41392
rect 104052 41318 106658 41370
rect 106710 41318 106722 41370
rect 106774 41318 106786 41370
rect 106838 41318 106850 41370
rect 106902 41318 106914 41370
rect 106966 41318 108836 41370
rect 104052 41296 108836 41318
rect 1104 40826 7912 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 7912 40826
rect 1104 40752 7912 40774
rect 104052 40826 108836 40848
rect 104052 40774 105922 40826
rect 105974 40774 105986 40826
rect 106038 40774 106050 40826
rect 106102 40774 106114 40826
rect 106166 40774 106178 40826
rect 106230 40774 108836 40826
rect 104052 40752 108836 40774
rect 1104 40282 7912 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 7912 40282
rect 1104 40208 7912 40230
rect 104052 40282 108836 40304
rect 104052 40230 106658 40282
rect 106710 40230 106722 40282
rect 106774 40230 106786 40282
rect 106838 40230 106850 40282
rect 106902 40230 106914 40282
rect 106966 40230 108836 40282
rect 104052 40208 108836 40230
rect 3418 39992 3424 40044
rect 3476 40032 3482 40044
rect 7558 40032 7564 40044
rect 3476 40004 7564 40032
rect 3476 39992 3482 40004
rect 7558 39992 7564 40004
rect 7616 39992 7622 40044
rect 7282 39788 7288 39840
rect 7340 39828 7346 39840
rect 7469 39831 7527 39837
rect 7469 39828 7481 39831
rect 7340 39800 7481 39828
rect 7340 39788 7346 39800
rect 7469 39797 7481 39800
rect 7515 39797 7527 39831
rect 7469 39791 7527 39797
rect 1104 39738 7912 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 7912 39738
rect 1104 39664 7912 39686
rect 104052 39738 108836 39760
rect 104052 39686 105922 39738
rect 105974 39686 105986 39738
rect 106038 39686 106050 39738
rect 106102 39686 106114 39738
rect 106166 39686 106178 39738
rect 106230 39686 108836 39738
rect 104052 39664 108836 39686
rect 1104 39194 7912 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 7912 39194
rect 1104 39120 7912 39142
rect 104052 39194 108836 39216
rect 104052 39142 106658 39194
rect 106710 39142 106722 39194
rect 106774 39142 106786 39194
rect 106838 39142 106850 39194
rect 106902 39142 106914 39194
rect 106966 39142 108836 39194
rect 104052 39120 108836 39142
rect 7558 38700 7564 38752
rect 7616 38700 7622 38752
rect 1104 38650 7912 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 7912 38650
rect 1104 38576 7912 38598
rect 104052 38650 108836 38672
rect 104052 38598 105922 38650
rect 105974 38598 105986 38650
rect 106038 38598 106050 38650
rect 106102 38598 106114 38650
rect 106166 38598 106178 38650
rect 106230 38598 108836 38650
rect 104052 38576 108836 38598
rect 1104 38106 7912 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 7912 38106
rect 1104 38032 7912 38054
rect 104052 38106 108836 38128
rect 104052 38054 106658 38106
rect 106710 38054 106722 38106
rect 106774 38054 106786 38106
rect 106838 38054 106850 38106
rect 106902 38054 106914 38106
rect 106966 38054 108836 38106
rect 104052 38032 108836 38054
rect 1104 37562 7912 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 7912 37562
rect 1104 37488 7912 37510
rect 104052 37562 108836 37584
rect 104052 37510 105922 37562
rect 105974 37510 105986 37562
rect 106038 37510 106050 37562
rect 106102 37510 106114 37562
rect 106166 37510 106178 37562
rect 106230 37510 108836 37562
rect 104052 37488 108836 37510
rect 1104 37018 7912 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 7912 37018
rect 1104 36944 7912 36966
rect 104052 37018 108836 37040
rect 104052 36966 106658 37018
rect 106710 36966 106722 37018
rect 106774 36966 106786 37018
rect 106838 36966 106850 37018
rect 106902 36966 106914 37018
rect 106966 36966 108836 37018
rect 104052 36944 108836 36966
rect 7558 36592 7564 36644
rect 7616 36592 7622 36644
rect 1104 36474 7912 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 7912 36474
rect 1104 36400 7912 36422
rect 104052 36474 108836 36496
rect 104052 36422 105922 36474
rect 105974 36422 105986 36474
rect 106038 36422 106050 36474
rect 106102 36422 106114 36474
rect 106166 36422 106178 36474
rect 106230 36422 108836 36474
rect 104052 36400 108836 36422
rect 1104 35930 7912 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 7912 35930
rect 1104 35856 7912 35878
rect 104052 35930 108836 35952
rect 104052 35878 106658 35930
rect 106710 35878 106722 35930
rect 106774 35878 106786 35930
rect 106838 35878 106850 35930
rect 106902 35878 106914 35930
rect 106966 35878 108836 35930
rect 104052 35856 108836 35878
rect 7466 35436 7472 35488
rect 7524 35436 7530 35488
rect 1104 35386 7912 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 7912 35386
rect 1104 35312 7912 35334
rect 104052 35386 108836 35408
rect 104052 35334 105922 35386
rect 105974 35334 105986 35386
rect 106038 35334 106050 35386
rect 106102 35334 106114 35386
rect 106166 35334 106178 35386
rect 106230 35334 108836 35386
rect 104052 35312 108836 35334
rect 1104 34842 7912 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 7912 34842
rect 1104 34768 7912 34790
rect 104052 34842 108836 34864
rect 104052 34790 106658 34842
rect 106710 34790 106722 34842
rect 106774 34790 106786 34842
rect 106838 34790 106850 34842
rect 106902 34790 106914 34842
rect 106966 34790 108836 34842
rect 104052 34768 108836 34790
rect 1104 34298 7912 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 7912 34298
rect 1104 34224 7912 34246
rect 104052 34298 108836 34320
rect 104052 34246 105922 34298
rect 105974 34246 105986 34298
rect 106038 34246 106050 34298
rect 106102 34246 106114 34298
rect 106166 34246 106178 34298
rect 106230 34246 108836 34298
rect 104052 34224 108836 34246
rect 7558 33872 7564 33924
rect 7616 33872 7622 33924
rect 1104 33754 7912 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 7912 33754
rect 1104 33680 7912 33702
rect 104052 33754 108836 33776
rect 104052 33702 106658 33754
rect 106710 33702 106722 33754
rect 106774 33702 106786 33754
rect 106838 33702 106850 33754
rect 106902 33702 106914 33754
rect 106966 33702 108836 33754
rect 104052 33680 108836 33702
rect 1104 33210 7912 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 7912 33210
rect 1104 33136 7912 33158
rect 104052 33210 108836 33232
rect 104052 33158 105922 33210
rect 105974 33158 105986 33210
rect 106038 33158 106050 33210
rect 106102 33158 106114 33210
rect 106166 33158 106178 33210
rect 106230 33158 108836 33210
rect 104052 33136 108836 33158
rect 1578 33056 1584 33108
rect 1636 33096 1642 33108
rect 7558 33096 7564 33108
rect 1636 33068 7564 33096
rect 1636 33056 1642 33068
rect 7558 33056 7564 33068
rect 7616 33056 7622 33108
rect 1104 32666 7912 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 7912 32666
rect 1104 32592 7912 32614
rect 104052 32666 108836 32688
rect 104052 32614 106658 32666
rect 106710 32614 106722 32666
rect 106774 32614 106786 32666
rect 106838 32614 106850 32666
rect 106902 32614 106914 32666
rect 106966 32614 108836 32666
rect 104052 32592 108836 32614
rect 1104 32122 7912 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 7912 32122
rect 1104 32048 7912 32070
rect 104052 32122 108836 32144
rect 104052 32070 105922 32122
rect 105974 32070 105986 32122
rect 106038 32070 106050 32122
rect 106102 32070 106114 32122
rect 106166 32070 106178 32122
rect 106230 32070 108836 32122
rect 104052 32048 108836 32070
rect 1104 31578 7912 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 7912 31578
rect 1104 31504 7912 31526
rect 104052 31578 108836 31600
rect 104052 31526 106658 31578
rect 106710 31526 106722 31578
rect 106774 31526 106786 31578
rect 106838 31526 106850 31578
rect 106902 31526 106914 31578
rect 106966 31526 108836 31578
rect 104052 31504 108836 31526
rect 1104 31034 7912 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 7912 31034
rect 1104 30960 7912 30982
rect 104052 31034 108836 31056
rect 104052 30982 105922 31034
rect 105974 30982 105986 31034
rect 106038 30982 106050 31034
rect 106102 30982 106114 31034
rect 106166 30982 106178 31034
rect 106230 30982 108836 31034
rect 104052 30960 108836 30982
rect 1104 30490 7912 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 7912 30490
rect 1104 30416 7912 30438
rect 104052 30490 108836 30512
rect 104052 30438 106658 30490
rect 106710 30438 106722 30490
rect 106774 30438 106786 30490
rect 106838 30438 106850 30490
rect 106902 30438 106914 30490
rect 106966 30438 108836 30490
rect 104052 30416 108836 30438
rect 1762 30268 1768 30320
rect 1820 30308 1826 30320
rect 7466 30308 7472 30320
rect 1820 30280 7472 30308
rect 1820 30268 1826 30280
rect 7466 30268 7472 30280
rect 7524 30268 7530 30320
rect 1104 29946 7912 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 7912 29946
rect 1104 29872 7912 29894
rect 104052 29946 108836 29968
rect 104052 29894 105922 29946
rect 105974 29894 105986 29946
rect 106038 29894 106050 29946
rect 106102 29894 106114 29946
rect 106166 29894 106178 29946
rect 106230 29894 108836 29946
rect 104052 29872 108836 29894
rect 1104 29402 7912 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 7912 29402
rect 1104 29328 7912 29350
rect 104052 29402 108836 29424
rect 104052 29350 106658 29402
rect 106710 29350 106722 29402
rect 106774 29350 106786 29402
rect 106838 29350 106850 29402
rect 106902 29350 106914 29402
rect 106966 29350 108836 29402
rect 104052 29328 108836 29350
rect 1104 28858 7912 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 7912 28858
rect 1104 28784 7912 28806
rect 104052 28858 108836 28880
rect 104052 28806 105922 28858
rect 105974 28806 105986 28858
rect 106038 28806 106050 28858
rect 106102 28806 106114 28858
rect 106166 28806 106178 28858
rect 106230 28806 108836 28858
rect 104052 28784 108836 28806
rect 1104 28314 7912 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 7912 28314
rect 1104 28240 7912 28262
rect 104052 28314 108836 28336
rect 104052 28262 106658 28314
rect 106710 28262 106722 28314
rect 106774 28262 106786 28314
rect 106838 28262 106850 28314
rect 106902 28262 106914 28314
rect 106966 28262 108836 28314
rect 104052 28240 108836 28262
rect 1104 27770 7912 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 7912 27770
rect 1104 27696 7912 27718
rect 104052 27770 108836 27792
rect 104052 27718 105922 27770
rect 105974 27718 105986 27770
rect 106038 27718 106050 27770
rect 106102 27718 106114 27770
rect 106166 27718 106178 27770
rect 106230 27718 108836 27770
rect 104052 27696 108836 27718
rect 1104 27226 7912 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 7912 27226
rect 1104 27152 7912 27174
rect 104052 27226 108836 27248
rect 104052 27174 106658 27226
rect 106710 27174 106722 27226
rect 106774 27174 106786 27226
rect 106838 27174 106850 27226
rect 106902 27174 106914 27226
rect 106966 27174 108836 27226
rect 104052 27152 108836 27174
rect 1104 26682 7912 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 7912 26682
rect 1104 26608 7912 26630
rect 104052 26682 108836 26704
rect 104052 26630 105922 26682
rect 105974 26630 105986 26682
rect 106038 26630 106050 26682
rect 106102 26630 106114 26682
rect 106166 26630 106178 26682
rect 106230 26630 108836 26682
rect 104052 26608 108836 26630
rect 1854 26256 1860 26308
rect 1912 26296 1918 26308
rect 7374 26296 7380 26308
rect 1912 26268 7380 26296
rect 1912 26256 1918 26268
rect 7374 26256 7380 26268
rect 7432 26256 7438 26308
rect 1104 26138 7912 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 7912 26138
rect 1104 26064 7912 26086
rect 104052 26138 108836 26160
rect 104052 26086 106658 26138
rect 106710 26086 106722 26138
rect 106774 26086 106786 26138
rect 106838 26086 106850 26138
rect 106902 26086 106914 26138
rect 106966 26086 108836 26138
rect 104052 26064 108836 26086
rect 1104 25594 7912 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 7912 25594
rect 1104 25520 7912 25542
rect 104052 25594 108836 25616
rect 104052 25542 105922 25594
rect 105974 25542 105986 25594
rect 106038 25542 106050 25594
rect 106102 25542 106114 25594
rect 106166 25542 106178 25594
rect 106230 25542 108836 25594
rect 104052 25520 108836 25542
rect 102594 25100 102600 25152
rect 102652 25140 102658 25152
rect 104345 25143 104403 25149
rect 104345 25140 104357 25143
rect 102652 25112 104357 25140
rect 102652 25100 102658 25112
rect 104345 25109 104357 25112
rect 104391 25109 104403 25143
rect 104345 25103 104403 25109
rect 1104 25050 7912 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 7912 25050
rect 1104 24976 7912 24998
rect 104052 25050 108836 25072
rect 104052 24998 106658 25050
rect 106710 24998 106722 25050
rect 106774 24998 106786 25050
rect 106838 24998 106850 25050
rect 106902 24998 106914 25050
rect 106966 24998 108836 25050
rect 104052 24976 108836 24998
rect 1104 24506 7912 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 7912 24506
rect 1104 24432 7912 24454
rect 104052 24506 108836 24528
rect 104052 24454 105922 24506
rect 105974 24454 105986 24506
rect 106038 24454 106050 24506
rect 106102 24454 106114 24506
rect 106166 24454 106178 24506
rect 106230 24454 108836 24506
rect 104052 24432 108836 24454
rect 2038 24012 2044 24064
rect 2096 24052 2102 24064
rect 7558 24052 7564 24064
rect 2096 24024 7564 24052
rect 2096 24012 2102 24024
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 1104 23962 7912 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 7912 23962
rect 1104 23888 7912 23910
rect 104052 23962 108836 23984
rect 104052 23910 106658 23962
rect 106710 23910 106722 23962
rect 106774 23910 106786 23962
rect 106838 23910 106850 23962
rect 106902 23910 106914 23962
rect 106966 23910 108836 23962
rect 104052 23888 108836 23910
rect 102778 23468 102784 23520
rect 102836 23508 102842 23520
rect 104345 23511 104403 23517
rect 104345 23508 104357 23511
rect 102836 23480 104357 23508
rect 102836 23468 102842 23480
rect 104345 23477 104357 23480
rect 104391 23477 104403 23511
rect 104345 23471 104403 23477
rect 1104 23418 7912 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 7912 23418
rect 1104 23344 7912 23366
rect 104052 23418 108836 23440
rect 104052 23366 105922 23418
rect 105974 23366 105986 23418
rect 106038 23366 106050 23418
rect 106102 23366 106114 23418
rect 106166 23366 106178 23418
rect 106230 23366 108836 23418
rect 104052 23344 108836 23366
rect 1104 22874 7912 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 7912 22874
rect 1104 22800 7912 22822
rect 104052 22874 108836 22896
rect 104052 22822 106658 22874
rect 106710 22822 106722 22874
rect 106774 22822 106786 22874
rect 106838 22822 106850 22874
rect 106902 22822 106914 22874
rect 106966 22822 108836 22874
rect 104052 22800 108836 22822
rect 102134 22720 102140 22772
rect 102192 22760 102198 22772
rect 104345 22763 104403 22769
rect 104345 22760 104357 22763
rect 102192 22732 104357 22760
rect 102192 22720 102198 22732
rect 104345 22729 104357 22732
rect 104391 22729 104403 22763
rect 104345 22723 104403 22729
rect 1104 22330 7912 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 7912 22330
rect 1104 22256 7912 22278
rect 104052 22330 108836 22352
rect 104052 22278 105922 22330
rect 105974 22278 105986 22330
rect 106038 22278 106050 22330
rect 106102 22278 106114 22330
rect 106166 22278 106178 22330
rect 106230 22278 108836 22330
rect 104052 22256 108836 22278
rect 1104 21786 7912 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 7912 21786
rect 1104 21712 7912 21734
rect 104052 21786 108836 21808
rect 104052 21734 106658 21786
rect 106710 21734 106722 21786
rect 106774 21734 106786 21786
rect 106838 21734 106850 21786
rect 106902 21734 106914 21786
rect 106966 21734 108836 21786
rect 104052 21712 108836 21734
rect 1104 21242 7912 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 7912 21242
rect 1104 21168 7912 21190
rect 104052 21242 108836 21264
rect 104052 21190 105922 21242
rect 105974 21190 105986 21242
rect 106038 21190 106050 21242
rect 106102 21190 106114 21242
rect 106166 21190 106178 21242
rect 106230 21190 108836 21242
rect 104052 21168 108836 21190
rect 1104 20698 7912 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 7912 20698
rect 1104 20624 7912 20646
rect 104052 20698 108836 20720
rect 104052 20646 106658 20698
rect 106710 20646 106722 20698
rect 106774 20646 106786 20698
rect 106838 20646 106850 20698
rect 106902 20646 106914 20698
rect 106966 20646 108836 20698
rect 104052 20624 108836 20646
rect 1104 20154 7912 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 7912 20154
rect 1104 20080 7912 20102
rect 104052 20154 108836 20176
rect 104052 20102 105922 20154
rect 105974 20102 105986 20154
rect 106038 20102 106050 20154
rect 106102 20102 106114 20154
rect 106166 20102 106178 20154
rect 106230 20102 108836 20154
rect 104052 20080 108836 20102
rect 1104 19610 7912 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 7912 19610
rect 1104 19536 7912 19558
rect 104052 19610 108836 19632
rect 104052 19558 106658 19610
rect 106710 19558 106722 19610
rect 106774 19558 106786 19610
rect 106838 19558 106850 19610
rect 106902 19558 106914 19610
rect 106966 19558 108836 19610
rect 104052 19536 108836 19558
rect 1104 19066 7912 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 7912 19066
rect 1104 18992 7912 19014
rect 104052 19066 108836 19088
rect 104052 19014 105922 19066
rect 105974 19014 105986 19066
rect 106038 19014 106050 19066
rect 106102 19014 106114 19066
rect 106166 19014 106178 19066
rect 106230 19014 108836 19066
rect 104052 18992 108836 19014
rect 1104 18522 7912 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 7912 18522
rect 1104 18448 7912 18470
rect 104052 18522 108836 18544
rect 104052 18470 106658 18522
rect 106710 18470 106722 18522
rect 106774 18470 106786 18522
rect 106838 18470 106850 18522
rect 106902 18470 106914 18522
rect 106966 18470 108836 18522
rect 104052 18448 108836 18470
rect 1104 17978 7912 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 7912 17978
rect 1104 17904 7912 17926
rect 104052 17978 108836 18000
rect 104052 17926 105922 17978
rect 105974 17926 105986 17978
rect 106038 17926 106050 17978
rect 106102 17926 106114 17978
rect 106166 17926 106178 17978
rect 106230 17926 108836 17978
rect 104052 17904 108836 17926
rect 1104 17434 7912 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 7912 17434
rect 1104 17360 7912 17382
rect 104052 17434 108836 17456
rect 104052 17382 106658 17434
rect 106710 17382 106722 17434
rect 106774 17382 106786 17434
rect 106838 17382 106850 17434
rect 106902 17382 106914 17434
rect 106966 17382 108836 17434
rect 104052 17360 108836 17382
rect 1104 16890 7912 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 7912 16890
rect 1104 16816 7912 16838
rect 104052 16890 108836 16912
rect 104052 16838 105922 16890
rect 105974 16838 105986 16890
rect 106038 16838 106050 16890
rect 106102 16838 106114 16890
rect 106166 16838 106178 16890
rect 106230 16838 108836 16890
rect 104052 16816 108836 16838
rect 1104 16346 7912 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 7912 16346
rect 1104 16272 7912 16294
rect 104052 16346 108836 16368
rect 104052 16294 106658 16346
rect 106710 16294 106722 16346
rect 106774 16294 106786 16346
rect 106838 16294 106850 16346
rect 106902 16294 106914 16346
rect 106966 16294 108836 16346
rect 104052 16272 108836 16294
rect 1104 15802 7912 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 7912 15802
rect 1104 15728 7912 15750
rect 104052 15802 108836 15824
rect 104052 15750 105922 15802
rect 105974 15750 105986 15802
rect 106038 15750 106050 15802
rect 106102 15750 106114 15802
rect 106166 15750 106178 15802
rect 106230 15750 108836 15802
rect 104052 15728 108836 15750
rect 7466 15308 7472 15360
rect 7524 15308 7530 15360
rect 1104 15258 7912 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 7912 15258
rect 1104 15184 7912 15206
rect 104052 15258 108836 15280
rect 104052 15206 106658 15258
rect 106710 15206 106722 15258
rect 106774 15206 106786 15258
rect 106838 15206 106850 15258
rect 106902 15206 106914 15258
rect 106966 15206 108836 15258
rect 104052 15184 108836 15206
rect 1104 14714 7912 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 7912 14714
rect 1104 14640 7912 14662
rect 104052 14714 108836 14736
rect 104052 14662 105922 14714
rect 105974 14662 105986 14714
rect 106038 14662 106050 14714
rect 106102 14662 106114 14714
rect 106166 14662 106178 14714
rect 106230 14662 108836 14714
rect 104052 14640 108836 14662
rect 1104 14170 7912 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 7912 14170
rect 1104 14096 7912 14118
rect 104052 14170 108836 14192
rect 104052 14118 106658 14170
rect 106710 14118 106722 14170
rect 106774 14118 106786 14170
rect 106838 14118 106850 14170
rect 106902 14118 106914 14170
rect 106966 14118 108836 14170
rect 104052 14096 108836 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1627 14028 1869 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1857 14025 1869 14028
rect 1903 14056 1915 14059
rect 3418 14056 3424 14068
rect 1903 14028 3424 14056
rect 1903 14025 1915 14028
rect 1857 14019 1915 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1949 13923 2007 13929
rect 1949 13920 1961 13923
rect 1544 13892 1961 13920
rect 1544 13880 1550 13892
rect 1949 13889 1961 13892
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 1104 13626 7912 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 7912 13626
rect 1104 13552 7912 13574
rect 104052 13626 108836 13648
rect 104052 13574 105922 13626
rect 105974 13574 105986 13626
rect 106038 13574 106050 13626
rect 106102 13574 106114 13626
rect 106166 13574 106178 13626
rect 106230 13574 108836 13626
rect 104052 13552 108836 13574
rect 1581 13515 1639 13521
rect 1581 13481 1593 13515
rect 1627 13512 1639 13515
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1627 13484 1869 13512
rect 1627 13481 1639 13484
rect 1581 13475 1639 13481
rect 1857 13481 1869 13484
rect 1903 13512 1915 13515
rect 2038 13512 2044 13524
rect 1903 13484 2044 13512
rect 1903 13481 1915 13484
rect 1857 13475 1915 13481
rect 2038 13472 2044 13484
rect 2096 13472 2102 13524
rect 1302 13200 1308 13252
rect 1360 13240 1366 13252
rect 1489 13243 1547 13249
rect 1489 13240 1501 13243
rect 1360 13212 1501 13240
rect 1360 13200 1366 13212
rect 1489 13209 1501 13212
rect 1535 13240 1547 13243
rect 1949 13243 2007 13249
rect 1949 13240 1961 13243
rect 1535 13212 1961 13240
rect 1535 13209 1547 13212
rect 1489 13203 1547 13209
rect 1949 13209 1961 13212
rect 1995 13209 2007 13243
rect 1949 13203 2007 13209
rect 1104 13082 7912 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 7912 13082
rect 1104 13008 7912 13030
rect 104052 13082 108836 13104
rect 104052 13030 106658 13082
rect 106710 13030 106722 13082
rect 106774 13030 106786 13082
rect 106838 13030 106850 13082
rect 106902 13030 106914 13082
rect 106966 13030 108836 13082
rect 104052 13008 108836 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 1854 12968 1860 12980
rect 1627 12940 1860 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 1486 12792 1492 12844
rect 1544 12832 1550 12844
rect 1949 12835 2007 12841
rect 1949 12832 1961 12835
rect 1544 12804 1961 12832
rect 1544 12792 1550 12804
rect 1949 12801 1961 12804
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 1104 12538 7912 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 7912 12538
rect 1104 12464 7912 12486
rect 104052 12538 108836 12560
rect 104052 12486 105922 12538
rect 105974 12486 105986 12538
rect 106038 12486 106050 12538
rect 106102 12486 106114 12538
rect 106166 12486 106178 12538
rect 106230 12486 108836 12538
rect 104052 12464 108836 12486
rect 1104 11994 7912 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 7912 11994
rect 1104 11920 7912 11942
rect 104052 11994 108836 12016
rect 104052 11942 106658 11994
rect 106710 11942 106722 11994
rect 106774 11942 106786 11994
rect 106838 11942 106850 11994
rect 106902 11942 106914 11994
rect 106966 11942 108836 11994
rect 104052 11920 108836 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 1762 11880 1768 11892
rect 1627 11852 1768 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 1762 11840 1768 11852
rect 1820 11840 1826 11892
rect 1210 11704 1216 11756
rect 1268 11744 1274 11756
rect 1489 11747 1547 11753
rect 1489 11744 1501 11747
rect 1268 11716 1501 11744
rect 1268 11704 1274 11716
rect 1489 11713 1501 11716
rect 1535 11744 1547 11747
rect 1949 11747 2007 11753
rect 1949 11744 1961 11747
rect 1535 11716 1961 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1949 11713 1961 11716
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 1104 11450 7912 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 7912 11450
rect 1104 11376 7912 11398
rect 104052 11450 108836 11472
rect 104052 11398 105922 11450
rect 105974 11398 105986 11450
rect 106038 11398 106050 11450
rect 106102 11398 106114 11450
rect 106166 11398 106178 11450
rect 106230 11398 108836 11450
rect 104052 11376 108836 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1857 11339 1915 11345
rect 1857 11336 1869 11339
rect 1627 11308 1869 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1857 11305 1869 11308
rect 1903 11336 1915 11339
rect 7282 11336 7288 11348
rect 1903 11308 7288 11336
rect 1903 11305 1915 11308
rect 1857 11299 1915 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 1486 11024 1492 11076
rect 1544 11064 1550 11076
rect 1949 11067 2007 11073
rect 1949 11064 1961 11067
rect 1544 11036 1961 11064
rect 1544 11024 1550 11036
rect 1949 11033 1961 11036
rect 1995 11033 2007 11067
rect 1949 11027 2007 11033
rect 1104 10906 7912 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 7912 10906
rect 1104 10832 7912 10854
rect 104052 10906 108836 10928
rect 104052 10854 106658 10906
rect 106710 10854 106722 10906
rect 106774 10854 106786 10906
rect 106838 10854 106850 10906
rect 106902 10854 106914 10906
rect 106966 10854 108836 10906
rect 104052 10832 108836 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 1765 10795 1823 10801
rect 1765 10792 1777 10795
rect 1636 10764 1777 10792
rect 1636 10752 1642 10764
rect 1765 10761 1777 10764
rect 1811 10761 1823 10795
rect 1765 10755 1823 10761
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 1489 10659 1547 10665
rect 1489 10656 1501 10659
rect 1360 10628 1501 10656
rect 1360 10616 1366 10628
rect 1489 10625 1501 10628
rect 1535 10656 1547 10659
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1535 10628 1961 10656
rect 1535 10625 1547 10628
rect 1489 10619 1547 10625
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 1104 10362 7912 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 7912 10362
rect 1104 10288 7912 10310
rect 104052 10362 108836 10384
rect 104052 10310 105922 10362
rect 105974 10310 105986 10362
rect 106038 10310 106050 10362
rect 106102 10310 106114 10362
rect 106166 10310 106178 10362
rect 106230 10310 108836 10362
rect 104052 10288 108836 10310
rect 1486 9936 1492 9988
rect 1544 9936 1550 9988
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 1857 9979 1915 9985
rect 1857 9976 1869 9979
rect 1719 9948 1869 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 1857 9945 1869 9948
rect 1903 9976 1915 9979
rect 1903 9948 6914 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 1504 9908 1532 9936
rect 1949 9911 2007 9917
rect 1949 9908 1961 9911
rect 1504 9880 1961 9908
rect 1949 9877 1961 9880
rect 1995 9877 2007 9911
rect 6886 9908 6914 9948
rect 29546 9908 29552 9920
rect 6886 9880 29552 9908
rect 1949 9871 2007 9877
rect 29546 9868 29552 9880
rect 29604 9868 29610 9920
rect 1104 9818 7912 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 7912 9818
rect 1104 9744 7912 9766
rect 104052 9818 108836 9840
rect 104052 9766 106658 9818
rect 106710 9766 106722 9818
rect 106774 9766 106786 9818
rect 106838 9766 106850 9818
rect 106902 9766 106914 9818
rect 106966 9766 108836 9818
rect 104052 9744 108836 9766
rect 9490 9596 9496 9648
rect 9548 9636 9554 9648
rect 16022 9636 16028 9648
rect 9548 9608 16028 9636
rect 9548 9596 9554 9608
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 16114 9568 16120 9580
rect 9640 9540 16120 9568
rect 9640 9528 9646 9540
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 1104 9274 7912 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 7912 9274
rect 1104 9200 7912 9222
rect 104052 9274 108836 9296
rect 104052 9222 105922 9274
rect 105974 9222 105986 9274
rect 106038 9222 106050 9274
rect 106102 9222 106114 9274
rect 106166 9222 106178 9274
rect 106230 9222 108836 9274
rect 104052 9200 108836 9222
rect 90818 9052 90824 9104
rect 90876 9092 90882 9104
rect 103974 9092 103980 9104
rect 90876 9064 103980 9092
rect 90876 9052 90882 9064
rect 103974 9052 103980 9064
rect 104032 9052 104038 9104
rect 90634 8984 90640 9036
rect 90692 9024 90698 9036
rect 103698 9024 103704 9036
rect 90692 8996 103704 9024
rect 90692 8984 90698 8996
rect 103698 8984 103704 8996
rect 103756 8984 103762 9036
rect 90542 8916 90548 8968
rect 90600 8956 90606 8968
rect 103606 8956 103612 8968
rect 90600 8928 103612 8956
rect 90600 8916 90606 8928
rect 103606 8916 103612 8928
rect 103664 8916 103670 8968
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 1489 8891 1547 8897
rect 1489 8888 1501 8891
rect 1268 8860 1501 8888
rect 1268 8848 1274 8860
rect 1489 8857 1501 8860
rect 1535 8857 1547 8891
rect 1489 8851 1547 8857
rect 1673 8891 1731 8897
rect 1673 8857 1685 8891
rect 1719 8888 1731 8891
rect 1857 8891 1915 8897
rect 1857 8888 1869 8891
rect 1719 8860 1869 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 1857 8857 1869 8860
rect 1903 8888 1915 8891
rect 1903 8860 6914 8888
rect 1903 8857 1915 8860
rect 1857 8851 1915 8857
rect 1504 8820 1532 8851
rect 1949 8823 2007 8829
rect 1949 8820 1961 8823
rect 1504 8792 1961 8820
rect 1949 8789 1961 8792
rect 1995 8789 2007 8823
rect 6886 8820 6914 8860
rect 26694 8820 26700 8832
rect 6886 8792 26700 8820
rect 1949 8783 2007 8789
rect 26694 8780 26700 8792
rect 26752 8780 26758 8832
rect 1104 8730 7912 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 7912 8730
rect 1104 8656 7912 8678
rect 104052 8730 108836 8752
rect 104052 8678 106658 8730
rect 106710 8678 106722 8730
rect 106774 8678 106786 8730
rect 106838 8678 106850 8730
rect 106902 8678 106914 8730
rect 106966 8678 108836 8730
rect 104052 8656 108836 8678
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8381 2007 8415
rect 1949 8375 2007 8381
rect 1964 8344 1992 8375
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 2096 8384 2237 8412
rect 2096 8372 2102 8384
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 2409 8347 2467 8353
rect 2409 8344 2421 8347
rect 1964 8316 2421 8344
rect 2409 8313 2421 8316
rect 2455 8344 2467 8347
rect 24670 8344 24676 8356
rect 2455 8316 24676 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 24670 8304 24676 8316
rect 24728 8304 24734 8356
rect 1104 8186 7912 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 7912 8186
rect 1104 8112 7912 8134
rect 104052 8186 108836 8208
rect 104052 8134 105922 8186
rect 105974 8134 105986 8186
rect 106038 8134 106050 8186
rect 106102 8134 106114 8186
rect 106166 8134 106178 8186
rect 106230 8134 108836 8186
rect 104052 8112 108836 8134
rect 1946 8032 1952 8084
rect 2004 8032 2010 8084
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 1504 7840 2145 7868
rect 1302 7760 1308 7812
rect 1360 7800 1366 7812
rect 1504 7809 1532 7840
rect 2133 7837 2145 7840
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 1489 7803 1547 7809
rect 1489 7800 1501 7803
rect 1360 7772 1501 7800
rect 1360 7760 1366 7772
rect 1489 7769 1501 7772
rect 1535 7769 1547 7803
rect 1489 7763 1547 7769
rect 1673 7803 1731 7809
rect 1673 7769 1685 7803
rect 1719 7800 1731 7803
rect 1857 7803 1915 7809
rect 1857 7800 1869 7803
rect 1719 7772 1869 7800
rect 1719 7769 1731 7772
rect 1673 7763 1731 7769
rect 1857 7769 1869 7772
rect 1903 7800 1915 7803
rect 1903 7772 6914 7800
rect 1903 7769 1915 7772
rect 1857 7763 1915 7769
rect 6886 7732 6914 7772
rect 30466 7732 30472 7744
rect 6886 7704 30472 7732
rect 30466 7692 30472 7704
rect 30524 7692 30530 7744
rect 1104 7642 108836 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 66314 7642
rect 66366 7590 66378 7642
rect 66430 7590 66442 7642
rect 66494 7590 66506 7642
rect 66558 7590 66570 7642
rect 66622 7590 97034 7642
rect 97086 7590 97098 7642
rect 97150 7590 97162 7642
rect 97214 7590 97226 7642
rect 97278 7590 97290 7642
rect 97342 7590 106658 7642
rect 106710 7590 106722 7642
rect 106774 7590 106786 7642
rect 106838 7590 106850 7642
rect 106902 7590 106914 7642
rect 106966 7590 108836 7642
rect 1104 7568 108836 7590
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 16080 7500 16129 7528
rect 16080 7488 16086 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16117 7491 16175 7497
rect 23474 7488 23480 7540
rect 23532 7488 23538 7540
rect 24670 7488 24676 7540
rect 24728 7488 24734 7540
rect 25774 7488 25780 7540
rect 25832 7528 25838 7540
rect 25869 7531 25927 7537
rect 25869 7528 25881 7531
rect 25832 7500 25881 7528
rect 25832 7488 25838 7500
rect 25869 7497 25881 7500
rect 25915 7497 25927 7531
rect 25869 7491 25927 7497
rect 26694 7488 26700 7540
rect 26752 7528 26758 7540
rect 26973 7531 27031 7537
rect 26973 7528 26985 7531
rect 26752 7500 26985 7528
rect 26752 7488 26758 7500
rect 26973 7497 26985 7500
rect 27019 7497 27031 7531
rect 26973 7491 27031 7497
rect 28166 7488 28172 7540
rect 28224 7488 28230 7540
rect 29546 7488 29552 7540
rect 29604 7488 29610 7540
rect 30466 7488 30472 7540
rect 30524 7488 30530 7540
rect 90542 7488 90548 7540
rect 90600 7488 90606 7540
rect 90634 7488 90640 7540
rect 90692 7528 90698 7540
rect 90729 7531 90787 7537
rect 90729 7528 90741 7531
rect 90692 7500 90741 7528
rect 90692 7488 90698 7500
rect 90729 7497 90741 7500
rect 90775 7497 90787 7531
rect 90729 7491 90787 7497
rect 90818 7488 90824 7540
rect 90876 7528 90882 7540
rect 90913 7531 90971 7537
rect 90913 7528 90925 7531
rect 90876 7500 90925 7528
rect 90876 7488 90882 7500
rect 90913 7497 90925 7500
rect 90959 7497 90971 7531
rect 90913 7491 90971 7497
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1489 7395 1547 7401
rect 1489 7392 1501 7395
rect 1360 7364 1501 7392
rect 1360 7352 1366 7364
rect 1489 7361 1501 7364
rect 1535 7392 1547 7395
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1535 7364 1961 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 1857 7259 1915 7265
rect 1857 7256 1869 7259
rect 1719 7228 1869 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 1857 7225 1869 7228
rect 1903 7256 1915 7259
rect 28166 7256 28172 7268
rect 1903 7228 28172 7256
rect 1903 7225 1915 7228
rect 1857 7219 1915 7225
rect 28166 7216 28172 7228
rect 28224 7216 28230 7268
rect 1104 7098 108836 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 105922 7098
rect 105974 7046 105986 7098
rect 106038 7046 106050 7098
rect 106102 7046 106114 7098
rect 106166 7046 106178 7098
rect 106230 7046 108836 7098
rect 1104 7024 108836 7046
rect 1104 6554 108836 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 66314 6554
rect 66366 6502 66378 6554
rect 66430 6502 66442 6554
rect 66494 6502 66506 6554
rect 66558 6502 66570 6554
rect 66622 6502 97034 6554
rect 97086 6502 97098 6554
rect 97150 6502 97162 6554
rect 97214 6502 97226 6554
rect 97278 6502 97290 6554
rect 97342 6502 108836 6554
rect 1104 6480 108836 6502
rect 1210 6264 1216 6316
rect 1268 6304 1274 6316
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 1268 6276 1501 6304
rect 1268 6264 1274 6276
rect 1489 6273 1501 6276
rect 1535 6304 1547 6307
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1535 6276 1961 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1673 6171 1731 6177
rect 1673 6137 1685 6171
rect 1719 6168 1731 6171
rect 1857 6171 1915 6177
rect 1857 6168 1869 6171
rect 1719 6140 1869 6168
rect 1719 6137 1731 6140
rect 1673 6131 1731 6137
rect 1857 6137 1869 6140
rect 1903 6168 1915 6171
rect 1903 6140 6914 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 6886 6100 6914 6140
rect 25866 6100 25872 6112
rect 6886 6072 25872 6100
rect 25866 6060 25872 6072
rect 25924 6060 25930 6112
rect 1104 6010 108836 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 108836 6010
rect 1104 5936 108836 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1765 5899 1823 5905
rect 1765 5896 1777 5899
rect 1627 5868 1777 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1765 5865 1777 5868
rect 1811 5896 1823 5899
rect 7466 5896 7472 5908
rect 1811 5868 7472 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1452 5664 1869 5692
rect 1452 5652 1458 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1104 5466 108836 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 66314 5466
rect 66366 5414 66378 5466
rect 66430 5414 66442 5466
rect 66494 5414 66506 5466
rect 66558 5414 66570 5466
rect 66622 5414 97034 5466
rect 97086 5414 97098 5466
rect 97150 5414 97162 5466
rect 97214 5414 97226 5466
rect 97278 5414 97290 5466
rect 97342 5414 108836 5466
rect 1104 5392 108836 5414
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 1360 5188 1501 5216
rect 1360 5176 1366 5188
rect 1489 5185 1501 5188
rect 1535 5216 1547 5219
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1535 5188 1961 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 1857 5083 1915 5089
rect 1857 5080 1869 5083
rect 1719 5052 1869 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 1857 5049 1869 5052
rect 1903 5080 1915 5083
rect 1903 5052 6914 5080
rect 1903 5049 1915 5052
rect 1857 5043 1915 5049
rect 6886 5012 6914 5052
rect 23474 5012 23480 5024
rect 6886 4984 23480 5012
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 1104 4922 108836 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 108836 4922
rect 1104 4848 108836 4870
rect 1104 4378 108836 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 66314 4378
rect 66366 4326 66378 4378
rect 66430 4326 66442 4378
rect 66494 4326 66506 4378
rect 66558 4326 66570 4378
rect 66622 4326 97034 4378
rect 97086 4326 97098 4378
rect 97150 4326 97162 4378
rect 97214 4326 97226 4378
rect 97278 4326 97290 4378
rect 97342 4326 108836 4378
rect 1104 4304 108836 4326
rect 1104 3834 108836 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 108836 3834
rect 1104 3760 108836 3782
rect 1104 3290 108836 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 66314 3290
rect 66366 3238 66378 3290
rect 66430 3238 66442 3290
rect 66494 3238 66506 3290
rect 66558 3238 66570 3290
rect 66622 3238 97034 3290
rect 97086 3238 97098 3290
rect 97150 3238 97162 3290
rect 97214 3238 97226 3290
rect 97278 3238 97290 3290
rect 97342 3238 108836 3290
rect 1104 3216 108836 3238
rect 1104 2746 108836 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 108836 2746
rect 1104 2672 108836 2694
rect 31662 2592 31668 2644
rect 31720 2592 31726 2644
rect 32950 2592 32956 2644
rect 33008 2592 33014 2644
rect 34238 2592 34244 2644
rect 34296 2592 34302 2644
rect 35434 2592 35440 2644
rect 35492 2632 35498 2644
rect 35529 2635 35587 2641
rect 35529 2632 35541 2635
rect 35492 2604 35541 2632
rect 35492 2592 35498 2604
rect 35529 2601 35541 2604
rect 35575 2601 35587 2635
rect 35529 2595 35587 2601
rect 36354 2592 36360 2644
rect 36412 2592 36418 2644
rect 37458 2592 37464 2644
rect 37516 2592 37522 2644
rect 38746 2592 38752 2644
rect 38804 2592 38810 2644
rect 39942 2592 39948 2644
rect 40000 2632 40006 2644
rect 40037 2635 40095 2641
rect 40037 2632 40049 2635
rect 40000 2604 40049 2632
rect 40000 2592 40006 2604
rect 40037 2601 40049 2604
rect 40083 2601 40095 2635
rect 40037 2595 40095 2601
rect 41322 2592 41328 2644
rect 41380 2592 41386 2644
rect 42150 2592 42156 2644
rect 42208 2592 42214 2644
rect 43438 2592 43444 2644
rect 43496 2592 43502 2644
rect 31849 2431 31907 2437
rect 31849 2428 31861 2431
rect 31588 2400 31861 2428
rect 31588 2304 31616 2400
rect 31849 2397 31861 2400
rect 31895 2397 31907 2431
rect 33137 2431 33195 2437
rect 33137 2428 33149 2431
rect 31849 2391 31907 2397
rect 32876 2400 33149 2428
rect 32876 2304 32904 2400
rect 33137 2397 33149 2400
rect 33183 2397 33195 2431
rect 34425 2431 34483 2437
rect 34425 2428 34437 2431
rect 33137 2391 33195 2397
rect 34164 2400 34437 2428
rect 34164 2304 34192 2400
rect 34425 2397 34437 2400
rect 34471 2397 34483 2431
rect 35713 2431 35771 2437
rect 35713 2428 35725 2431
rect 34425 2391 34483 2397
rect 35452 2400 35725 2428
rect 35452 2304 35480 2400
rect 35713 2397 35725 2400
rect 35759 2397 35771 2431
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35713 2391 35771 2397
rect 36096 2400 36185 2428
rect 36096 2304 36124 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 37645 2431 37703 2437
rect 37645 2428 37657 2431
rect 36173 2391 36231 2397
rect 37384 2400 37657 2428
rect 37384 2304 37412 2400
rect 37645 2397 37657 2400
rect 37691 2397 37703 2431
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 37645 2391 37703 2397
rect 38672 2400 38945 2428
rect 38672 2304 38700 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 38933 2391 38991 2397
rect 39960 2400 40233 2428
rect 39960 2304 39988 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 41509 2431 41567 2437
rect 41509 2428 41521 2431
rect 40221 2391 40279 2397
rect 41248 2400 41521 2428
rect 41248 2304 41276 2400
rect 41509 2397 41521 2400
rect 41555 2397 41567 2431
rect 41969 2431 42027 2437
rect 41969 2428 41981 2431
rect 41509 2391 41567 2397
rect 41892 2400 41981 2428
rect 41892 2304 41920 2400
rect 41969 2397 41981 2400
rect 42015 2397 42027 2431
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 41969 2391 42027 2397
rect 43180 2400 43269 2428
rect 43180 2304 43208 2400
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 43257 2391 43315 2397
rect 31570 2252 31576 2304
rect 31628 2252 31634 2304
rect 32858 2252 32864 2304
rect 32916 2252 32922 2304
rect 34146 2252 34152 2304
rect 34204 2252 34210 2304
rect 35434 2252 35440 2304
rect 35492 2252 35498 2304
rect 36078 2252 36084 2304
rect 36136 2252 36142 2304
rect 37366 2252 37372 2304
rect 37424 2252 37430 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 39942 2252 39948 2304
rect 40000 2252 40006 2304
rect 41230 2252 41236 2304
rect 41288 2252 41294 2304
rect 41874 2252 41880 2304
rect 41932 2252 41938 2304
rect 43162 2252 43168 2304
rect 43220 2252 43226 2304
rect 1104 2202 108836 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 66314 2202
rect 66366 2150 66378 2202
rect 66430 2150 66442 2202
rect 66494 2150 66506 2202
rect 66558 2150 66570 2202
rect 66622 2150 97034 2202
rect 97086 2150 97098 2202
rect 97150 2150 97162 2202
rect 97214 2150 97226 2202
rect 97278 2150 97290 2202
rect 97342 2150 108836 2202
rect 1104 2128 108836 2150
<< via1 >>
rect 4214 147398 4266 147450
rect 4278 147398 4330 147450
rect 4342 147398 4394 147450
rect 4406 147398 4458 147450
rect 4470 147398 4522 147450
rect 34934 147398 34986 147450
rect 34998 147398 35050 147450
rect 35062 147398 35114 147450
rect 35126 147398 35178 147450
rect 35190 147398 35242 147450
rect 65654 147398 65706 147450
rect 65718 147398 65770 147450
rect 65782 147398 65834 147450
rect 65846 147398 65898 147450
rect 65910 147398 65962 147450
rect 96374 147398 96426 147450
rect 96438 147398 96490 147450
rect 96502 147398 96554 147450
rect 96566 147398 96618 147450
rect 96630 147398 96682 147450
rect 4874 146854 4926 146906
rect 4938 146854 4990 146906
rect 5002 146854 5054 146906
rect 5066 146854 5118 146906
rect 5130 146854 5182 146906
rect 35594 146854 35646 146906
rect 35658 146854 35710 146906
rect 35722 146854 35774 146906
rect 35786 146854 35838 146906
rect 35850 146854 35902 146906
rect 66314 146854 66366 146906
rect 66378 146854 66430 146906
rect 66442 146854 66494 146906
rect 66506 146854 66558 146906
rect 66570 146854 66622 146906
rect 97034 146854 97086 146906
rect 97098 146854 97150 146906
rect 97162 146854 97214 146906
rect 97226 146854 97278 146906
rect 97290 146854 97342 146906
rect 4214 146310 4266 146362
rect 4278 146310 4330 146362
rect 4342 146310 4394 146362
rect 4406 146310 4458 146362
rect 4470 146310 4522 146362
rect 34934 146310 34986 146362
rect 34998 146310 35050 146362
rect 35062 146310 35114 146362
rect 35126 146310 35178 146362
rect 35190 146310 35242 146362
rect 65654 146310 65706 146362
rect 65718 146310 65770 146362
rect 65782 146310 65834 146362
rect 65846 146310 65898 146362
rect 65910 146310 65962 146362
rect 96374 146310 96426 146362
rect 96438 146310 96490 146362
rect 96502 146310 96554 146362
rect 96566 146310 96618 146362
rect 96630 146310 96682 146362
rect 4874 145766 4926 145818
rect 4938 145766 4990 145818
rect 5002 145766 5054 145818
rect 5066 145766 5118 145818
rect 5130 145766 5182 145818
rect 35594 145766 35646 145818
rect 35658 145766 35710 145818
rect 35722 145766 35774 145818
rect 35786 145766 35838 145818
rect 35850 145766 35902 145818
rect 66314 145766 66366 145818
rect 66378 145766 66430 145818
rect 66442 145766 66494 145818
rect 66506 145766 66558 145818
rect 66570 145766 66622 145818
rect 97034 145766 97086 145818
rect 97098 145766 97150 145818
rect 97162 145766 97214 145818
rect 97226 145766 97278 145818
rect 97290 145766 97342 145818
rect 4214 145222 4266 145274
rect 4278 145222 4330 145274
rect 4342 145222 4394 145274
rect 4406 145222 4458 145274
rect 4470 145222 4522 145274
rect 34934 145222 34986 145274
rect 34998 145222 35050 145274
rect 35062 145222 35114 145274
rect 35126 145222 35178 145274
rect 35190 145222 35242 145274
rect 65654 145222 65706 145274
rect 65718 145222 65770 145274
rect 65782 145222 65834 145274
rect 65846 145222 65898 145274
rect 65910 145222 65962 145274
rect 96374 145222 96426 145274
rect 96438 145222 96490 145274
rect 96502 145222 96554 145274
rect 96566 145222 96618 145274
rect 96630 145222 96682 145274
rect 4874 144678 4926 144730
rect 4938 144678 4990 144730
rect 5002 144678 5054 144730
rect 5066 144678 5118 144730
rect 5130 144678 5182 144730
rect 35594 144678 35646 144730
rect 35658 144678 35710 144730
rect 35722 144678 35774 144730
rect 35786 144678 35838 144730
rect 35850 144678 35902 144730
rect 66314 144678 66366 144730
rect 66378 144678 66430 144730
rect 66442 144678 66494 144730
rect 66506 144678 66558 144730
rect 66570 144678 66622 144730
rect 97034 144678 97086 144730
rect 97098 144678 97150 144730
rect 97162 144678 97214 144730
rect 97226 144678 97278 144730
rect 97290 144678 97342 144730
rect 4214 144134 4266 144186
rect 4278 144134 4330 144186
rect 4342 144134 4394 144186
rect 4406 144134 4458 144186
rect 4470 144134 4522 144186
rect 34934 144134 34986 144186
rect 34998 144134 35050 144186
rect 35062 144134 35114 144186
rect 35126 144134 35178 144186
rect 35190 144134 35242 144186
rect 65654 144134 65706 144186
rect 65718 144134 65770 144186
rect 65782 144134 65834 144186
rect 65846 144134 65898 144186
rect 65910 144134 65962 144186
rect 96374 144134 96426 144186
rect 96438 144134 96490 144186
rect 96502 144134 96554 144186
rect 96566 144134 96618 144186
rect 96630 144134 96682 144186
rect 4874 143590 4926 143642
rect 4938 143590 4990 143642
rect 5002 143590 5054 143642
rect 5066 143590 5118 143642
rect 5130 143590 5182 143642
rect 35594 143590 35646 143642
rect 35658 143590 35710 143642
rect 35722 143590 35774 143642
rect 35786 143590 35838 143642
rect 35850 143590 35902 143642
rect 66314 143590 66366 143642
rect 66378 143590 66430 143642
rect 66442 143590 66494 143642
rect 66506 143590 66558 143642
rect 66570 143590 66622 143642
rect 97034 143590 97086 143642
rect 97098 143590 97150 143642
rect 97162 143590 97214 143642
rect 97226 143590 97278 143642
rect 97290 143590 97342 143642
rect 4214 143046 4266 143098
rect 4278 143046 4330 143098
rect 4342 143046 4394 143098
rect 4406 143046 4458 143098
rect 4470 143046 4522 143098
rect 34934 143046 34986 143098
rect 34998 143046 35050 143098
rect 35062 143046 35114 143098
rect 35126 143046 35178 143098
rect 35190 143046 35242 143098
rect 65654 143046 65706 143098
rect 65718 143046 65770 143098
rect 65782 143046 65834 143098
rect 65846 143046 65898 143098
rect 65910 143046 65962 143098
rect 96374 143046 96426 143098
rect 96438 143046 96490 143098
rect 96502 143046 96554 143098
rect 96566 143046 96618 143098
rect 96630 143046 96682 143098
rect 4874 142502 4926 142554
rect 4938 142502 4990 142554
rect 5002 142502 5054 142554
rect 5066 142502 5118 142554
rect 5130 142502 5182 142554
rect 35594 142502 35646 142554
rect 35658 142502 35710 142554
rect 35722 142502 35774 142554
rect 35786 142502 35838 142554
rect 35850 142502 35902 142554
rect 66314 142502 66366 142554
rect 66378 142502 66430 142554
rect 66442 142502 66494 142554
rect 66506 142502 66558 142554
rect 66570 142502 66622 142554
rect 97034 142502 97086 142554
rect 97098 142502 97150 142554
rect 97162 142502 97214 142554
rect 97226 142502 97278 142554
rect 97290 142502 97342 142554
rect 4214 141958 4266 142010
rect 4278 141958 4330 142010
rect 4342 141958 4394 142010
rect 4406 141958 4458 142010
rect 4470 141958 4522 142010
rect 34934 141958 34986 142010
rect 34998 141958 35050 142010
rect 35062 141958 35114 142010
rect 35126 141958 35178 142010
rect 35190 141958 35242 142010
rect 65654 141958 65706 142010
rect 65718 141958 65770 142010
rect 65782 141958 65834 142010
rect 65846 141958 65898 142010
rect 65910 141958 65962 142010
rect 96374 141958 96426 142010
rect 96438 141958 96490 142010
rect 96502 141958 96554 142010
rect 96566 141958 96618 142010
rect 96630 141958 96682 142010
rect 4874 141414 4926 141466
rect 4938 141414 4990 141466
rect 5002 141414 5054 141466
rect 5066 141414 5118 141466
rect 5130 141414 5182 141466
rect 35594 141414 35646 141466
rect 35658 141414 35710 141466
rect 35722 141414 35774 141466
rect 35786 141414 35838 141466
rect 35850 141414 35902 141466
rect 66314 141414 66366 141466
rect 66378 141414 66430 141466
rect 66442 141414 66494 141466
rect 66506 141414 66558 141466
rect 66570 141414 66622 141466
rect 97034 141414 97086 141466
rect 97098 141414 97150 141466
rect 97162 141414 97214 141466
rect 97226 141414 97278 141466
rect 97290 141414 97342 141466
rect 4214 140870 4266 140922
rect 4278 140870 4330 140922
rect 4342 140870 4394 140922
rect 4406 140870 4458 140922
rect 4470 140870 4522 140922
rect 34934 140870 34986 140922
rect 34998 140870 35050 140922
rect 35062 140870 35114 140922
rect 35126 140870 35178 140922
rect 35190 140870 35242 140922
rect 65654 140870 65706 140922
rect 65718 140870 65770 140922
rect 65782 140870 65834 140922
rect 65846 140870 65898 140922
rect 65910 140870 65962 140922
rect 96374 140870 96426 140922
rect 96438 140870 96490 140922
rect 96502 140870 96554 140922
rect 96566 140870 96618 140922
rect 96630 140870 96682 140922
rect 4874 140326 4926 140378
rect 4938 140326 4990 140378
rect 5002 140326 5054 140378
rect 5066 140326 5118 140378
rect 5130 140326 5182 140378
rect 35594 140326 35646 140378
rect 35658 140326 35710 140378
rect 35722 140326 35774 140378
rect 35786 140326 35838 140378
rect 35850 140326 35902 140378
rect 66314 140326 66366 140378
rect 66378 140326 66430 140378
rect 66442 140326 66494 140378
rect 66506 140326 66558 140378
rect 66570 140326 66622 140378
rect 97034 140326 97086 140378
rect 97098 140326 97150 140378
rect 97162 140326 97214 140378
rect 97226 140326 97278 140378
rect 97290 140326 97342 140378
rect 4214 139782 4266 139834
rect 4278 139782 4330 139834
rect 4342 139782 4394 139834
rect 4406 139782 4458 139834
rect 4470 139782 4522 139834
rect 34934 139782 34986 139834
rect 34998 139782 35050 139834
rect 35062 139782 35114 139834
rect 35126 139782 35178 139834
rect 35190 139782 35242 139834
rect 65654 139782 65706 139834
rect 65718 139782 65770 139834
rect 65782 139782 65834 139834
rect 65846 139782 65898 139834
rect 65910 139782 65962 139834
rect 96374 139782 96426 139834
rect 96438 139782 96490 139834
rect 96502 139782 96554 139834
rect 96566 139782 96618 139834
rect 96630 139782 96682 139834
rect 4874 139238 4926 139290
rect 4938 139238 4990 139290
rect 5002 139238 5054 139290
rect 5066 139238 5118 139290
rect 5130 139238 5182 139290
rect 35594 139238 35646 139290
rect 35658 139238 35710 139290
rect 35722 139238 35774 139290
rect 35786 139238 35838 139290
rect 35850 139238 35902 139290
rect 66314 139238 66366 139290
rect 66378 139238 66430 139290
rect 66442 139238 66494 139290
rect 66506 139238 66558 139290
rect 66570 139238 66622 139290
rect 97034 139238 97086 139290
rect 97098 139238 97150 139290
rect 97162 139238 97214 139290
rect 97226 139238 97278 139290
rect 97290 139238 97342 139290
rect 4214 138694 4266 138746
rect 4278 138694 4330 138746
rect 4342 138694 4394 138746
rect 4406 138694 4458 138746
rect 4470 138694 4522 138746
rect 34934 138694 34986 138746
rect 34998 138694 35050 138746
rect 35062 138694 35114 138746
rect 35126 138694 35178 138746
rect 35190 138694 35242 138746
rect 65654 138694 65706 138746
rect 65718 138694 65770 138746
rect 65782 138694 65834 138746
rect 65846 138694 65898 138746
rect 65910 138694 65962 138746
rect 96374 138694 96426 138746
rect 96438 138694 96490 138746
rect 96502 138694 96554 138746
rect 96566 138694 96618 138746
rect 96630 138694 96682 138746
rect 4874 138150 4926 138202
rect 4938 138150 4990 138202
rect 5002 138150 5054 138202
rect 5066 138150 5118 138202
rect 5130 138150 5182 138202
rect 35594 138150 35646 138202
rect 35658 138150 35710 138202
rect 35722 138150 35774 138202
rect 35786 138150 35838 138202
rect 35850 138150 35902 138202
rect 66314 138150 66366 138202
rect 66378 138150 66430 138202
rect 66442 138150 66494 138202
rect 66506 138150 66558 138202
rect 66570 138150 66622 138202
rect 97034 138150 97086 138202
rect 97098 138150 97150 138202
rect 97162 138150 97214 138202
rect 97226 138150 97278 138202
rect 97290 138150 97342 138202
rect 4214 137606 4266 137658
rect 4278 137606 4330 137658
rect 4342 137606 4394 137658
rect 4406 137606 4458 137658
rect 4470 137606 4522 137658
rect 34934 137606 34986 137658
rect 34998 137606 35050 137658
rect 35062 137606 35114 137658
rect 35126 137606 35178 137658
rect 35190 137606 35242 137658
rect 65654 137606 65706 137658
rect 65718 137606 65770 137658
rect 65782 137606 65834 137658
rect 65846 137606 65898 137658
rect 65910 137606 65962 137658
rect 96374 137606 96426 137658
rect 96438 137606 96490 137658
rect 96502 137606 96554 137658
rect 96566 137606 96618 137658
rect 96630 137606 96682 137658
rect 4874 137062 4926 137114
rect 4938 137062 4990 137114
rect 5002 137062 5054 137114
rect 5066 137062 5118 137114
rect 5130 137062 5182 137114
rect 35594 137062 35646 137114
rect 35658 137062 35710 137114
rect 35722 137062 35774 137114
rect 35786 137062 35838 137114
rect 35850 137062 35902 137114
rect 66314 137062 66366 137114
rect 66378 137062 66430 137114
rect 66442 137062 66494 137114
rect 66506 137062 66558 137114
rect 66570 137062 66622 137114
rect 97034 137062 97086 137114
rect 97098 137062 97150 137114
rect 97162 137062 97214 137114
rect 97226 137062 97278 137114
rect 97290 137062 97342 137114
rect 63592 136620 63644 136672
rect 102140 136824 102192 136876
rect 95976 136620 96028 136672
rect 4214 136518 4266 136570
rect 4278 136518 4330 136570
rect 4342 136518 4394 136570
rect 4406 136518 4458 136570
rect 4470 136518 4522 136570
rect 34934 136518 34986 136570
rect 34998 136518 35050 136570
rect 35062 136518 35114 136570
rect 35126 136518 35178 136570
rect 35190 136518 35242 136570
rect 65654 136518 65706 136570
rect 65718 136518 65770 136570
rect 65782 136518 65834 136570
rect 65846 136518 65898 136570
rect 65910 136518 65962 136570
rect 96374 136518 96426 136570
rect 96438 136518 96490 136570
rect 96502 136518 96554 136570
rect 96566 136518 96618 136570
rect 96630 136518 96682 136570
rect 105922 136518 105974 136570
rect 105986 136518 106038 136570
rect 106050 136518 106102 136570
rect 106114 136518 106166 136570
rect 106178 136518 106230 136570
rect 35992 136212 36044 136264
rect 34152 136187 34204 136196
rect 34152 136153 34161 136187
rect 34161 136153 34195 136187
rect 34195 136153 34204 136187
rect 34152 136144 34204 136153
rect 34980 136187 35032 136196
rect 34980 136153 34989 136187
rect 34989 136153 35023 136187
rect 35023 136153 35032 136187
rect 34980 136144 35032 136153
rect 38568 136212 38620 136264
rect 38752 136144 38804 136196
rect 43168 136187 43220 136196
rect 43168 136153 43177 136187
rect 43177 136153 43211 136187
rect 43211 136153 43220 136187
rect 43168 136144 43220 136153
rect 48504 136144 48556 136196
rect 51080 136144 51132 136196
rect 55404 136187 55456 136196
rect 55404 136153 55413 136187
rect 55413 136153 55447 136187
rect 55447 136153 55456 136187
rect 55404 136144 55456 136153
rect 57980 136187 58032 136196
rect 57980 136153 57989 136187
rect 57989 136153 58023 136187
rect 58023 136153 58032 136187
rect 57980 136144 58032 136153
rect 60556 136187 60608 136196
rect 60556 136153 60565 136187
rect 60565 136153 60599 136187
rect 60599 136153 60608 136187
rect 60556 136144 60608 136153
rect 36084 136119 36136 136128
rect 36084 136085 36093 136119
rect 36093 136085 36127 136119
rect 36127 136085 36136 136119
rect 36084 136076 36136 136085
rect 43076 136119 43128 136128
rect 43076 136085 43085 136119
rect 43085 136085 43119 136119
rect 43119 136085 43128 136119
rect 43076 136076 43128 136085
rect 46112 136119 46164 136128
rect 46112 136085 46121 136119
rect 46121 136085 46155 136119
rect 46155 136085 46164 136119
rect 46112 136076 46164 136085
rect 47676 136119 47728 136128
rect 47676 136085 47685 136119
rect 47685 136085 47719 136119
rect 47719 136085 47728 136119
rect 47676 136076 47728 136085
rect 50252 136119 50304 136128
rect 50252 136085 50261 136119
rect 50261 136085 50295 136119
rect 50295 136085 50304 136119
rect 50252 136076 50304 136085
rect 55772 136119 55824 136128
rect 55772 136085 55781 136119
rect 55781 136085 55815 136119
rect 55815 136085 55824 136119
rect 55772 136076 55824 136085
rect 58348 136119 58400 136128
rect 58348 136085 58357 136119
rect 58357 136085 58391 136119
rect 58391 136085 58400 136119
rect 58348 136076 58400 136085
rect 63132 136187 63184 136196
rect 63132 136153 63141 136187
rect 63141 136153 63175 136187
rect 63175 136153 63184 136187
rect 63132 136144 63184 136153
rect 72516 136187 72568 136196
rect 72516 136153 72525 136187
rect 72525 136153 72559 136187
rect 72559 136153 72568 136187
rect 72516 136144 72568 136153
rect 72700 136144 72752 136196
rect 77392 136187 77444 136196
rect 77392 136153 77401 136187
rect 77401 136153 77435 136187
rect 77435 136153 77444 136187
rect 77392 136144 77444 136153
rect 60924 136119 60976 136128
rect 60924 136085 60933 136119
rect 60933 136085 60967 136119
rect 60967 136085 60976 136119
rect 60924 136076 60976 136085
rect 63500 136119 63552 136128
rect 63500 136085 63509 136119
rect 63509 136085 63543 136119
rect 63543 136085 63552 136119
rect 63500 136076 63552 136085
rect 63592 136119 63644 136128
rect 63592 136085 63601 136119
rect 63601 136085 63635 136119
rect 63635 136085 63644 136119
rect 63592 136076 63644 136085
rect 68560 136119 68612 136128
rect 68560 136085 68569 136119
rect 68569 136085 68603 136119
rect 68603 136085 68612 136119
rect 68560 136076 68612 136085
rect 72884 136119 72936 136128
rect 72884 136085 72893 136119
rect 72893 136085 72927 136119
rect 72927 136085 72936 136119
rect 72884 136076 72936 136085
rect 73804 136119 73856 136128
rect 73804 136085 73813 136119
rect 73813 136085 73847 136119
rect 73847 136085 73856 136119
rect 73804 136076 73856 136085
rect 77760 136119 77812 136128
rect 77760 136085 77769 136119
rect 77769 136085 77803 136119
rect 77803 136085 77812 136119
rect 77760 136076 77812 136085
rect 86316 136119 86368 136128
rect 86316 136085 86325 136119
rect 86325 136085 86359 136119
rect 86359 136085 86368 136119
rect 86316 136076 86368 136085
rect 87328 136119 87380 136128
rect 87328 136085 87337 136119
rect 87337 136085 87371 136119
rect 87371 136085 87380 136119
rect 87328 136076 87380 136085
rect 95976 136119 96028 136128
rect 95976 136085 95985 136119
rect 95985 136085 96019 136119
rect 96019 136085 96028 136119
rect 95976 136076 96028 136085
rect 104348 136076 104400 136128
rect 4874 135974 4926 136026
rect 4938 135974 4990 136026
rect 5002 135974 5054 136026
rect 5066 135974 5118 136026
rect 5130 135974 5182 136026
rect 35594 135974 35646 136026
rect 35658 135974 35710 136026
rect 35722 135974 35774 136026
rect 35786 135974 35838 136026
rect 35850 135974 35902 136026
rect 66314 135974 66366 136026
rect 66378 135974 66430 136026
rect 66442 135974 66494 136026
rect 66506 135974 66558 136026
rect 66570 135974 66622 136026
rect 97034 135974 97086 136026
rect 97098 135974 97150 136026
rect 97162 135974 97214 136026
rect 97226 135974 97278 136026
rect 97290 135974 97342 136026
rect 106658 135974 106710 136026
rect 106722 135974 106774 136026
rect 106786 135974 106838 136026
rect 106850 135974 106902 136026
rect 106914 135974 106966 136026
rect 9588 135872 9640 135924
rect 47676 135872 47728 135924
rect 55772 135872 55824 135924
rect 103704 135872 103756 135924
rect 8208 135804 8260 135856
rect 43076 135804 43128 135856
rect 58348 135804 58400 135856
rect 102232 135804 102284 135856
rect 8024 135736 8076 135788
rect 36084 135736 36136 135788
rect 60924 135736 60976 135788
rect 103796 135736 103848 135788
rect 63500 135668 63552 135720
rect 103612 135668 103664 135720
rect 72884 135600 72936 135652
rect 103520 135600 103572 135652
rect 8116 135532 8168 135584
rect 50252 135532 50304 135584
rect 73804 135532 73856 135584
rect 104624 135532 104676 135584
rect 4214 135430 4266 135482
rect 4278 135430 4330 135482
rect 4342 135430 4394 135482
rect 4406 135430 4458 135482
rect 4470 135430 4522 135482
rect 77760 135464 77812 135516
rect 102784 135464 102836 135516
rect 86316 135396 86368 135448
rect 102324 135396 102376 135448
rect 105922 135430 105974 135482
rect 105986 135430 106038 135482
rect 106050 135430 106102 135482
rect 106114 135430 106166 135482
rect 106178 135430 106230 135482
rect 4874 134886 4926 134938
rect 4938 134886 4990 134938
rect 5002 134886 5054 134938
rect 5066 134886 5118 134938
rect 5130 134886 5182 134938
rect 106658 134886 106710 134938
rect 106722 134886 106774 134938
rect 106786 134886 106838 134938
rect 106850 134886 106902 134938
rect 106914 134886 106966 134938
rect 8944 134580 8996 134632
rect 34152 134580 34204 134632
rect 9036 134512 9088 134564
rect 34980 134512 35032 134564
rect 4214 134342 4266 134394
rect 4278 134342 4330 134394
rect 4342 134342 4394 134394
rect 4406 134342 4458 134394
rect 4470 134342 4522 134394
rect 105922 134342 105974 134394
rect 105986 134342 106038 134394
rect 106050 134342 106102 134394
rect 106114 134342 106166 134394
rect 106178 134342 106230 134394
rect 87328 133900 87380 133952
rect 104072 133900 104124 133952
rect 4874 133798 4926 133850
rect 4938 133798 4990 133850
rect 5002 133798 5054 133850
rect 5066 133798 5118 133850
rect 5130 133798 5182 133850
rect 106658 133798 106710 133850
rect 106722 133798 106774 133850
rect 106786 133798 106838 133850
rect 106850 133798 106902 133850
rect 106914 133798 106966 133850
rect 7380 133696 7432 133748
rect 46112 133696 46164 133748
rect 68560 133696 68612 133748
rect 104532 133696 104584 133748
rect 4214 133254 4266 133306
rect 4278 133254 4330 133306
rect 4342 133254 4394 133306
rect 4406 133254 4458 133306
rect 4470 133254 4522 133306
rect 105922 133254 105974 133306
rect 105986 133254 106038 133306
rect 106050 133254 106102 133306
rect 106114 133254 106166 133306
rect 106178 133254 106230 133306
rect 4874 132710 4926 132762
rect 4938 132710 4990 132762
rect 5002 132710 5054 132762
rect 5066 132710 5118 132762
rect 5130 132710 5182 132762
rect 106658 132710 106710 132762
rect 106722 132710 106774 132762
rect 106786 132710 106838 132762
rect 106850 132710 106902 132762
rect 106914 132710 106966 132762
rect 4214 132166 4266 132218
rect 4278 132166 4330 132218
rect 4342 132166 4394 132218
rect 4406 132166 4458 132218
rect 4470 132166 4522 132218
rect 105922 132166 105974 132218
rect 105986 132166 106038 132218
rect 106050 132166 106102 132218
rect 106114 132166 106166 132218
rect 106178 132166 106230 132218
rect 4874 131622 4926 131674
rect 4938 131622 4990 131674
rect 5002 131622 5054 131674
rect 5066 131622 5118 131674
rect 5130 131622 5182 131674
rect 106658 131622 106710 131674
rect 106722 131622 106774 131674
rect 106786 131622 106838 131674
rect 106850 131622 106902 131674
rect 106914 131622 106966 131674
rect 4214 131078 4266 131130
rect 4278 131078 4330 131130
rect 4342 131078 4394 131130
rect 4406 131078 4458 131130
rect 4470 131078 4522 131130
rect 105922 131078 105974 131130
rect 105986 131078 106038 131130
rect 106050 131078 106102 131130
rect 106114 131078 106166 131130
rect 106178 131078 106230 131130
rect 4874 130534 4926 130586
rect 4938 130534 4990 130586
rect 5002 130534 5054 130586
rect 5066 130534 5118 130586
rect 5130 130534 5182 130586
rect 106658 130534 106710 130586
rect 106722 130534 106774 130586
rect 106786 130534 106838 130586
rect 106850 130534 106902 130586
rect 106914 130534 106966 130586
rect 4214 129990 4266 130042
rect 4278 129990 4330 130042
rect 4342 129990 4394 130042
rect 4406 129990 4458 130042
rect 4470 129990 4522 130042
rect 105922 129990 105974 130042
rect 105986 129990 106038 130042
rect 106050 129990 106102 130042
rect 106114 129990 106166 130042
rect 106178 129990 106230 130042
rect 103888 129752 103940 129804
rect 4874 129446 4926 129498
rect 4938 129446 4990 129498
rect 5002 129446 5054 129498
rect 5066 129446 5118 129498
rect 5130 129446 5182 129498
rect 106658 129446 106710 129498
rect 106722 129446 106774 129498
rect 106786 129446 106838 129498
rect 106850 129446 106902 129498
rect 106914 129446 106966 129498
rect 4214 128902 4266 128954
rect 4278 128902 4330 128954
rect 4342 128902 4394 128954
rect 4406 128902 4458 128954
rect 4470 128902 4522 128954
rect 105922 128902 105974 128954
rect 105986 128902 106038 128954
rect 106050 128902 106102 128954
rect 106114 128902 106166 128954
rect 106178 128902 106230 128954
rect 4874 128358 4926 128410
rect 4938 128358 4990 128410
rect 5002 128358 5054 128410
rect 5066 128358 5118 128410
rect 5130 128358 5182 128410
rect 106658 128358 106710 128410
rect 106722 128358 106774 128410
rect 106786 128358 106838 128410
rect 106850 128358 106902 128410
rect 106914 128358 106966 128410
rect 4214 127814 4266 127866
rect 4278 127814 4330 127866
rect 4342 127814 4394 127866
rect 4406 127814 4458 127866
rect 4470 127814 4522 127866
rect 105922 127814 105974 127866
rect 105986 127814 106038 127866
rect 106050 127814 106102 127866
rect 106114 127814 106166 127866
rect 106178 127814 106230 127866
rect 4874 127270 4926 127322
rect 4938 127270 4990 127322
rect 5002 127270 5054 127322
rect 5066 127270 5118 127322
rect 5130 127270 5182 127322
rect 106658 127270 106710 127322
rect 106722 127270 106774 127322
rect 106786 127270 106838 127322
rect 106850 127270 106902 127322
rect 106914 127270 106966 127322
rect 4214 126726 4266 126778
rect 4278 126726 4330 126778
rect 4342 126726 4394 126778
rect 4406 126726 4458 126778
rect 4470 126726 4522 126778
rect 105922 126726 105974 126778
rect 105986 126726 106038 126778
rect 106050 126726 106102 126778
rect 106114 126726 106166 126778
rect 106178 126726 106230 126778
rect 4874 126182 4926 126234
rect 4938 126182 4990 126234
rect 5002 126182 5054 126234
rect 5066 126182 5118 126234
rect 5130 126182 5182 126234
rect 106658 126182 106710 126234
rect 106722 126182 106774 126234
rect 106786 126182 106838 126234
rect 106850 126182 106902 126234
rect 106914 126182 106966 126234
rect 4214 125638 4266 125690
rect 4278 125638 4330 125690
rect 4342 125638 4394 125690
rect 4406 125638 4458 125690
rect 4470 125638 4522 125690
rect 105922 125638 105974 125690
rect 105986 125638 106038 125690
rect 106050 125638 106102 125690
rect 106114 125638 106166 125690
rect 106178 125638 106230 125690
rect 4874 125094 4926 125146
rect 4938 125094 4990 125146
rect 5002 125094 5054 125146
rect 5066 125094 5118 125146
rect 5130 125094 5182 125146
rect 106658 125094 106710 125146
rect 106722 125094 106774 125146
rect 106786 125094 106838 125146
rect 106850 125094 106902 125146
rect 106914 125094 106966 125146
rect 4214 124550 4266 124602
rect 4278 124550 4330 124602
rect 4342 124550 4394 124602
rect 4406 124550 4458 124602
rect 4470 124550 4522 124602
rect 105922 124550 105974 124602
rect 105986 124550 106038 124602
rect 106050 124550 106102 124602
rect 106114 124550 106166 124602
rect 106178 124550 106230 124602
rect 4874 124006 4926 124058
rect 4938 124006 4990 124058
rect 5002 124006 5054 124058
rect 5066 124006 5118 124058
rect 5130 124006 5182 124058
rect 106658 124006 106710 124058
rect 106722 124006 106774 124058
rect 106786 124006 106838 124058
rect 106850 124006 106902 124058
rect 106914 124006 106966 124058
rect 4214 123462 4266 123514
rect 4278 123462 4330 123514
rect 4342 123462 4394 123514
rect 4406 123462 4458 123514
rect 4470 123462 4522 123514
rect 105922 123462 105974 123514
rect 105986 123462 106038 123514
rect 106050 123462 106102 123514
rect 106114 123462 106166 123514
rect 106178 123462 106230 123514
rect 4874 122918 4926 122970
rect 4938 122918 4990 122970
rect 5002 122918 5054 122970
rect 5066 122918 5118 122970
rect 5130 122918 5182 122970
rect 106658 122918 106710 122970
rect 106722 122918 106774 122970
rect 106786 122918 106838 122970
rect 106850 122918 106902 122970
rect 106914 122918 106966 122970
rect 4214 122374 4266 122426
rect 4278 122374 4330 122426
rect 4342 122374 4394 122426
rect 4406 122374 4458 122426
rect 4470 122374 4522 122426
rect 105922 122374 105974 122426
rect 105986 122374 106038 122426
rect 106050 122374 106102 122426
rect 106114 122374 106166 122426
rect 106178 122374 106230 122426
rect 4874 121830 4926 121882
rect 4938 121830 4990 121882
rect 5002 121830 5054 121882
rect 5066 121830 5118 121882
rect 5130 121830 5182 121882
rect 106658 121830 106710 121882
rect 106722 121830 106774 121882
rect 106786 121830 106838 121882
rect 106850 121830 106902 121882
rect 106914 121830 106966 121882
rect 4214 121286 4266 121338
rect 4278 121286 4330 121338
rect 4342 121286 4394 121338
rect 4406 121286 4458 121338
rect 4470 121286 4522 121338
rect 105922 121286 105974 121338
rect 105986 121286 106038 121338
rect 106050 121286 106102 121338
rect 106114 121286 106166 121338
rect 106178 121286 106230 121338
rect 4874 120742 4926 120794
rect 4938 120742 4990 120794
rect 5002 120742 5054 120794
rect 5066 120742 5118 120794
rect 5130 120742 5182 120794
rect 106658 120742 106710 120794
rect 106722 120742 106774 120794
rect 106786 120742 106838 120794
rect 106850 120742 106902 120794
rect 106914 120742 106966 120794
rect 4214 120198 4266 120250
rect 4278 120198 4330 120250
rect 4342 120198 4394 120250
rect 4406 120198 4458 120250
rect 4470 120198 4522 120250
rect 105922 120198 105974 120250
rect 105986 120198 106038 120250
rect 106050 120198 106102 120250
rect 106114 120198 106166 120250
rect 106178 120198 106230 120250
rect 4874 119654 4926 119706
rect 4938 119654 4990 119706
rect 5002 119654 5054 119706
rect 5066 119654 5118 119706
rect 5130 119654 5182 119706
rect 106658 119654 106710 119706
rect 106722 119654 106774 119706
rect 106786 119654 106838 119706
rect 106850 119654 106902 119706
rect 106914 119654 106966 119706
rect 4214 119110 4266 119162
rect 4278 119110 4330 119162
rect 4342 119110 4394 119162
rect 4406 119110 4458 119162
rect 4470 119110 4522 119162
rect 105922 119110 105974 119162
rect 105986 119110 106038 119162
rect 106050 119110 106102 119162
rect 106114 119110 106166 119162
rect 106178 119110 106230 119162
rect 4874 118566 4926 118618
rect 4938 118566 4990 118618
rect 5002 118566 5054 118618
rect 5066 118566 5118 118618
rect 5130 118566 5182 118618
rect 106658 118566 106710 118618
rect 106722 118566 106774 118618
rect 106786 118566 106838 118618
rect 106850 118566 106902 118618
rect 106914 118566 106966 118618
rect 7380 118464 7432 118516
rect 4214 118022 4266 118074
rect 4278 118022 4330 118074
rect 4342 118022 4394 118074
rect 4406 118022 4458 118074
rect 4470 118022 4522 118074
rect 105922 118022 105974 118074
rect 105986 118022 106038 118074
rect 106050 118022 106102 118074
rect 106114 118022 106166 118074
rect 106178 118022 106230 118074
rect 7472 117716 7524 117768
rect 7380 117648 7432 117700
rect 7288 117580 7340 117632
rect 4874 117478 4926 117530
rect 4938 117478 4990 117530
rect 5002 117478 5054 117530
rect 5066 117478 5118 117530
rect 5130 117478 5182 117530
rect 106658 117478 106710 117530
rect 106722 117478 106774 117530
rect 106786 117478 106838 117530
rect 106850 117478 106902 117530
rect 106914 117478 106966 117530
rect 7288 117079 7340 117088
rect 7288 117045 7297 117079
rect 7297 117045 7331 117079
rect 7331 117045 7340 117079
rect 7288 117036 7340 117045
rect 7472 117079 7524 117088
rect 7472 117045 7481 117079
rect 7481 117045 7515 117079
rect 7515 117045 7524 117079
rect 7472 117036 7524 117045
rect 4214 116934 4266 116986
rect 4278 116934 4330 116986
rect 4342 116934 4394 116986
rect 4406 116934 4458 116986
rect 4470 116934 4522 116986
rect 105922 116934 105974 116986
rect 105986 116934 106038 116986
rect 106050 116934 106102 116986
rect 106114 116934 106166 116986
rect 106178 116934 106230 116986
rect 4874 116390 4926 116442
rect 4938 116390 4990 116442
rect 5002 116390 5054 116442
rect 5066 116390 5118 116442
rect 5130 116390 5182 116442
rect 106658 116390 106710 116442
rect 106722 116390 106774 116442
rect 106786 116390 106838 116442
rect 106850 116390 106902 116442
rect 106914 116390 106966 116442
rect 4214 115846 4266 115898
rect 4278 115846 4330 115898
rect 4342 115846 4394 115898
rect 4406 115846 4458 115898
rect 4470 115846 4522 115898
rect 105922 115846 105974 115898
rect 105986 115846 106038 115898
rect 106050 115846 106102 115898
rect 106114 115846 106166 115898
rect 106178 115846 106230 115898
rect 4874 115302 4926 115354
rect 4938 115302 4990 115354
rect 5002 115302 5054 115354
rect 5066 115302 5118 115354
rect 5130 115302 5182 115354
rect 106658 115302 106710 115354
rect 106722 115302 106774 115354
rect 106786 115302 106838 115354
rect 106850 115302 106902 115354
rect 106914 115302 106966 115354
rect 4214 114758 4266 114810
rect 4278 114758 4330 114810
rect 4342 114758 4394 114810
rect 4406 114758 4458 114810
rect 4470 114758 4522 114810
rect 105922 114758 105974 114810
rect 105986 114758 106038 114810
rect 106050 114758 106102 114810
rect 106114 114758 106166 114810
rect 106178 114758 106230 114810
rect 4874 114214 4926 114266
rect 4938 114214 4990 114266
rect 5002 114214 5054 114266
rect 5066 114214 5118 114266
rect 5130 114214 5182 114266
rect 106658 114214 106710 114266
rect 106722 114214 106774 114266
rect 106786 114214 106838 114266
rect 106850 114214 106902 114266
rect 106914 114214 106966 114266
rect 4214 113670 4266 113722
rect 4278 113670 4330 113722
rect 4342 113670 4394 113722
rect 4406 113670 4458 113722
rect 4470 113670 4522 113722
rect 105922 113670 105974 113722
rect 105986 113670 106038 113722
rect 106050 113670 106102 113722
rect 106114 113670 106166 113722
rect 106178 113670 106230 113722
rect 104348 113568 104400 113620
rect 105636 113568 105688 113620
rect 104348 113475 104400 113484
rect 104348 113441 104357 113475
rect 104357 113441 104391 113475
rect 104391 113441 104400 113475
rect 104348 113432 104400 113441
rect 104532 113296 104584 113348
rect 102876 113228 102928 113280
rect 4874 113126 4926 113178
rect 4938 113126 4990 113178
rect 5002 113126 5054 113178
rect 5066 113126 5118 113178
rect 5130 113126 5182 113178
rect 106658 113126 106710 113178
rect 106722 113126 106774 113178
rect 106786 113126 106838 113178
rect 106850 113126 106902 113178
rect 106914 113126 106966 113178
rect 104532 113024 104584 113076
rect 4214 112582 4266 112634
rect 4278 112582 4330 112634
rect 4342 112582 4394 112634
rect 4406 112582 4458 112634
rect 4470 112582 4522 112634
rect 105922 112582 105974 112634
rect 105986 112582 106038 112634
rect 106050 112582 106102 112634
rect 106114 112582 106166 112634
rect 106178 112582 106230 112634
rect 4874 112038 4926 112090
rect 4938 112038 4990 112090
rect 5002 112038 5054 112090
rect 5066 112038 5118 112090
rect 5130 112038 5182 112090
rect 106658 112038 106710 112090
rect 106722 112038 106774 112090
rect 106786 112038 106838 112090
rect 106850 112038 106902 112090
rect 106914 112038 106966 112090
rect 4214 111494 4266 111546
rect 4278 111494 4330 111546
rect 4342 111494 4394 111546
rect 4406 111494 4458 111546
rect 4470 111494 4522 111546
rect 105922 111494 105974 111546
rect 105986 111494 106038 111546
rect 106050 111494 106102 111546
rect 106114 111494 106166 111546
rect 106178 111494 106230 111546
rect 9496 111324 9548 111376
rect 1308 111188 1360 111240
rect 4874 110950 4926 111002
rect 4938 110950 4990 111002
rect 5002 110950 5054 111002
rect 5066 110950 5118 111002
rect 5130 110950 5182 111002
rect 106658 110950 106710 111002
rect 106722 110950 106774 111002
rect 106786 110950 106838 111002
rect 106850 110950 106902 111002
rect 106914 110950 106966 111002
rect 4214 110406 4266 110458
rect 4278 110406 4330 110458
rect 4342 110406 4394 110458
rect 4406 110406 4458 110458
rect 4470 110406 4522 110458
rect 105922 110406 105974 110458
rect 105986 110406 106038 110458
rect 106050 110406 106102 110458
rect 106114 110406 106166 110458
rect 106178 110406 106230 110458
rect 4874 109862 4926 109914
rect 4938 109862 4990 109914
rect 5002 109862 5054 109914
rect 5066 109862 5118 109914
rect 5130 109862 5182 109914
rect 106658 109862 106710 109914
rect 106722 109862 106774 109914
rect 106786 109862 106838 109914
rect 106850 109862 106902 109914
rect 106914 109862 106966 109914
rect 1308 109624 1360 109676
rect 9496 109488 9548 109540
rect 4214 109318 4266 109370
rect 4278 109318 4330 109370
rect 4342 109318 4394 109370
rect 4406 109318 4458 109370
rect 4470 109318 4522 109370
rect 105922 109318 105974 109370
rect 105986 109318 106038 109370
rect 106050 109318 106102 109370
rect 106114 109318 106166 109370
rect 106178 109318 106230 109370
rect 4874 108774 4926 108826
rect 4938 108774 4990 108826
rect 5002 108774 5054 108826
rect 5066 108774 5118 108826
rect 5130 108774 5182 108826
rect 106658 108774 106710 108826
rect 106722 108774 106774 108826
rect 106786 108774 106838 108826
rect 106850 108774 106902 108826
rect 106914 108774 106966 108826
rect 1308 108536 1360 108588
rect 9496 108400 9548 108452
rect 4214 108230 4266 108282
rect 4278 108230 4330 108282
rect 4342 108230 4394 108282
rect 4406 108230 4458 108282
rect 4470 108230 4522 108282
rect 105922 108230 105974 108282
rect 105986 108230 106038 108282
rect 106050 108230 106102 108282
rect 106114 108230 106166 108282
rect 106178 108230 106230 108282
rect 4874 107686 4926 107738
rect 4938 107686 4990 107738
rect 5002 107686 5054 107738
rect 5066 107686 5118 107738
rect 5130 107686 5182 107738
rect 106658 107686 106710 107738
rect 106722 107686 106774 107738
rect 106786 107686 106838 107738
rect 106850 107686 106902 107738
rect 106914 107686 106966 107738
rect 4214 107142 4266 107194
rect 4278 107142 4330 107194
rect 4342 107142 4394 107194
rect 4406 107142 4458 107194
rect 4470 107142 4522 107194
rect 105922 107142 105974 107194
rect 105986 107142 106038 107194
rect 106050 107142 106102 107194
rect 106114 107142 106166 107194
rect 106178 107142 106230 107194
rect 105636 107083 105688 107092
rect 105636 107049 105645 107083
rect 105645 107049 105679 107083
rect 105679 107049 105688 107083
rect 105636 107040 105688 107049
rect 105820 107040 105872 107092
rect 9496 106972 9548 107024
rect 1216 106836 1268 106888
rect 105084 106768 105136 106820
rect 4874 106598 4926 106650
rect 4938 106598 4990 106650
rect 5002 106598 5054 106650
rect 5066 106598 5118 106650
rect 5130 106598 5182 106650
rect 106658 106598 106710 106650
rect 106722 106598 106774 106650
rect 106786 106598 106838 106650
rect 106850 106598 106902 106650
rect 106914 106598 106966 106650
rect 4214 106054 4266 106106
rect 4278 106054 4330 106106
rect 4342 106054 4394 106106
rect 4406 106054 4458 106106
rect 4470 106054 4522 106106
rect 105922 106054 105974 106106
rect 105986 106054 106038 106106
rect 106050 106054 106102 106106
rect 106114 106054 106166 106106
rect 106178 106054 106230 106106
rect 9496 105884 9548 105936
rect 1308 105748 1360 105800
rect 4874 105510 4926 105562
rect 4938 105510 4990 105562
rect 5002 105510 5054 105562
rect 5066 105510 5118 105562
rect 5130 105510 5182 105562
rect 106658 105510 106710 105562
rect 106722 105510 106774 105562
rect 106786 105510 106838 105562
rect 106850 105510 106902 105562
rect 106914 105510 106966 105562
rect 4214 104966 4266 105018
rect 4278 104966 4330 105018
rect 4342 104966 4394 105018
rect 4406 104966 4458 105018
rect 4470 104966 4522 105018
rect 105922 104966 105974 105018
rect 105986 104966 106038 105018
rect 106050 104966 106102 105018
rect 106114 104966 106166 105018
rect 106178 104966 106230 105018
rect 4874 104422 4926 104474
rect 4938 104422 4990 104474
rect 5002 104422 5054 104474
rect 5066 104422 5118 104474
rect 5130 104422 5182 104474
rect 106658 104422 106710 104474
rect 106722 104422 106774 104474
rect 106786 104422 106838 104474
rect 106850 104422 106902 104474
rect 106914 104422 106966 104474
rect 1308 104184 1360 104236
rect 9496 104048 9548 104100
rect 4214 103878 4266 103930
rect 4278 103878 4330 103930
rect 4342 103878 4394 103930
rect 4406 103878 4458 103930
rect 4470 103878 4522 103930
rect 105922 103878 105974 103930
rect 105986 103878 106038 103930
rect 106050 103878 106102 103930
rect 106114 103878 106166 103930
rect 106178 103878 106230 103930
rect 4874 103334 4926 103386
rect 4938 103334 4990 103386
rect 5002 103334 5054 103386
rect 5066 103334 5118 103386
rect 5130 103334 5182 103386
rect 106658 103334 106710 103386
rect 106722 103334 106774 103386
rect 106786 103334 106838 103386
rect 106850 103334 106902 103386
rect 106914 103334 106966 103386
rect 4214 102790 4266 102842
rect 4278 102790 4330 102842
rect 4342 102790 4394 102842
rect 4406 102790 4458 102842
rect 4470 102790 4522 102842
rect 105922 102790 105974 102842
rect 105986 102790 106038 102842
rect 106050 102790 106102 102842
rect 106114 102790 106166 102842
rect 106178 102790 106230 102842
rect 4874 102246 4926 102298
rect 4938 102246 4990 102298
rect 5002 102246 5054 102298
rect 5066 102246 5118 102298
rect 5130 102246 5182 102298
rect 106658 102246 106710 102298
rect 106722 102246 106774 102298
rect 106786 102246 106838 102298
rect 106850 102246 106902 102298
rect 106914 102246 106966 102298
rect 7288 102144 7340 102196
rect 9128 102144 9180 102196
rect 4214 101702 4266 101754
rect 4278 101702 4330 101754
rect 4342 101702 4394 101754
rect 4406 101702 4458 101754
rect 4470 101702 4522 101754
rect 105922 101702 105974 101754
rect 105986 101702 106038 101754
rect 106050 101702 106102 101754
rect 106114 101702 106166 101754
rect 106178 101702 106230 101754
rect 4874 101158 4926 101210
rect 4938 101158 4990 101210
rect 5002 101158 5054 101210
rect 5066 101158 5118 101210
rect 5130 101158 5182 101210
rect 106658 101158 106710 101210
rect 106722 101158 106774 101210
rect 106786 101158 106838 101210
rect 106850 101158 106902 101210
rect 106914 101158 106966 101210
rect 7380 101056 7432 101108
rect 9036 101056 9088 101108
rect 104624 101031 104676 101040
rect 104624 100997 104658 101031
rect 104658 100997 104676 101031
rect 104624 100988 104676 100997
rect 105820 100852 105872 100904
rect 105636 100784 105688 100836
rect 105820 100759 105872 100768
rect 105820 100725 105829 100759
rect 105829 100725 105863 100759
rect 105863 100725 105872 100759
rect 105820 100716 105872 100725
rect 4214 100614 4266 100666
rect 4278 100614 4330 100666
rect 4342 100614 4394 100666
rect 4406 100614 4458 100666
rect 4470 100614 4522 100666
rect 105922 100614 105974 100666
rect 105986 100614 106038 100666
rect 106050 100614 106102 100666
rect 106114 100614 106166 100666
rect 106178 100614 106230 100666
rect 104624 100512 104676 100564
rect 7472 100308 7524 100360
rect 7380 100240 7432 100292
rect 7288 100172 7340 100224
rect 4874 100070 4926 100122
rect 4938 100070 4990 100122
rect 5002 100070 5054 100122
rect 5066 100070 5118 100122
rect 5130 100070 5182 100122
rect 106658 100070 106710 100122
rect 106722 100070 106774 100122
rect 106786 100070 106838 100122
rect 106850 100070 106902 100122
rect 106914 100070 106966 100122
rect 7472 100011 7524 100020
rect 7472 99977 7481 100011
rect 7481 99977 7515 100011
rect 7515 99977 7524 100011
rect 7472 99968 7524 99977
rect 7288 99671 7340 99680
rect 7288 99637 7297 99671
rect 7297 99637 7331 99671
rect 7331 99637 7340 99671
rect 7288 99628 7340 99637
rect 4214 99526 4266 99578
rect 4278 99526 4330 99578
rect 4342 99526 4394 99578
rect 4406 99526 4458 99578
rect 4470 99526 4522 99578
rect 105922 99526 105974 99578
rect 105986 99526 106038 99578
rect 106050 99526 106102 99578
rect 106114 99526 106166 99578
rect 106178 99526 106230 99578
rect 4874 98982 4926 99034
rect 4938 98982 4990 99034
rect 5002 98982 5054 99034
rect 5066 98982 5118 99034
rect 5130 98982 5182 99034
rect 106658 98982 106710 99034
rect 106722 98982 106774 99034
rect 106786 98982 106838 99034
rect 106850 98982 106902 99034
rect 106914 98982 106966 99034
rect 4214 98438 4266 98490
rect 4278 98438 4330 98490
rect 4342 98438 4394 98490
rect 4406 98438 4458 98490
rect 4470 98438 4522 98490
rect 105922 98438 105974 98490
rect 105986 98438 106038 98490
rect 106050 98438 106102 98490
rect 106114 98438 106166 98490
rect 106178 98438 106230 98490
rect 4874 97894 4926 97946
rect 4938 97894 4990 97946
rect 5002 97894 5054 97946
rect 5066 97894 5118 97946
rect 5130 97894 5182 97946
rect 106658 97894 106710 97946
rect 106722 97894 106774 97946
rect 106786 97894 106838 97946
rect 106850 97894 106902 97946
rect 106914 97894 106966 97946
rect 4214 97350 4266 97402
rect 4278 97350 4330 97402
rect 4342 97350 4394 97402
rect 4406 97350 4458 97402
rect 4470 97350 4522 97402
rect 105922 97350 105974 97402
rect 105986 97350 106038 97402
rect 106050 97350 106102 97402
rect 106114 97350 106166 97402
rect 106178 97350 106230 97402
rect 4874 96806 4926 96858
rect 4938 96806 4990 96858
rect 5002 96806 5054 96858
rect 5066 96806 5118 96858
rect 5130 96806 5182 96858
rect 106658 96806 106710 96858
rect 106722 96806 106774 96858
rect 106786 96806 106838 96858
rect 106850 96806 106902 96858
rect 106914 96806 106966 96858
rect 102784 96568 102836 96620
rect 4214 96262 4266 96314
rect 4278 96262 4330 96314
rect 4342 96262 4394 96314
rect 4406 96262 4458 96314
rect 4470 96262 4522 96314
rect 104348 96543 104400 96552
rect 104348 96509 104357 96543
rect 104357 96509 104391 96543
rect 104391 96509 104400 96543
rect 104348 96500 104400 96509
rect 104348 96364 104400 96416
rect 105636 96432 105688 96484
rect 105728 96407 105780 96416
rect 105728 96373 105737 96407
rect 105737 96373 105771 96407
rect 105771 96373 105780 96407
rect 105728 96364 105780 96373
rect 105922 96262 105974 96314
rect 105986 96262 106038 96314
rect 106050 96262 106102 96314
rect 106114 96262 106166 96314
rect 106178 96262 106230 96314
rect 102968 96092 103020 96144
rect 105728 96092 105780 96144
rect 4874 95718 4926 95770
rect 4938 95718 4990 95770
rect 5002 95718 5054 95770
rect 5066 95718 5118 95770
rect 5130 95718 5182 95770
rect 106658 95718 106710 95770
rect 106722 95718 106774 95770
rect 106786 95718 106838 95770
rect 106850 95718 106902 95770
rect 106914 95718 106966 95770
rect 7472 95659 7524 95668
rect 7472 95625 7481 95659
rect 7481 95625 7515 95659
rect 7515 95625 7524 95659
rect 7472 95616 7524 95625
rect 4214 95174 4266 95226
rect 4278 95174 4330 95226
rect 4342 95174 4394 95226
rect 4406 95174 4458 95226
rect 4470 95174 4522 95226
rect 102508 95140 102560 95192
rect 105922 95174 105974 95226
rect 105986 95174 106038 95226
rect 106050 95174 106102 95226
rect 106114 95174 106166 95226
rect 106178 95174 106230 95226
rect 7472 94979 7524 94988
rect 7472 94945 7481 94979
rect 7481 94945 7515 94979
rect 7515 94945 7524 94979
rect 7472 94936 7524 94945
rect 5816 94843 5868 94852
rect 5816 94809 5825 94843
rect 5825 94809 5859 94843
rect 5859 94809 5868 94843
rect 5816 94800 5868 94809
rect 4874 94630 4926 94682
rect 4938 94630 4990 94682
rect 5002 94630 5054 94682
rect 5066 94630 5118 94682
rect 5130 94630 5182 94682
rect 106658 94630 106710 94682
rect 106722 94630 106774 94682
rect 106786 94630 106838 94682
rect 106850 94630 106902 94682
rect 106914 94630 106966 94682
rect 7472 94392 7524 94444
rect 4214 94086 4266 94138
rect 4278 94086 4330 94138
rect 4342 94086 4394 94138
rect 4406 94086 4458 94138
rect 4470 94086 4522 94138
rect 105922 94086 105974 94138
rect 105986 94086 106038 94138
rect 106050 94086 106102 94138
rect 106114 94086 106166 94138
rect 106178 94086 106230 94138
rect 7472 93780 7524 93832
rect 7104 93644 7156 93696
rect 4874 93542 4926 93594
rect 4938 93542 4990 93594
rect 5002 93542 5054 93594
rect 5066 93542 5118 93594
rect 5130 93542 5182 93594
rect 8944 93712 8996 93764
rect 102416 93644 102468 93696
rect 106658 93542 106710 93594
rect 106722 93542 106774 93594
rect 106786 93542 106838 93594
rect 106850 93542 106902 93594
rect 106914 93542 106966 93594
rect 7104 93143 7156 93152
rect 7104 93109 7113 93143
rect 7113 93109 7147 93143
rect 7147 93109 7156 93143
rect 7104 93100 7156 93109
rect 7472 93143 7524 93152
rect 7472 93109 7481 93143
rect 7481 93109 7515 93143
rect 7515 93109 7524 93143
rect 7472 93100 7524 93109
rect 4214 92998 4266 93050
rect 4278 92998 4330 93050
rect 4342 92998 4394 93050
rect 4406 92998 4458 93050
rect 4470 92998 4522 93050
rect 105922 92998 105974 93050
rect 105986 92998 106038 93050
rect 106050 92998 106102 93050
rect 106114 92998 106166 93050
rect 106178 92998 106230 93050
rect 103888 92556 103940 92608
rect 4874 92454 4926 92506
rect 4938 92454 4990 92506
rect 5002 92454 5054 92506
rect 5066 92454 5118 92506
rect 5130 92454 5182 92506
rect 106658 92454 106710 92506
rect 106722 92454 106774 92506
rect 106786 92454 106838 92506
rect 106850 92454 106902 92506
rect 106914 92454 106966 92506
rect 4214 91910 4266 91962
rect 4278 91910 4330 91962
rect 4342 91910 4394 91962
rect 4406 91910 4458 91962
rect 4470 91910 4522 91962
rect 105922 91910 105974 91962
rect 105986 91910 106038 91962
rect 106050 91910 106102 91962
rect 106114 91910 106166 91962
rect 106178 91910 106230 91962
rect 4874 91366 4926 91418
rect 4938 91366 4990 91418
rect 5002 91366 5054 91418
rect 5066 91366 5118 91418
rect 5130 91366 5182 91418
rect 102784 91060 102836 91112
rect 105084 91579 105136 91588
rect 105084 91545 105093 91579
rect 105093 91545 105127 91579
rect 105127 91545 105136 91579
rect 105084 91536 105136 91545
rect 106658 91366 106710 91418
rect 106722 91366 106774 91418
rect 106786 91366 106838 91418
rect 106850 91366 106902 91418
rect 106914 91366 106966 91418
rect 4214 90822 4266 90874
rect 4278 90822 4330 90874
rect 4342 90822 4394 90874
rect 4406 90822 4458 90874
rect 4470 90822 4522 90874
rect 105922 90822 105974 90874
rect 105986 90822 106038 90874
rect 106050 90822 106102 90874
rect 106114 90822 106166 90874
rect 106178 90822 106230 90874
rect 4874 90278 4926 90330
rect 4938 90278 4990 90330
rect 5002 90278 5054 90330
rect 5066 90278 5118 90330
rect 5130 90278 5182 90330
rect 106658 90278 106710 90330
rect 106722 90278 106774 90330
rect 106786 90278 106838 90330
rect 106850 90278 106902 90330
rect 106914 90278 106966 90330
rect 4214 89734 4266 89786
rect 4278 89734 4330 89786
rect 4342 89734 4394 89786
rect 4406 89734 4458 89786
rect 4470 89734 4522 89786
rect 105922 89734 105974 89786
rect 105986 89734 106038 89786
rect 106050 89734 106102 89786
rect 106114 89734 106166 89786
rect 106178 89734 106230 89786
rect 4874 89190 4926 89242
rect 4938 89190 4990 89242
rect 5002 89190 5054 89242
rect 5066 89190 5118 89242
rect 5130 89190 5182 89242
rect 106658 89190 106710 89242
rect 106722 89190 106774 89242
rect 106786 89190 106838 89242
rect 106850 89190 106902 89242
rect 106914 89190 106966 89242
rect 1308 88952 1360 89004
rect 7564 88816 7616 88868
rect 4214 88646 4266 88698
rect 4278 88646 4330 88698
rect 4342 88646 4394 88698
rect 4406 88646 4458 88698
rect 4470 88646 4522 88698
rect 105922 88646 105974 88698
rect 105986 88646 106038 88698
rect 106050 88646 106102 88698
rect 106114 88646 106166 88698
rect 106178 88646 106230 88698
rect 4874 88102 4926 88154
rect 4938 88102 4990 88154
rect 5002 88102 5054 88154
rect 5066 88102 5118 88154
rect 5130 88102 5182 88154
rect 106658 88102 106710 88154
rect 106722 88102 106774 88154
rect 106786 88102 106838 88154
rect 106850 88102 106902 88154
rect 106914 88102 106966 88154
rect 1216 87864 1268 87916
rect 8944 87728 8996 87780
rect 4214 87558 4266 87610
rect 4278 87558 4330 87610
rect 4342 87558 4394 87610
rect 4406 87558 4458 87610
rect 4470 87558 4522 87610
rect 105922 87558 105974 87610
rect 105986 87558 106038 87610
rect 106050 87558 106102 87610
rect 106114 87558 106166 87610
rect 106178 87558 106230 87610
rect 1216 87184 1268 87236
rect 1860 87159 1912 87168
rect 1860 87125 1869 87159
rect 1869 87125 1903 87159
rect 1903 87125 1912 87159
rect 1860 87116 1912 87125
rect 4874 87014 4926 87066
rect 4938 87014 4990 87066
rect 5002 87014 5054 87066
rect 5066 87014 5118 87066
rect 5130 87014 5182 87066
rect 106658 87014 106710 87066
rect 106722 87014 106774 87066
rect 106786 87014 106838 87066
rect 106850 87014 106902 87066
rect 106914 87014 106966 87066
rect 1308 86776 1360 86828
rect 8392 86640 8444 86692
rect 4214 86470 4266 86522
rect 4278 86470 4330 86522
rect 4342 86470 4394 86522
rect 4406 86470 4458 86522
rect 4470 86470 4522 86522
rect 105922 86470 105974 86522
rect 105986 86470 106038 86522
rect 106050 86470 106102 86522
rect 106114 86470 106166 86522
rect 106178 86470 106230 86522
rect 1308 86164 1360 86216
rect 5540 86028 5592 86080
rect 4874 85926 4926 85978
rect 4938 85926 4990 85978
rect 5002 85926 5054 85978
rect 5066 85926 5118 85978
rect 5130 85926 5182 85978
rect 106658 85926 106710 85978
rect 106722 85926 106774 85978
rect 106786 85926 106838 85978
rect 106850 85926 106902 85978
rect 106914 85926 106966 85978
rect 1860 85552 1912 85604
rect 8576 85552 8628 85604
rect 4214 85382 4266 85434
rect 4278 85382 4330 85434
rect 4342 85382 4394 85434
rect 4406 85382 4458 85434
rect 4470 85382 4522 85434
rect 105922 85382 105974 85434
rect 105986 85382 106038 85434
rect 106050 85382 106102 85434
rect 106114 85382 106166 85434
rect 106178 85382 106230 85434
rect 1216 85008 1268 85060
rect 2044 84940 2096 84992
rect 4874 84838 4926 84890
rect 4938 84838 4990 84890
rect 5002 84838 5054 84890
rect 5066 84838 5118 84890
rect 5130 84838 5182 84890
rect 106658 84838 106710 84890
rect 106722 84838 106774 84890
rect 106786 84838 106838 84890
rect 106850 84838 106902 84890
rect 106914 84838 106966 84890
rect 1308 84600 1360 84652
rect 1860 84464 1912 84516
rect 4214 84294 4266 84346
rect 4278 84294 4330 84346
rect 4342 84294 4394 84346
rect 4406 84294 4458 84346
rect 4470 84294 4522 84346
rect 105922 84294 105974 84346
rect 105986 84294 106038 84346
rect 106050 84294 106102 84346
rect 106114 84294 106166 84346
rect 106178 84294 106230 84346
rect 1860 84124 1912 84176
rect 9312 84124 9364 84176
rect 1308 83988 1360 84040
rect 2504 83852 2556 83904
rect 4874 83750 4926 83802
rect 4938 83750 4990 83802
rect 5002 83750 5054 83802
rect 5066 83750 5118 83802
rect 5130 83750 5182 83802
rect 106658 83750 106710 83802
rect 106722 83750 106774 83802
rect 106786 83750 106838 83802
rect 106850 83750 106902 83802
rect 106914 83750 106966 83802
rect 1308 83512 1360 83564
rect 2044 83444 2096 83496
rect 9220 83444 9272 83496
rect 2044 83308 2096 83360
rect 4214 83206 4266 83258
rect 4278 83206 4330 83258
rect 4342 83206 4394 83258
rect 4406 83206 4458 83258
rect 4470 83206 4522 83258
rect 105922 83206 105974 83258
rect 105986 83206 106038 83258
rect 106050 83206 106102 83258
rect 106114 83206 106166 83258
rect 106178 83206 106230 83258
rect 4874 82662 4926 82714
rect 4938 82662 4990 82714
rect 5002 82662 5054 82714
rect 5066 82662 5118 82714
rect 5130 82662 5182 82714
rect 106658 82662 106710 82714
rect 106722 82662 106774 82714
rect 106786 82662 106838 82714
rect 106850 82662 106902 82714
rect 106914 82662 106966 82714
rect 1216 82424 1268 82476
rect 2688 82220 2740 82272
rect 5264 82356 5316 82408
rect 5816 82220 5868 82272
rect 6184 82220 6236 82272
rect 4214 82118 4266 82170
rect 4278 82118 4330 82170
rect 4342 82118 4394 82170
rect 4406 82118 4458 82170
rect 4470 82118 4522 82170
rect 105922 82118 105974 82170
rect 105986 82118 106038 82170
rect 106050 82118 106102 82170
rect 106114 82118 106166 82170
rect 106178 82118 106230 82170
rect 1216 81744 1268 81796
rect 1860 81719 1912 81728
rect 1860 81685 1869 81719
rect 1869 81685 1903 81719
rect 1903 81685 1912 81719
rect 1860 81676 1912 81685
rect 4874 81574 4926 81626
rect 4938 81574 4990 81626
rect 5002 81574 5054 81626
rect 5066 81574 5118 81626
rect 5130 81574 5182 81626
rect 106658 81574 106710 81626
rect 106722 81574 106774 81626
rect 106786 81574 106838 81626
rect 106850 81574 106902 81626
rect 106914 81574 106966 81626
rect 1308 81336 1360 81388
rect 2044 81268 2096 81320
rect 9772 81268 9824 81320
rect 9588 81200 9640 81252
rect 4214 81030 4266 81082
rect 4278 81030 4330 81082
rect 4342 81030 4394 81082
rect 4406 81030 4458 81082
rect 4470 81030 4522 81082
rect 105922 81030 105974 81082
rect 105986 81030 106038 81082
rect 106050 81030 106102 81082
rect 106114 81030 106166 81082
rect 106178 81030 106230 81082
rect 1860 80792 1912 80844
rect 9680 80792 9732 80844
rect 1308 80724 1360 80776
rect 2688 80724 2740 80776
rect 9864 80724 9916 80776
rect 107752 80724 107804 80776
rect 108488 80767 108540 80776
rect 108488 80733 108497 80767
rect 108497 80733 108531 80767
rect 108531 80733 108540 80767
rect 108488 80724 108540 80733
rect 2504 80656 2556 80708
rect 9956 80656 10008 80708
rect 5540 80588 5592 80640
rect 4874 80486 4926 80538
rect 4938 80486 4990 80538
rect 5002 80486 5054 80538
rect 5066 80486 5118 80538
rect 5130 80486 5182 80538
rect 106658 80486 106710 80538
rect 106722 80486 106774 80538
rect 106786 80486 106838 80538
rect 106850 80486 106902 80538
rect 106914 80486 106966 80538
rect 1308 80316 1360 80368
rect 108488 80359 108540 80368
rect 108488 80325 108497 80359
rect 108497 80325 108531 80359
rect 108531 80325 108540 80359
rect 108488 80316 108540 80325
rect 101956 80044 102008 80096
rect 105820 80044 105872 80096
rect 4214 79942 4266 79994
rect 4278 79942 4330 79994
rect 4342 79942 4394 79994
rect 4406 79942 4458 79994
rect 4470 79942 4522 79994
rect 9956 79976 10008 80028
rect 43260 79976 43312 80028
rect 9772 79908 9824 79960
rect 40960 79908 41012 79960
rect 105922 79942 105974 79994
rect 105986 79942 106038 79994
rect 106050 79942 106102 79994
rect 106114 79942 106166 79994
rect 106178 79942 106230 79994
rect 9864 79840 9916 79892
rect 39764 79840 39816 79892
rect 7564 79772 7616 79824
rect 36268 79772 36320 79824
rect 9680 79704 9732 79756
rect 38660 79704 38712 79756
rect 8944 79636 8996 79688
rect 33968 79636 34020 79688
rect 98000 79636 98052 79688
rect 1216 79568 1268 79620
rect 8576 79568 8628 79620
rect 31668 79568 31720 79620
rect 37464 79500 37516 79552
rect 108396 79543 108448 79552
rect 108396 79509 108405 79543
rect 108405 79509 108439 79543
rect 108439 79509 108448 79543
rect 108396 79500 108448 79509
rect 4874 79398 4926 79450
rect 4938 79398 4990 79450
rect 5002 79398 5054 79450
rect 5066 79398 5118 79450
rect 5130 79398 5182 79450
rect 92112 79432 92164 79484
rect 102876 79432 102928 79484
rect 90272 79364 90324 79416
rect 102968 79364 103020 79416
rect 106658 79398 106710 79450
rect 106722 79398 106774 79450
rect 106786 79398 106838 79450
rect 106850 79398 106902 79450
rect 106914 79398 106966 79450
rect 73804 79296 73856 79348
rect 102784 79296 102836 79348
rect 1308 79160 1360 79212
rect 96804 79160 96856 79212
rect 42156 78956 42208 79008
rect 108396 78999 108448 79008
rect 108396 78965 108405 78999
rect 108405 78965 108439 78999
rect 108439 78965 108448 78999
rect 108396 78956 108448 78965
rect 4214 78854 4266 78906
rect 4278 78854 4330 78906
rect 4342 78854 4394 78906
rect 4406 78854 4458 78906
rect 4470 78854 4522 78906
rect 105922 78854 105974 78906
rect 105986 78854 106038 78906
rect 106050 78854 106102 78906
rect 106114 78854 106166 78906
rect 106178 78854 106230 78906
rect 7288 78616 7340 78668
rect 14004 78616 14056 78668
rect 95884 78616 95936 78668
rect 102048 78616 102100 78668
rect 107660 78548 107712 78600
rect 1308 78480 1360 78532
rect 29552 78412 29604 78464
rect 108396 78455 108448 78464
rect 108396 78421 108405 78455
rect 108405 78421 108439 78455
rect 108439 78421 108448 78455
rect 108396 78412 108448 78421
rect 4874 78310 4926 78362
rect 4938 78310 4990 78362
rect 5002 78310 5054 78362
rect 5066 78310 5118 78362
rect 5130 78310 5182 78362
rect 106658 78310 106710 78362
rect 106722 78310 106774 78362
rect 106786 78310 106838 78362
rect 106850 78310 106902 78362
rect 106914 78310 106966 78362
rect 91928 78140 91980 78192
rect 102324 78140 102376 78192
rect 1308 78072 1360 78124
rect 2044 78072 2096 78124
rect 35348 78072 35400 78124
rect 108212 78115 108264 78124
rect 108212 78081 108221 78115
rect 108221 78081 108255 78115
rect 108255 78081 108264 78115
rect 108212 78072 108264 78081
rect 16212 78004 16264 78056
rect 25412 78004 25464 78056
rect 92388 78004 92440 78056
rect 102416 78004 102468 78056
rect 7104 77936 7156 77988
rect 17132 77936 17184 77988
rect 89904 77936 89956 77988
rect 102140 77936 102192 77988
rect 26056 77868 26108 77920
rect 87236 77868 87288 77920
rect 101956 77868 102008 77920
rect 108396 77911 108448 77920
rect 108396 77877 108405 77911
rect 108405 77877 108439 77911
rect 108439 77877 108448 77911
rect 108396 77868 108448 77877
rect 4214 77766 4266 77818
rect 4278 77766 4330 77818
rect 4342 77766 4394 77818
rect 4406 77766 4458 77818
rect 4470 77766 4522 77818
rect 34934 77766 34986 77818
rect 34998 77766 35050 77818
rect 35062 77766 35114 77818
rect 35126 77766 35178 77818
rect 35190 77766 35242 77818
rect 65654 77766 65706 77818
rect 65718 77766 65770 77818
rect 65782 77766 65834 77818
rect 65846 77766 65898 77818
rect 65910 77766 65962 77818
rect 96374 77766 96426 77818
rect 96438 77766 96490 77818
rect 96502 77766 96554 77818
rect 96566 77766 96618 77818
rect 96630 77766 96682 77818
rect 105922 77766 105974 77818
rect 105986 77766 106038 77818
rect 106050 77766 106102 77818
rect 106114 77766 106166 77818
rect 106178 77766 106230 77818
rect 8024 77664 8076 77716
rect 11060 77596 11112 77648
rect 16120 77664 16172 77716
rect 26056 77707 26108 77716
rect 26056 77673 26065 77707
rect 26065 77673 26099 77707
rect 26099 77673 26108 77707
rect 26056 77664 26108 77673
rect 26976 77707 27028 77716
rect 26976 77673 26985 77707
rect 26985 77673 27019 77707
rect 27019 77673 27028 77707
rect 26976 77664 27028 77673
rect 28172 77707 28224 77716
rect 28172 77673 28181 77707
rect 28181 77673 28215 77707
rect 28215 77673 28224 77707
rect 28172 77664 28224 77673
rect 29552 77707 29604 77716
rect 29552 77673 29561 77707
rect 29561 77673 29595 77707
rect 29595 77673 29604 77707
rect 29552 77664 29604 77673
rect 30472 77707 30524 77716
rect 30472 77673 30481 77707
rect 30481 77673 30515 77707
rect 30515 77673 30524 77707
rect 30472 77664 30524 77673
rect 31760 77707 31812 77716
rect 31760 77673 31769 77707
rect 31769 77673 31803 77707
rect 31803 77673 31812 77707
rect 31760 77664 31812 77673
rect 32864 77707 32916 77716
rect 32864 77673 32873 77707
rect 32873 77673 32907 77707
rect 32907 77673 32916 77707
rect 32864 77664 32916 77673
rect 33968 77707 34020 77716
rect 33968 77673 33977 77707
rect 33977 77673 34011 77707
rect 34011 77673 34020 77707
rect 33968 77664 34020 77673
rect 35348 77664 35400 77716
rect 36268 77664 36320 77716
rect 37464 77707 37516 77716
rect 37464 77673 37473 77707
rect 37473 77673 37507 77707
rect 37507 77673 37516 77707
rect 37464 77664 37516 77673
rect 38660 77707 38712 77716
rect 38660 77673 38669 77707
rect 38669 77673 38703 77707
rect 38703 77673 38712 77707
rect 38660 77664 38712 77673
rect 39764 77664 39816 77716
rect 40960 77664 41012 77716
rect 42156 77707 42208 77716
rect 42156 77673 42165 77707
rect 42165 77673 42199 77707
rect 42199 77673 42208 77707
rect 42156 77664 42208 77673
rect 43260 77664 43312 77716
rect 91192 77664 91244 77716
rect 94872 77664 94924 77716
rect 97908 77664 97960 77716
rect 99104 77664 99156 77716
rect 104348 77664 104400 77716
rect 27528 77596 27580 77648
rect 87236 77639 87288 77648
rect 19892 77460 19944 77512
rect 55036 77460 55088 77512
rect 14648 77367 14700 77376
rect 14648 77333 14657 77367
rect 14657 77333 14691 77367
rect 14691 77333 14700 77367
rect 14648 77324 14700 77333
rect 16212 77435 16264 77444
rect 16212 77401 16221 77435
rect 16221 77401 16255 77435
rect 16255 77401 16264 77435
rect 16212 77392 16264 77401
rect 55128 77435 55180 77444
rect 55128 77401 55137 77435
rect 55137 77401 55171 77435
rect 55171 77401 55180 77435
rect 55128 77392 55180 77401
rect 20720 77324 20772 77376
rect 23480 77367 23532 77376
rect 23480 77333 23489 77367
rect 23489 77333 23523 77367
rect 23523 77333 23532 77367
rect 23480 77324 23532 77333
rect 55036 77324 55088 77376
rect 59268 77324 59320 77376
rect 82820 77324 82872 77376
rect 86408 77571 86460 77580
rect 86408 77537 86417 77571
rect 86417 77537 86451 77571
rect 86451 77537 86460 77571
rect 86408 77528 86460 77537
rect 87236 77605 87245 77639
rect 87245 77605 87279 77639
rect 87279 77605 87288 77639
rect 87236 77596 87288 77605
rect 89628 77596 89680 77648
rect 89720 77596 89772 77648
rect 89812 77596 89864 77648
rect 89904 77528 89956 77580
rect 90548 77596 90600 77648
rect 91928 77596 91980 77648
rect 96528 77596 96580 77648
rect 108212 77596 108264 77648
rect 84016 77367 84068 77376
rect 84016 77333 84025 77367
rect 84025 77333 84059 77367
rect 84059 77333 84068 77367
rect 84016 77324 84068 77333
rect 85856 77324 85908 77376
rect 86776 77324 86828 77376
rect 89628 77392 89680 77444
rect 92480 77460 92532 77512
rect 105084 77528 105136 77580
rect 93952 77460 94004 77512
rect 94872 77503 94924 77512
rect 94872 77469 94881 77503
rect 94881 77469 94915 77503
rect 94915 77469 94924 77503
rect 94872 77460 94924 77469
rect 96896 77460 96948 77512
rect 91468 77435 91520 77444
rect 91468 77401 91477 77435
rect 91477 77401 91511 77435
rect 91511 77401 91520 77435
rect 91468 77392 91520 77401
rect 92020 77392 92072 77444
rect 95240 77392 95292 77444
rect 97908 77392 97960 77444
rect 89812 77324 89864 77376
rect 90088 77324 90140 77376
rect 91560 77367 91612 77376
rect 91560 77333 91569 77367
rect 91569 77333 91603 77367
rect 91603 77333 91612 77367
rect 91560 77324 91612 77333
rect 92204 77324 92256 77376
rect 92572 77324 92624 77376
rect 93952 77324 94004 77376
rect 97632 77324 97684 77376
rect 99104 77367 99156 77376
rect 99104 77333 99113 77367
rect 99113 77333 99147 77367
rect 99147 77333 99156 77367
rect 99104 77324 99156 77333
rect 4874 77222 4926 77274
rect 4938 77222 4990 77274
rect 5002 77222 5054 77274
rect 5066 77222 5118 77274
rect 5130 77222 5182 77274
rect 35594 77222 35646 77274
rect 35658 77222 35710 77274
rect 35722 77222 35774 77274
rect 35786 77222 35838 77274
rect 35850 77222 35902 77274
rect 66314 77222 66366 77274
rect 66378 77222 66430 77274
rect 66442 77222 66494 77274
rect 66506 77222 66558 77274
rect 66570 77222 66622 77274
rect 97034 77222 97086 77274
rect 97098 77222 97150 77274
rect 97162 77222 97214 77274
rect 97226 77222 97278 77274
rect 97290 77222 97342 77274
rect 106658 77222 106710 77274
rect 106722 77222 106774 77274
rect 106786 77222 106838 77274
rect 106850 77222 106902 77274
rect 106914 77222 106966 77274
rect 2044 77120 2096 77172
rect 8116 77120 8168 77172
rect 46940 77120 46992 77172
rect 86408 77120 86460 77172
rect 20720 77052 20772 77104
rect 24676 77095 24728 77104
rect 24676 77061 24685 77095
rect 24685 77061 24719 77095
rect 24719 77061 24728 77095
rect 24676 77052 24728 77061
rect 25228 77052 25280 77104
rect 1216 76984 1268 77036
rect 22468 77027 22520 77036
rect 22468 76993 22477 77027
rect 22477 76993 22511 77027
rect 22511 76993 22520 77027
rect 22468 76984 22520 76993
rect 8208 76916 8260 76968
rect 9128 76848 9180 76900
rect 25228 76891 25280 76900
rect 25228 76857 25237 76891
rect 25237 76857 25271 76891
rect 25271 76857 25280 76891
rect 25228 76848 25280 76857
rect 32956 76984 33008 77036
rect 26332 76916 26384 76968
rect 89720 77120 89772 77172
rect 90364 77120 90416 77172
rect 95240 77120 95292 77172
rect 88432 76984 88484 77036
rect 90272 76984 90324 77036
rect 90364 77027 90416 77036
rect 90364 76993 90373 77027
rect 90373 76993 90407 77027
rect 90407 76993 90416 77027
rect 90364 76984 90416 76993
rect 90548 77027 90600 77036
rect 90548 76993 90557 77027
rect 90557 76993 90591 77027
rect 90591 76993 90600 77027
rect 90548 76984 90600 76993
rect 41328 76848 41380 76900
rect 89260 76916 89312 76968
rect 91928 77027 91980 77036
rect 91928 76993 91937 77027
rect 91937 76993 91971 77027
rect 91971 76993 91980 77027
rect 91928 76984 91980 76993
rect 92112 77027 92164 77036
rect 92112 76993 92121 77027
rect 92121 76993 92155 77027
rect 92155 76993 92164 77027
rect 92112 76984 92164 76993
rect 22376 76780 22428 76832
rect 25412 76823 25464 76832
rect 25412 76789 25421 76823
rect 25421 76789 25455 76823
rect 25455 76789 25464 76823
rect 25412 76780 25464 76789
rect 26332 76823 26384 76832
rect 26332 76789 26341 76823
rect 26341 76789 26375 76823
rect 26375 76789 26384 76823
rect 26332 76780 26384 76789
rect 55036 76823 55088 76832
rect 55036 76789 55045 76823
rect 55045 76789 55079 76823
rect 55079 76789 55088 76823
rect 55036 76780 55088 76789
rect 90456 76823 90508 76832
rect 90456 76789 90465 76823
rect 90465 76789 90499 76823
rect 90499 76789 90508 76823
rect 90456 76780 90508 76789
rect 92572 76780 92624 76832
rect 93952 77027 94004 77036
rect 93952 76993 93961 77027
rect 93961 76993 93995 77027
rect 93995 76993 94004 77027
rect 96896 77120 96948 77172
rect 97632 77163 97684 77172
rect 97632 77129 97641 77163
rect 97641 77129 97675 77163
rect 97675 77129 97684 77163
rect 97632 77120 97684 77129
rect 96528 77052 96580 77104
rect 98736 77052 98788 77104
rect 93952 76984 94004 76993
rect 99104 77027 99156 77036
rect 99104 76993 99113 77027
rect 99113 76993 99147 77027
rect 99147 76993 99156 77027
rect 99104 76984 99156 76993
rect 99288 77027 99340 77036
rect 99288 76993 99297 77027
rect 99297 76993 99331 77027
rect 99331 76993 99340 77027
rect 99288 76984 99340 76993
rect 99196 76916 99248 76968
rect 100116 76984 100168 77036
rect 100760 76984 100812 77036
rect 100576 76916 100628 76968
rect 107660 76848 107712 76900
rect 108396 76891 108448 76900
rect 108396 76857 108405 76891
rect 108405 76857 108439 76891
rect 108439 76857 108448 76891
rect 108396 76848 108448 76857
rect 94044 76823 94096 76832
rect 94044 76789 94053 76823
rect 94053 76789 94087 76823
rect 94087 76789 94096 76823
rect 94044 76780 94096 76789
rect 98460 76780 98512 76832
rect 101036 76780 101088 76832
rect 4214 76678 4266 76730
rect 4278 76678 4330 76730
rect 4342 76678 4394 76730
rect 4406 76678 4458 76730
rect 4470 76678 4522 76730
rect 34934 76678 34986 76730
rect 34998 76678 35050 76730
rect 35062 76678 35114 76730
rect 35126 76678 35178 76730
rect 35190 76678 35242 76730
rect 65654 76678 65706 76730
rect 65718 76678 65770 76730
rect 65782 76678 65834 76730
rect 65846 76678 65898 76730
rect 65910 76678 65962 76730
rect 96374 76678 96426 76730
rect 96438 76678 96490 76730
rect 96502 76678 96554 76730
rect 96566 76678 96618 76730
rect 96630 76678 96682 76730
rect 9404 76576 9456 76628
rect 19340 76508 19392 76560
rect 14004 76440 14056 76492
rect 26332 76440 26384 76492
rect 14556 76372 14608 76424
rect 17132 76372 17184 76424
rect 27528 76440 27580 76492
rect 41328 76619 41380 76628
rect 41328 76585 41337 76619
rect 41337 76585 41371 76619
rect 41371 76585 41380 76619
rect 41328 76576 41380 76585
rect 46940 76619 46992 76628
rect 46940 76585 46949 76619
rect 46949 76585 46983 76619
rect 46983 76585 46992 76619
rect 46940 76576 46992 76585
rect 58624 76576 58676 76628
rect 59268 76576 59320 76628
rect 68928 76576 68980 76628
rect 92480 76576 92532 76628
rect 98000 76576 98052 76628
rect 99104 76576 99156 76628
rect 95424 76508 95476 76560
rect 99288 76508 99340 76560
rect 82544 76440 82596 76492
rect 82728 76440 82780 76492
rect 85856 76440 85908 76492
rect 98276 76440 98328 76492
rect 848 76236 900 76288
rect 23572 76279 23624 76288
rect 23572 76245 23581 76279
rect 23581 76245 23615 76279
rect 23615 76245 23624 76279
rect 23572 76236 23624 76245
rect 24860 76236 24912 76288
rect 28448 76236 28500 76288
rect 28540 76279 28592 76288
rect 28540 76245 28549 76279
rect 28549 76245 28583 76279
rect 28583 76245 28592 76279
rect 28540 76236 28592 76245
rect 30288 76304 30340 76356
rect 55036 76372 55088 76424
rect 86868 76372 86920 76424
rect 33048 76236 33100 76288
rect 39856 76279 39908 76288
rect 39856 76245 39865 76279
rect 39865 76245 39899 76279
rect 39899 76245 39908 76279
rect 39856 76236 39908 76245
rect 46940 76304 46992 76356
rect 61016 76347 61068 76356
rect 61016 76313 61050 76347
rect 61050 76313 61068 76347
rect 61016 76304 61068 76313
rect 63132 76347 63184 76356
rect 63132 76313 63166 76347
rect 63166 76313 63184 76347
rect 63132 76304 63184 76313
rect 65984 76304 66036 76356
rect 67916 76347 67968 76356
rect 67916 76313 67950 76347
rect 67950 76313 67968 76347
rect 67916 76304 67968 76313
rect 69112 76347 69164 76356
rect 69112 76313 69121 76347
rect 69121 76313 69155 76347
rect 69155 76313 69164 76347
rect 69112 76304 69164 76313
rect 41328 76236 41380 76288
rect 42892 76279 42944 76288
rect 42892 76245 42901 76279
rect 42901 76245 42935 76279
rect 42935 76245 42944 76279
rect 42892 76236 42944 76245
rect 45468 76279 45520 76288
rect 45468 76245 45477 76279
rect 45477 76245 45511 76279
rect 45511 76245 45520 76279
rect 45468 76236 45520 76245
rect 62120 76279 62172 76288
rect 62120 76245 62129 76279
rect 62129 76245 62163 76279
rect 62163 76245 62172 76279
rect 62120 76236 62172 76245
rect 64236 76279 64288 76288
rect 64236 76245 64245 76279
rect 64245 76245 64279 76279
rect 64279 76245 64288 76279
rect 64236 76236 64288 76245
rect 74540 76236 74592 76288
rect 82544 76279 82596 76288
rect 82544 76245 82553 76279
rect 82553 76245 82587 76279
rect 82587 76245 82596 76279
rect 82544 76236 82596 76245
rect 83096 76279 83148 76288
rect 83096 76245 83105 76279
rect 83105 76245 83139 76279
rect 83139 76245 83148 76279
rect 83096 76236 83148 76245
rect 83464 76279 83516 76288
rect 83464 76245 83473 76279
rect 83473 76245 83507 76279
rect 83507 76245 83516 76279
rect 83464 76236 83516 76245
rect 83648 76279 83700 76288
rect 83648 76245 83657 76279
rect 83657 76245 83691 76279
rect 83691 76245 83700 76279
rect 83648 76236 83700 76245
rect 84844 76347 84896 76356
rect 84844 76313 84862 76347
rect 84862 76313 84896 76347
rect 84844 76304 84896 76313
rect 98460 76415 98512 76424
rect 98460 76381 98469 76415
rect 98469 76381 98503 76415
rect 98503 76381 98512 76415
rect 98460 76372 98512 76381
rect 98644 76415 98696 76424
rect 98644 76381 98653 76415
rect 98653 76381 98687 76415
rect 98687 76381 98696 76415
rect 98644 76372 98696 76381
rect 99012 76415 99064 76424
rect 99012 76381 99021 76415
rect 99021 76381 99055 76415
rect 99055 76381 99064 76415
rect 99012 76372 99064 76381
rect 93492 76304 93544 76356
rect 97724 76304 97776 76356
rect 98184 76304 98236 76356
rect 99196 76304 99248 76356
rect 100944 76440 100996 76492
rect 101036 76483 101088 76492
rect 101036 76449 101045 76483
rect 101045 76449 101079 76483
rect 101079 76449 101088 76483
rect 101036 76440 101088 76449
rect 100392 76372 100444 76424
rect 101128 76415 101180 76424
rect 101128 76381 101137 76415
rect 101137 76381 101171 76415
rect 101171 76381 101180 76415
rect 101128 76372 101180 76381
rect 92572 76279 92624 76288
rect 92572 76245 92581 76279
rect 92581 76245 92615 76279
rect 92615 76245 92624 76279
rect 92572 76236 92624 76245
rect 99564 76304 99616 76356
rect 100024 76236 100076 76288
rect 107936 76236 107988 76288
rect 108396 76279 108448 76288
rect 108396 76245 108405 76279
rect 108405 76245 108439 76279
rect 108439 76245 108448 76279
rect 108396 76236 108448 76245
rect 4874 76134 4926 76186
rect 4938 76134 4990 76186
rect 5002 76134 5054 76186
rect 5066 76134 5118 76186
rect 5130 76134 5182 76186
rect 35594 76134 35646 76186
rect 35658 76134 35710 76186
rect 35722 76134 35774 76186
rect 35786 76134 35838 76186
rect 35850 76134 35902 76186
rect 66314 76134 66366 76186
rect 66378 76134 66430 76186
rect 66442 76134 66494 76186
rect 66506 76134 66558 76186
rect 66570 76134 66622 76186
rect 97034 76134 97086 76186
rect 97098 76134 97150 76186
rect 97162 76134 97214 76186
rect 97226 76134 97278 76186
rect 97290 76134 97342 76186
rect 14648 76075 14700 76084
rect 14648 76041 14657 76075
rect 14657 76041 14691 76075
rect 14691 76041 14700 76075
rect 14648 76032 14700 76041
rect 16304 75964 16356 76016
rect 11060 75896 11112 75948
rect 14556 75896 14608 75948
rect 16580 76032 16632 76084
rect 22284 76032 22336 76084
rect 23572 76032 23624 76084
rect 30564 76032 30616 76084
rect 62120 76032 62172 76084
rect 68468 76032 68520 76084
rect 83648 76032 83700 76084
rect 84844 76032 84896 76084
rect 90456 76032 90508 76084
rect 93492 76032 93544 76084
rect 100576 76032 100628 76084
rect 100760 76075 100812 76084
rect 100760 76041 100769 76075
rect 100769 76041 100803 76075
rect 100803 76041 100812 76075
rect 100760 76032 100812 76041
rect 108396 76075 108448 76084
rect 108396 76041 108405 76075
rect 108405 76041 108439 76075
rect 108439 76041 108448 76075
rect 108396 76032 108448 76041
rect 64236 75964 64288 76016
rect 70124 75964 70176 76016
rect 90272 76007 90324 76016
rect 90272 75973 90281 76007
rect 90281 75973 90315 76007
rect 90315 75973 90324 76007
rect 90272 75964 90324 75973
rect 83464 75896 83516 75948
rect 93400 75964 93452 76016
rect 94044 75964 94096 76016
rect 98460 75964 98512 76016
rect 91192 75896 91244 75948
rect 96896 75896 96948 75948
rect 97724 75896 97776 75948
rect 18052 75828 18104 75880
rect 19340 75760 19392 75812
rect 88248 75760 88300 75812
rect 89720 75760 89772 75812
rect 1492 75735 1544 75744
rect 1492 75701 1501 75735
rect 1501 75701 1535 75735
rect 1535 75701 1544 75735
rect 1492 75692 1544 75701
rect 88064 75692 88116 75744
rect 89904 75735 89956 75744
rect 89904 75701 89913 75735
rect 89913 75701 89947 75735
rect 89947 75701 89956 75735
rect 89904 75692 89956 75701
rect 90088 75735 90140 75744
rect 90088 75701 90097 75735
rect 90097 75701 90131 75735
rect 90131 75701 90140 75735
rect 90088 75692 90140 75701
rect 92572 75692 92624 75744
rect 95424 75871 95476 75880
rect 95424 75837 95433 75871
rect 95433 75837 95467 75871
rect 95467 75837 95476 75871
rect 95424 75828 95476 75837
rect 98000 75828 98052 75880
rect 98552 75939 98604 75948
rect 98552 75905 98561 75939
rect 98561 75905 98595 75939
rect 98595 75905 98604 75939
rect 98552 75896 98604 75905
rect 98644 75939 98696 75948
rect 98644 75905 98653 75939
rect 98653 75905 98687 75939
rect 98687 75905 98696 75939
rect 98644 75896 98696 75905
rect 98736 75939 98788 75948
rect 98736 75905 98745 75939
rect 98745 75905 98779 75939
rect 98779 75905 98788 75939
rect 98736 75896 98788 75905
rect 99012 75896 99064 75948
rect 98460 75828 98512 75880
rect 98184 75760 98236 75812
rect 98644 75760 98696 75812
rect 99564 75896 99616 75948
rect 100024 75896 100076 75948
rect 100208 75828 100260 75880
rect 100392 75871 100444 75880
rect 100392 75837 100401 75871
rect 100401 75837 100435 75871
rect 100435 75837 100444 75871
rect 100392 75828 100444 75837
rect 101680 75828 101732 75880
rect 104072 75828 104124 75880
rect 100300 75760 100352 75812
rect 97540 75692 97592 75744
rect 98368 75735 98420 75744
rect 98368 75701 98377 75735
rect 98377 75701 98411 75735
rect 98411 75701 98420 75735
rect 98368 75692 98420 75701
rect 99104 75735 99156 75744
rect 99104 75701 99113 75735
rect 99113 75701 99147 75735
rect 99147 75701 99156 75735
rect 99104 75692 99156 75701
rect 99196 75692 99248 75744
rect 107936 75692 107988 75744
rect 4214 75590 4266 75642
rect 4278 75590 4330 75642
rect 4342 75590 4394 75642
rect 4406 75590 4458 75642
rect 4470 75590 4522 75642
rect 34934 75590 34986 75642
rect 34998 75590 35050 75642
rect 35062 75590 35114 75642
rect 35126 75590 35178 75642
rect 35190 75590 35242 75642
rect 65654 75590 65706 75642
rect 65718 75590 65770 75642
rect 65782 75590 65834 75642
rect 65846 75590 65898 75642
rect 65910 75590 65962 75642
rect 96374 75590 96426 75642
rect 96438 75590 96490 75642
rect 96502 75590 96554 75642
rect 96566 75590 96618 75642
rect 96630 75590 96682 75642
rect 22284 75531 22336 75540
rect 22284 75497 22293 75531
rect 22293 75497 22327 75531
rect 22327 75497 22336 75531
rect 22284 75488 22336 75497
rect 90272 75488 90324 75540
rect 91008 75488 91060 75540
rect 96804 75488 96856 75540
rect 98000 75488 98052 75540
rect 88248 75420 88300 75472
rect 97724 75420 97776 75472
rect 98644 75488 98696 75540
rect 99196 75488 99248 75540
rect 101680 75488 101732 75540
rect 99288 75420 99340 75472
rect 103520 75463 103572 75472
rect 103520 75429 103529 75463
rect 103529 75429 103563 75463
rect 103563 75429 103572 75463
rect 103520 75420 103572 75429
rect 18144 75284 18196 75336
rect 22376 75327 22428 75336
rect 22376 75293 22385 75327
rect 22385 75293 22419 75327
rect 22419 75293 22428 75327
rect 22376 75284 22428 75293
rect 19156 75216 19208 75268
rect 848 75148 900 75200
rect 22376 75148 22428 75200
rect 24768 75148 24820 75200
rect 86868 75284 86920 75336
rect 88156 75259 88208 75268
rect 88156 75225 88165 75259
rect 88165 75225 88199 75259
rect 88199 75225 88208 75259
rect 88156 75216 88208 75225
rect 87788 75148 87840 75200
rect 89628 75216 89680 75268
rect 90732 75259 90784 75268
rect 90732 75225 90741 75259
rect 90741 75225 90775 75259
rect 90775 75225 90784 75259
rect 90732 75216 90784 75225
rect 89904 75148 89956 75200
rect 93400 75395 93452 75404
rect 93400 75361 93409 75395
rect 93409 75361 93443 75395
rect 93443 75361 93452 75395
rect 93400 75352 93452 75361
rect 96896 75352 96948 75404
rect 91468 75216 91520 75268
rect 92388 75216 92440 75268
rect 91376 75148 91428 75200
rect 92572 75148 92624 75200
rect 98276 75327 98328 75336
rect 98276 75293 98285 75327
rect 98285 75293 98319 75327
rect 98319 75293 98328 75327
rect 98276 75284 98328 75293
rect 98368 75327 98420 75336
rect 98368 75293 98377 75327
rect 98377 75293 98411 75327
rect 98411 75293 98420 75327
rect 98368 75284 98420 75293
rect 100944 75352 100996 75404
rect 101404 75352 101456 75404
rect 101956 75395 102008 75404
rect 101956 75361 101965 75395
rect 101965 75361 101999 75395
rect 101999 75361 102008 75395
rect 101956 75352 102008 75361
rect 93032 75216 93084 75268
rect 96804 75148 96856 75200
rect 97908 75216 97960 75268
rect 98736 75216 98788 75268
rect 99380 75284 99432 75336
rect 100024 75284 100076 75336
rect 103152 75352 103204 75404
rect 103336 75352 103388 75404
rect 99472 75216 99524 75268
rect 99932 75216 99984 75268
rect 100392 75216 100444 75268
rect 102968 75327 103020 75336
rect 102968 75293 102977 75327
rect 102977 75293 103011 75327
rect 103011 75293 103020 75327
rect 102968 75284 103020 75293
rect 97448 75191 97500 75200
rect 97448 75157 97457 75191
rect 97457 75157 97491 75191
rect 97491 75157 97500 75191
rect 97448 75148 97500 75157
rect 98000 75148 98052 75200
rect 98184 75148 98236 75200
rect 100300 75148 100352 75200
rect 100484 75191 100536 75200
rect 100484 75157 100493 75191
rect 100493 75157 100527 75191
rect 100527 75157 100536 75191
rect 100484 75148 100536 75157
rect 101220 75191 101272 75200
rect 101220 75157 101229 75191
rect 101229 75157 101263 75191
rect 101263 75157 101272 75191
rect 101220 75148 101272 75157
rect 101956 75216 102008 75268
rect 102876 75216 102928 75268
rect 103060 75191 103112 75200
rect 103060 75157 103069 75191
rect 103069 75157 103103 75191
rect 103103 75157 103112 75191
rect 103060 75148 103112 75157
rect 103336 75216 103388 75268
rect 104164 75488 104216 75540
rect 104808 75488 104860 75540
rect 103980 75420 104032 75472
rect 104164 75327 104216 75336
rect 104164 75293 104173 75327
rect 104173 75293 104207 75327
rect 104207 75293 104216 75327
rect 104164 75284 104216 75293
rect 104072 75216 104124 75268
rect 104348 75191 104400 75200
rect 104348 75157 104357 75191
rect 104357 75157 104391 75191
rect 104391 75157 104400 75191
rect 104348 75148 104400 75157
rect 104440 75191 104492 75200
rect 104440 75157 104449 75191
rect 104449 75157 104483 75191
rect 104483 75157 104492 75191
rect 104440 75148 104492 75157
rect 107752 75284 107804 75336
rect 105268 75191 105320 75200
rect 105268 75157 105277 75191
rect 105277 75157 105311 75191
rect 105311 75157 105320 75191
rect 105268 75148 105320 75157
rect 108396 75191 108448 75200
rect 108396 75157 108405 75191
rect 108405 75157 108439 75191
rect 108439 75157 108448 75191
rect 108396 75148 108448 75157
rect 4874 75046 4926 75098
rect 4938 75046 4990 75098
rect 5002 75046 5054 75098
rect 5066 75046 5118 75098
rect 5130 75046 5182 75098
rect 35594 75046 35646 75098
rect 35658 75046 35710 75098
rect 35722 75046 35774 75098
rect 35786 75046 35838 75098
rect 35850 75046 35902 75098
rect 66314 75046 66366 75098
rect 66378 75046 66430 75098
rect 66442 75046 66494 75098
rect 66506 75046 66558 75098
rect 66570 75046 66622 75098
rect 97034 75046 97086 75098
rect 97098 75046 97150 75098
rect 97162 75046 97214 75098
rect 97226 75046 97278 75098
rect 97290 75046 97342 75098
rect 18052 74987 18104 74996
rect 18052 74953 18061 74987
rect 18061 74953 18095 74987
rect 18095 74953 18104 74987
rect 18052 74944 18104 74953
rect 18972 74944 19024 74996
rect 19892 74944 19944 74996
rect 86868 74944 86920 74996
rect 19156 74876 19208 74928
rect 85672 74876 85724 74928
rect 87788 74919 87840 74928
rect 87788 74885 87797 74919
rect 87797 74885 87831 74919
rect 87831 74885 87840 74919
rect 87788 74876 87840 74885
rect 88156 74944 88208 74996
rect 88708 74944 88760 74996
rect 89628 74987 89680 74996
rect 89628 74953 89637 74987
rect 89637 74953 89671 74987
rect 89671 74953 89680 74987
rect 89628 74944 89680 74953
rect 89720 74944 89772 74996
rect 91836 74944 91888 74996
rect 93308 74944 93360 74996
rect 88340 74919 88392 74928
rect 19892 74851 19944 74860
rect 19892 74817 19901 74851
rect 19901 74817 19935 74851
rect 19935 74817 19944 74851
rect 19892 74808 19944 74817
rect 88340 74885 88349 74919
rect 88349 74885 88383 74919
rect 88383 74885 88392 74919
rect 88340 74876 88392 74885
rect 93952 74876 94004 74928
rect 18144 74783 18196 74792
rect 18144 74749 18153 74783
rect 18153 74749 18187 74783
rect 18187 74749 18196 74783
rect 18144 74740 18196 74749
rect 28540 74740 28592 74792
rect 88156 74740 88208 74792
rect 85948 74604 86000 74656
rect 91468 74851 91520 74860
rect 91468 74817 91477 74851
rect 91477 74817 91511 74851
rect 91511 74817 91520 74851
rect 91468 74808 91520 74817
rect 89904 74740 89956 74792
rect 90732 74740 90784 74792
rect 91836 74851 91888 74860
rect 91836 74817 91845 74851
rect 91845 74817 91879 74851
rect 91879 74817 91888 74851
rect 91836 74808 91888 74817
rect 92388 74851 92440 74860
rect 92388 74817 92397 74851
rect 92397 74817 92431 74851
rect 92431 74817 92440 74851
rect 92388 74808 92440 74817
rect 94044 74808 94096 74860
rect 96896 74944 96948 74996
rect 97448 74944 97500 74996
rect 97908 74944 97960 74996
rect 97356 74851 97408 74860
rect 97356 74817 97365 74851
rect 97365 74817 97399 74851
rect 97399 74817 97408 74851
rect 97356 74808 97408 74817
rect 96712 74783 96764 74792
rect 96712 74749 96721 74783
rect 96721 74749 96755 74783
rect 96755 74749 96764 74783
rect 96712 74740 96764 74749
rect 97540 74851 97592 74860
rect 97540 74817 97549 74851
rect 97549 74817 97583 74851
rect 97583 74817 97592 74851
rect 97540 74808 97592 74817
rect 97724 74851 97776 74860
rect 97724 74817 97733 74851
rect 97733 74817 97767 74851
rect 97767 74817 97776 74851
rect 97724 74808 97776 74817
rect 98552 74876 98604 74928
rect 98368 74808 98420 74860
rect 99104 74944 99156 74996
rect 99472 74876 99524 74928
rect 99288 74851 99340 74860
rect 99288 74817 99297 74851
rect 99297 74817 99331 74851
rect 99331 74817 99340 74851
rect 99288 74808 99340 74817
rect 100116 74944 100168 74996
rect 100944 74987 100996 74996
rect 100944 74953 100959 74987
rect 100959 74953 100993 74987
rect 100993 74953 100996 74987
rect 100944 74944 100996 74953
rect 101220 74944 101272 74996
rect 101864 74944 101916 74996
rect 99932 74851 99984 74860
rect 99932 74817 99941 74851
rect 99941 74817 99975 74851
rect 99975 74817 99984 74851
rect 99932 74808 99984 74817
rect 100024 74808 100076 74860
rect 100208 74851 100260 74860
rect 100208 74817 100217 74851
rect 100217 74817 100251 74851
rect 100251 74817 100260 74851
rect 100208 74808 100260 74817
rect 100300 74851 100352 74860
rect 100300 74817 100309 74851
rect 100309 74817 100343 74851
rect 100343 74817 100352 74851
rect 100300 74808 100352 74817
rect 100484 74851 100536 74860
rect 100484 74817 100493 74851
rect 100493 74817 100527 74851
rect 100527 74817 100536 74851
rect 100484 74808 100536 74817
rect 97908 74740 97960 74792
rect 88708 74672 88760 74724
rect 99196 74740 99248 74792
rect 99472 74783 99524 74792
rect 99472 74749 99481 74783
rect 99481 74749 99515 74783
rect 99515 74749 99524 74783
rect 99472 74740 99524 74749
rect 98460 74672 98512 74724
rect 99840 74740 99892 74792
rect 100668 74808 100720 74860
rect 101128 74851 101180 74860
rect 101128 74817 101137 74851
rect 101137 74817 101171 74851
rect 101171 74817 101180 74851
rect 101128 74808 101180 74817
rect 101404 74851 101456 74860
rect 101404 74817 101413 74851
rect 101413 74817 101447 74851
rect 101447 74817 101456 74851
rect 101404 74808 101456 74817
rect 101956 74851 102008 74860
rect 101956 74817 101965 74851
rect 101965 74817 101999 74851
rect 101999 74817 102008 74851
rect 101956 74808 102008 74817
rect 102048 74851 102100 74860
rect 102048 74817 102057 74851
rect 102057 74817 102091 74851
rect 102091 74817 102100 74851
rect 102048 74808 102100 74817
rect 104072 74987 104124 74996
rect 104072 74953 104081 74987
rect 104081 74953 104115 74987
rect 104115 74953 104124 74987
rect 104072 74944 104124 74953
rect 102968 74876 103020 74928
rect 100208 74672 100260 74724
rect 102508 74808 102560 74860
rect 102876 74740 102928 74792
rect 103428 74808 103480 74860
rect 103796 74876 103848 74928
rect 104440 74919 104492 74928
rect 104440 74885 104449 74919
rect 104449 74885 104483 74919
rect 104483 74885 104492 74919
rect 104440 74876 104492 74885
rect 103980 74808 104032 74860
rect 104072 74808 104124 74860
rect 104808 74808 104860 74860
rect 104624 74740 104676 74792
rect 104992 74740 105044 74792
rect 103704 74672 103756 74724
rect 104348 74672 104400 74724
rect 88984 74647 89036 74656
rect 88984 74613 88993 74647
rect 88993 74613 89027 74647
rect 89027 74613 89036 74647
rect 88984 74604 89036 74613
rect 91284 74647 91336 74656
rect 91284 74613 91293 74647
rect 91293 74613 91327 74647
rect 91327 74613 91336 74647
rect 91284 74604 91336 74613
rect 91468 74604 91520 74656
rect 94412 74604 94464 74656
rect 96896 74604 96948 74656
rect 97356 74604 97408 74656
rect 97816 74604 97868 74656
rect 97908 74604 97960 74656
rect 99656 74604 99708 74656
rect 100300 74604 100352 74656
rect 100760 74647 100812 74656
rect 100760 74613 100769 74647
rect 100769 74613 100803 74647
rect 100803 74613 100812 74647
rect 100760 74604 100812 74613
rect 103152 74604 103204 74656
rect 103428 74604 103480 74656
rect 103612 74647 103664 74656
rect 103612 74613 103621 74647
rect 103621 74613 103655 74647
rect 103655 74613 103664 74647
rect 103612 74604 103664 74613
rect 103980 74604 104032 74656
rect 105360 74604 105412 74656
rect 4214 74502 4266 74554
rect 4278 74502 4330 74554
rect 4342 74502 4394 74554
rect 4406 74502 4458 74554
rect 4470 74502 4522 74554
rect 34934 74502 34986 74554
rect 34998 74502 35050 74554
rect 35062 74502 35114 74554
rect 35126 74502 35178 74554
rect 35190 74502 35242 74554
rect 65654 74502 65706 74554
rect 65718 74502 65770 74554
rect 65782 74502 65834 74554
rect 65846 74502 65898 74554
rect 65910 74502 65962 74554
rect 96374 74502 96426 74554
rect 96438 74502 96490 74554
rect 96502 74502 96554 74554
rect 96566 74502 96618 74554
rect 96630 74502 96682 74554
rect 35440 74400 35492 74452
rect 75092 74443 75144 74452
rect 75092 74409 75101 74443
rect 75101 74409 75135 74443
rect 75135 74409 75144 74443
rect 75092 74400 75144 74409
rect 82544 74400 82596 74452
rect 85672 74443 85724 74452
rect 85672 74409 85681 74443
rect 85681 74409 85715 74443
rect 85715 74409 85724 74443
rect 85672 74400 85724 74409
rect 85948 74443 86000 74452
rect 85948 74409 85957 74443
rect 85957 74409 85991 74443
rect 85991 74409 86000 74443
rect 85948 74400 86000 74409
rect 87144 74400 87196 74452
rect 88156 74400 88208 74452
rect 91192 74400 91244 74452
rect 93032 74400 93084 74452
rect 96712 74443 96764 74452
rect 96712 74409 96721 74443
rect 96721 74409 96755 74443
rect 96755 74409 96764 74443
rect 96712 74400 96764 74409
rect 98368 74400 98420 74452
rect 99288 74400 99340 74452
rect 101956 74400 102008 74452
rect 103428 74400 103480 74452
rect 848 74332 900 74384
rect 84292 74332 84344 74384
rect 88340 74307 88392 74316
rect 88340 74273 88349 74307
rect 88349 74273 88383 74307
rect 88383 74273 88392 74307
rect 88340 74264 88392 74273
rect 98644 74332 98696 74384
rect 100392 74375 100444 74384
rect 100392 74341 100401 74375
rect 100401 74341 100435 74375
rect 100435 74341 100444 74375
rect 100392 74332 100444 74341
rect 102048 74332 102100 74384
rect 102140 74332 102192 74384
rect 104164 74332 104216 74384
rect 104532 74332 104584 74384
rect 96804 74264 96856 74316
rect 98000 74264 98052 74316
rect 23388 74128 23440 74180
rect 24768 74239 24820 74248
rect 24768 74205 24777 74239
rect 24777 74205 24811 74239
rect 24811 74205 24820 74239
rect 28264 74239 28316 74248
rect 24768 74196 24820 74205
rect 28264 74205 28273 74239
rect 28273 74205 28307 74239
rect 28307 74205 28316 74239
rect 28264 74196 28316 74205
rect 25044 74128 25096 74180
rect 29644 74103 29696 74112
rect 29644 74069 29653 74103
rect 29653 74069 29687 74103
rect 29687 74069 29696 74103
rect 29644 74060 29696 74069
rect 74172 74196 74224 74248
rect 78772 74196 78824 74248
rect 85120 74196 85172 74248
rect 85948 74196 86000 74248
rect 87144 74239 87196 74248
rect 87144 74205 87153 74239
rect 87153 74205 87187 74239
rect 87187 74205 87196 74239
rect 87144 74196 87196 74205
rect 91192 74196 91244 74248
rect 97448 74196 97500 74248
rect 97908 74239 97960 74248
rect 97908 74205 97912 74239
rect 97912 74205 97946 74239
rect 97946 74205 97960 74239
rect 97908 74196 97960 74205
rect 99932 74264 99984 74316
rect 98276 74239 98328 74248
rect 98276 74205 98284 74239
rect 98284 74205 98318 74239
rect 98318 74205 98328 74239
rect 98276 74196 98328 74205
rect 98644 74196 98696 74248
rect 100208 74239 100260 74248
rect 100208 74205 100217 74239
rect 100217 74205 100251 74239
rect 100251 74205 100260 74239
rect 100208 74196 100260 74205
rect 100760 74264 100812 74316
rect 101864 74264 101916 74316
rect 103060 74264 103112 74316
rect 100576 74239 100628 74248
rect 100576 74205 100585 74239
rect 100585 74205 100619 74239
rect 100619 74205 100628 74239
rect 100576 74196 100628 74205
rect 101312 74239 101364 74248
rect 101312 74205 101321 74239
rect 101321 74205 101355 74239
rect 101355 74205 101364 74239
rect 101312 74196 101364 74205
rect 101680 74196 101732 74248
rect 103520 74264 103572 74316
rect 105360 74307 105412 74316
rect 105360 74273 105369 74307
rect 105369 74273 105403 74307
rect 105403 74273 105412 74307
rect 105360 74264 105412 74273
rect 105452 74307 105504 74316
rect 105452 74273 105461 74307
rect 105461 74273 105495 74307
rect 105495 74273 105504 74307
rect 105452 74264 105504 74273
rect 103244 74239 103296 74248
rect 103244 74205 103253 74239
rect 103253 74205 103287 74239
rect 103287 74205 103296 74239
rect 103244 74196 103296 74205
rect 104440 74239 104492 74248
rect 104440 74205 104449 74239
rect 104449 74205 104483 74239
rect 104483 74205 104492 74239
rect 104440 74196 104492 74205
rect 104900 74196 104952 74248
rect 105268 74239 105320 74248
rect 105268 74205 105277 74239
rect 105277 74205 105311 74239
rect 105311 74205 105320 74239
rect 105268 74196 105320 74205
rect 36176 74060 36228 74112
rect 88800 74060 88852 74112
rect 91376 74060 91428 74112
rect 97724 74103 97776 74112
rect 97724 74069 97733 74103
rect 97733 74069 97767 74103
rect 97767 74069 97776 74103
rect 97724 74060 97776 74069
rect 99196 74128 99248 74180
rect 99748 74128 99800 74180
rect 98920 74060 98972 74112
rect 99932 74060 99984 74112
rect 101588 74060 101640 74112
rect 101956 74060 102008 74112
rect 102876 74060 102928 74112
rect 104348 74128 104400 74180
rect 104992 74060 105044 74112
rect 108396 74103 108448 74112
rect 108396 74069 108405 74103
rect 108405 74069 108439 74103
rect 108439 74069 108448 74103
rect 108396 74060 108448 74069
rect 4874 73958 4926 74010
rect 4938 73958 4990 74010
rect 5002 73958 5054 74010
rect 5066 73958 5118 74010
rect 5130 73958 5182 74010
rect 35594 73958 35646 74010
rect 35658 73958 35710 74010
rect 35722 73958 35774 74010
rect 35786 73958 35838 74010
rect 35850 73958 35902 74010
rect 66314 73958 66366 74010
rect 66378 73958 66430 74010
rect 66442 73958 66494 74010
rect 66506 73958 66558 74010
rect 66570 73958 66622 74010
rect 97034 73958 97086 74010
rect 97098 73958 97150 74010
rect 97162 73958 97214 74010
rect 97226 73958 97278 74010
rect 97290 73958 97342 74010
rect 9588 73856 9640 73908
rect 23388 73788 23440 73840
rect 29644 73788 29696 73840
rect 39856 73856 39908 73908
rect 68468 73899 68520 73908
rect 68468 73865 68477 73899
rect 68477 73865 68511 73899
rect 68511 73865 68520 73899
rect 68468 73856 68520 73865
rect 70124 73899 70176 73908
rect 70124 73865 70133 73899
rect 70133 73865 70167 73899
rect 70167 73865 70176 73899
rect 70124 73856 70176 73865
rect 74540 73856 74592 73908
rect 75092 73899 75144 73908
rect 848 73584 900 73636
rect 1860 73559 1912 73568
rect 1860 73525 1869 73559
rect 1869 73525 1903 73559
rect 1903 73525 1912 73559
rect 1860 73516 1912 73525
rect 6184 73516 6236 73568
rect 18972 73763 19024 73772
rect 18972 73729 18981 73763
rect 18981 73729 19015 73763
rect 19015 73729 19024 73763
rect 18972 73720 19024 73729
rect 28264 73720 28316 73772
rect 38844 73720 38896 73772
rect 74724 73788 74776 73840
rect 68560 73763 68612 73772
rect 68560 73729 68569 73763
rect 68569 73729 68603 73763
rect 68603 73729 68612 73763
rect 68560 73720 68612 73729
rect 69020 73720 69072 73772
rect 74172 73720 74224 73772
rect 74540 73763 74592 73772
rect 74540 73729 74549 73763
rect 74549 73729 74583 73763
rect 74583 73729 74592 73763
rect 74540 73720 74592 73729
rect 11704 73652 11756 73704
rect 24676 73652 24728 73704
rect 24768 73695 24820 73704
rect 24768 73661 24777 73695
rect 24777 73661 24811 73695
rect 24811 73661 24820 73695
rect 24768 73652 24820 73661
rect 25044 73695 25096 73704
rect 25044 73661 25053 73695
rect 25053 73661 25087 73695
rect 25087 73661 25096 73695
rect 25044 73652 25096 73661
rect 31760 73652 31812 73704
rect 33048 73652 33100 73704
rect 37924 73652 37976 73704
rect 68284 73695 68336 73704
rect 68284 73661 68293 73695
rect 68293 73661 68327 73695
rect 68327 73661 68336 73695
rect 68284 73652 68336 73661
rect 72424 73652 72476 73704
rect 75092 73865 75101 73899
rect 75101 73865 75135 73899
rect 75135 73865 75144 73899
rect 75092 73856 75144 73865
rect 74908 73788 74960 73840
rect 88708 73856 88760 73908
rect 13820 73584 13872 73636
rect 18972 73516 19024 73568
rect 22928 73516 22980 73568
rect 27896 73559 27948 73568
rect 27896 73525 27905 73559
rect 27905 73525 27939 73559
rect 27939 73525 27948 73559
rect 27896 73516 27948 73525
rect 29368 73516 29420 73568
rect 56140 73516 56192 73568
rect 73160 73584 73212 73636
rect 73804 73584 73856 73636
rect 84292 73720 84344 73772
rect 85120 73763 85172 73772
rect 85120 73729 85129 73763
rect 85129 73729 85163 73763
rect 85163 73729 85172 73763
rect 85120 73720 85172 73729
rect 91376 73856 91428 73908
rect 93308 73899 93360 73908
rect 93308 73865 93317 73899
rect 93317 73865 93351 73899
rect 93351 73865 93360 73899
rect 93308 73856 93360 73865
rect 89536 73788 89588 73840
rect 91008 73831 91060 73840
rect 91008 73797 91017 73831
rect 91017 73797 91051 73831
rect 91051 73797 91060 73831
rect 91008 73788 91060 73797
rect 98184 73856 98236 73908
rect 98828 73899 98880 73908
rect 98828 73865 98837 73899
rect 98837 73865 98871 73899
rect 98871 73865 98880 73899
rect 98828 73856 98880 73865
rect 98920 73856 98972 73908
rect 99748 73856 99800 73908
rect 99932 73856 99984 73908
rect 100300 73856 100352 73908
rect 91284 73720 91336 73772
rect 78588 73652 78640 73704
rect 85580 73652 85632 73704
rect 70584 73559 70636 73568
rect 70584 73525 70593 73559
rect 70593 73525 70627 73559
rect 70627 73525 70636 73559
rect 70584 73516 70636 73525
rect 89076 73695 89128 73704
rect 89076 73661 89085 73695
rect 89085 73661 89119 73695
rect 89119 73661 89128 73695
rect 89076 73652 89128 73661
rect 97816 73788 97868 73840
rect 98276 73788 98328 73840
rect 93308 73720 93360 73772
rect 86040 73516 86092 73568
rect 89628 73516 89680 73568
rect 91468 73584 91520 73636
rect 93860 73720 93912 73772
rect 94412 73763 94464 73772
rect 94412 73729 94421 73763
rect 94421 73729 94455 73763
rect 94455 73729 94464 73763
rect 94412 73720 94464 73729
rect 97448 73720 97500 73772
rect 98460 73720 98512 73772
rect 99012 73720 99064 73772
rect 98368 73652 98420 73704
rect 99288 73763 99340 73772
rect 99288 73729 99297 73763
rect 99297 73729 99331 73763
rect 99331 73729 99340 73763
rect 99288 73720 99340 73729
rect 99380 73720 99432 73772
rect 100576 73788 100628 73840
rect 101128 73788 101180 73840
rect 102140 73856 102192 73908
rect 103428 73856 103480 73908
rect 104440 73856 104492 73908
rect 105452 73856 105504 73908
rect 101588 73788 101640 73840
rect 102876 73788 102928 73840
rect 100484 73763 100536 73772
rect 100484 73729 100493 73763
rect 100493 73729 100527 73763
rect 100527 73729 100536 73763
rect 100484 73720 100536 73729
rect 100760 73720 100812 73772
rect 101772 73720 101824 73772
rect 98644 73627 98696 73636
rect 98644 73593 98653 73627
rect 98653 73593 98687 73627
rect 98687 73593 98696 73627
rect 98644 73584 98696 73593
rect 98736 73584 98788 73636
rect 99656 73652 99708 73704
rect 99472 73627 99524 73636
rect 99472 73593 99481 73627
rect 99481 73593 99515 73627
rect 99515 73593 99524 73627
rect 99472 73584 99524 73593
rect 100300 73695 100352 73704
rect 100300 73661 100309 73695
rect 100309 73661 100343 73695
rect 100343 73661 100352 73695
rect 100300 73652 100352 73661
rect 100392 73695 100444 73704
rect 100392 73661 100401 73695
rect 100401 73661 100435 73695
rect 100435 73661 100444 73695
rect 100392 73652 100444 73661
rect 101312 73584 101364 73636
rect 91376 73559 91428 73568
rect 91376 73525 91385 73559
rect 91385 73525 91419 73559
rect 91419 73525 91428 73559
rect 91376 73516 91428 73525
rect 91836 73516 91888 73568
rect 93584 73559 93636 73568
rect 93584 73525 93593 73559
rect 93593 73525 93627 73559
rect 93627 73525 93636 73559
rect 93584 73516 93636 73525
rect 93952 73559 94004 73568
rect 93952 73525 93961 73559
rect 93961 73525 93995 73559
rect 93995 73525 94004 73559
rect 93952 73516 94004 73525
rect 100116 73516 100168 73568
rect 100300 73516 100352 73568
rect 102784 73720 102836 73772
rect 103060 73720 103112 73772
rect 103520 73788 103572 73840
rect 104624 73831 104676 73840
rect 104624 73797 104633 73831
rect 104633 73797 104667 73831
rect 104667 73797 104676 73831
rect 104624 73788 104676 73797
rect 105912 73856 105964 73908
rect 103428 73763 103480 73772
rect 103428 73729 103437 73763
rect 103437 73729 103471 73763
rect 103471 73729 103480 73763
rect 103428 73720 103480 73729
rect 103612 73652 103664 73704
rect 103796 73584 103848 73636
rect 104716 73763 104768 73772
rect 104716 73729 104730 73763
rect 104730 73729 104764 73763
rect 104764 73729 104768 73763
rect 104716 73720 104768 73729
rect 105176 73763 105228 73772
rect 105176 73729 105185 73763
rect 105185 73729 105219 73763
rect 105219 73729 105228 73763
rect 105176 73720 105228 73729
rect 105360 73763 105412 73772
rect 105360 73729 105369 73763
rect 105369 73729 105403 73763
rect 105403 73729 105412 73763
rect 105360 73720 105412 73729
rect 105544 73720 105596 73772
rect 108488 73763 108540 73772
rect 108488 73729 108497 73763
rect 108497 73729 108531 73763
rect 108531 73729 108540 73763
rect 108488 73720 108540 73729
rect 104900 73652 104952 73704
rect 104624 73584 104676 73636
rect 105268 73584 105320 73636
rect 103520 73516 103572 73568
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 34934 73414 34986 73466
rect 34998 73414 35050 73466
rect 35062 73414 35114 73466
rect 35126 73414 35178 73466
rect 35190 73414 35242 73466
rect 65654 73414 65706 73466
rect 65718 73414 65770 73466
rect 65782 73414 65834 73466
rect 65846 73414 65898 73466
rect 65910 73414 65962 73466
rect 96374 73414 96426 73466
rect 96438 73414 96490 73466
rect 96502 73414 96554 73466
rect 96566 73414 96618 73466
rect 96630 73414 96682 73466
rect 1860 73312 1912 73364
rect 22928 73176 22980 73228
rect 25044 73312 25096 73364
rect 70584 73312 70636 73364
rect 78588 73312 78640 73364
rect 69112 73244 69164 73296
rect 848 72972 900 73024
rect 29368 73176 29420 73228
rect 37924 73219 37976 73228
rect 37924 73185 37933 73219
rect 37933 73185 37967 73219
rect 37967 73185 37976 73219
rect 37924 73176 37976 73185
rect 68284 73176 68336 73228
rect 72424 73219 72476 73228
rect 72424 73185 72433 73219
rect 72433 73185 72467 73219
rect 72467 73185 72476 73219
rect 72424 73176 72476 73185
rect 24768 73108 24820 73160
rect 27896 72972 27948 73024
rect 35440 72972 35492 73024
rect 37740 73015 37792 73024
rect 37740 72981 37749 73015
rect 37749 72981 37783 73015
rect 37783 72981 37792 73015
rect 37740 72972 37792 72981
rect 37832 73015 37884 73024
rect 37832 72981 37841 73015
rect 37841 72981 37875 73015
rect 37875 72981 37884 73015
rect 37832 72972 37884 72981
rect 45468 73108 45520 73160
rect 68928 73108 68980 73160
rect 72884 73176 72936 73228
rect 78772 73287 78824 73296
rect 78772 73253 78781 73287
rect 78781 73253 78815 73287
rect 78815 73253 78824 73287
rect 78772 73244 78824 73253
rect 88156 73355 88208 73364
rect 88156 73321 88165 73355
rect 88165 73321 88199 73355
rect 88199 73321 88208 73355
rect 88156 73312 88208 73321
rect 93308 73312 93360 73364
rect 98552 73355 98604 73364
rect 98552 73321 98561 73355
rect 98561 73321 98595 73355
rect 98595 73321 98604 73355
rect 98552 73312 98604 73321
rect 99288 73312 99340 73364
rect 99564 73355 99616 73364
rect 99564 73321 99573 73355
rect 99573 73321 99607 73355
rect 99607 73321 99616 73355
rect 99564 73312 99616 73321
rect 100300 73312 100352 73364
rect 100392 73312 100444 73364
rect 93860 73176 93912 73228
rect 97724 73244 97776 73296
rect 98460 73244 98512 73296
rect 100116 73244 100168 73296
rect 101864 73312 101916 73364
rect 89536 73108 89588 73160
rect 96896 73108 96948 73160
rect 99932 73176 99984 73228
rect 101588 73244 101640 73296
rect 101772 73244 101824 73296
rect 103336 73355 103388 73364
rect 103336 73321 103345 73355
rect 103345 73321 103379 73355
rect 103379 73321 103388 73355
rect 103336 73312 103388 73321
rect 103152 73244 103204 73296
rect 104624 73312 104676 73364
rect 103980 73244 104032 73296
rect 105452 73244 105504 73296
rect 70216 73083 70268 73092
rect 70216 73049 70225 73083
rect 70225 73049 70259 73083
rect 70259 73049 70268 73083
rect 70216 73040 70268 73049
rect 70400 73040 70452 73092
rect 81992 73040 82044 73092
rect 97540 73108 97592 73160
rect 97724 73151 97776 73160
rect 97724 73117 97733 73151
rect 97733 73117 97767 73151
rect 97767 73117 97776 73151
rect 97724 73108 97776 73117
rect 98092 73151 98144 73160
rect 98092 73117 98101 73151
rect 98101 73117 98135 73151
rect 98135 73117 98144 73151
rect 98092 73108 98144 73117
rect 98184 73151 98236 73160
rect 98184 73117 98193 73151
rect 98193 73117 98227 73151
rect 98227 73117 98236 73151
rect 98184 73108 98236 73117
rect 42708 72972 42760 73024
rect 69112 72972 69164 73024
rect 73068 73015 73120 73024
rect 73068 72981 73077 73015
rect 73077 72981 73111 73015
rect 73111 72981 73120 73015
rect 73068 72972 73120 72981
rect 96160 72972 96212 73024
rect 97448 73015 97500 73024
rect 97448 72981 97457 73015
rect 97457 72981 97491 73015
rect 97491 72981 97500 73015
rect 97448 72972 97500 72981
rect 97540 72972 97592 73024
rect 97908 73040 97960 73092
rect 98276 72972 98328 73024
rect 99656 73108 99708 73160
rect 100208 73108 100260 73160
rect 100668 73108 100720 73160
rect 101864 73176 101916 73228
rect 102784 73219 102836 73228
rect 102784 73185 102793 73219
rect 102793 73185 102827 73219
rect 102827 73185 102836 73219
rect 102784 73176 102836 73185
rect 103796 73176 103848 73228
rect 104440 73176 104492 73228
rect 103244 73108 103296 73160
rect 99196 73015 99248 73024
rect 99196 72981 99205 73015
rect 99205 72981 99239 73015
rect 99239 72981 99248 73015
rect 99196 72972 99248 72981
rect 100484 72972 100536 73024
rect 101220 73083 101272 73092
rect 101220 73049 101229 73083
rect 101229 73049 101263 73083
rect 101263 73049 101272 73083
rect 101220 73040 101272 73049
rect 102508 73083 102560 73092
rect 102508 73049 102517 73083
rect 102517 73049 102551 73083
rect 102551 73049 102560 73083
rect 102508 73040 102560 73049
rect 104624 73108 104676 73160
rect 105636 73151 105688 73160
rect 105636 73117 105645 73151
rect 105645 73117 105679 73151
rect 105679 73117 105688 73151
rect 105636 73108 105688 73117
rect 101496 72972 101548 73024
rect 101772 72972 101824 73024
rect 108120 73108 108172 73160
rect 108488 73151 108540 73160
rect 108488 73117 108497 73151
rect 108497 73117 108531 73151
rect 108531 73117 108540 73151
rect 108488 73108 108540 73117
rect 104256 73015 104308 73024
rect 104256 72981 104265 73015
rect 104265 72981 104299 73015
rect 104299 72981 104308 73015
rect 104256 72972 104308 72981
rect 105268 72972 105320 73024
rect 105636 72972 105688 73024
rect 4874 72870 4926 72922
rect 4938 72870 4990 72922
rect 5002 72870 5054 72922
rect 5066 72870 5118 72922
rect 5130 72870 5182 72922
rect 35594 72870 35646 72922
rect 35658 72870 35710 72922
rect 35722 72870 35774 72922
rect 35786 72870 35838 72922
rect 35850 72870 35902 72922
rect 66314 72870 66366 72922
rect 66378 72870 66430 72922
rect 66442 72870 66494 72922
rect 66506 72870 66558 72922
rect 66570 72870 66622 72922
rect 97034 72870 97086 72922
rect 97098 72870 97150 72922
rect 97162 72870 97214 72922
rect 97226 72870 97278 72922
rect 97290 72870 97342 72922
rect 37832 72768 37884 72820
rect 42892 72768 42944 72820
rect 69112 72811 69164 72820
rect 37740 72700 37792 72752
rect 42432 72700 42484 72752
rect 11704 72632 11756 72684
rect 69112 72777 69121 72811
rect 69121 72777 69155 72811
rect 69155 72777 69164 72811
rect 69112 72768 69164 72777
rect 73068 72768 73120 72820
rect 85580 72768 85632 72820
rect 86684 72768 86736 72820
rect 85488 72700 85540 72752
rect 97908 72768 97960 72820
rect 98184 72768 98236 72820
rect 100024 72811 100076 72820
rect 100024 72777 100033 72811
rect 100033 72777 100067 72811
rect 100067 72777 100076 72811
rect 100024 72768 100076 72777
rect 100852 72811 100904 72820
rect 100852 72777 100861 72811
rect 100861 72777 100895 72811
rect 100895 72777 100904 72811
rect 100852 72768 100904 72777
rect 101220 72768 101272 72820
rect 103796 72768 103848 72820
rect 104624 72768 104676 72820
rect 105176 72768 105228 72820
rect 105360 72811 105412 72820
rect 105360 72777 105369 72811
rect 105369 72777 105403 72811
rect 105403 72777 105412 72811
rect 105360 72768 105412 72777
rect 105452 72768 105504 72820
rect 106004 72768 106056 72820
rect 94504 72700 94556 72752
rect 96068 72700 96120 72752
rect 97632 72743 97684 72752
rect 97632 72709 97641 72743
rect 97641 72709 97675 72743
rect 97675 72709 97684 72743
rect 97632 72700 97684 72709
rect 848 72428 900 72480
rect 86040 72471 86092 72480
rect 86040 72437 86049 72471
rect 86049 72437 86083 72471
rect 86083 72437 86092 72471
rect 86040 72428 86092 72437
rect 97724 72632 97776 72684
rect 98460 72700 98512 72752
rect 86224 72564 86276 72616
rect 86684 72607 86736 72616
rect 86684 72573 86693 72607
rect 86693 72573 86727 72607
rect 86727 72573 86736 72607
rect 86684 72564 86736 72573
rect 98368 72632 98420 72684
rect 98736 72675 98788 72684
rect 98736 72641 98745 72675
rect 98745 72641 98779 72675
rect 98779 72641 98788 72675
rect 98736 72632 98788 72641
rect 100392 72675 100444 72684
rect 100392 72641 100401 72675
rect 100401 72641 100435 72675
rect 100435 72641 100444 72675
rect 100392 72632 100444 72641
rect 89076 72428 89128 72480
rect 98092 72564 98144 72616
rect 98552 72564 98604 72616
rect 99564 72564 99616 72616
rect 100024 72564 100076 72616
rect 102784 72743 102836 72752
rect 102784 72709 102793 72743
rect 102793 72709 102827 72743
rect 102827 72709 102836 72743
rect 102784 72700 102836 72709
rect 100668 72632 100720 72684
rect 101128 72675 101180 72684
rect 101128 72641 101137 72675
rect 101137 72641 101171 72675
rect 101171 72641 101180 72675
rect 101128 72632 101180 72641
rect 101588 72675 101640 72684
rect 101588 72641 101597 72675
rect 101597 72641 101631 72675
rect 101631 72641 101640 72675
rect 101588 72632 101640 72641
rect 98276 72496 98328 72548
rect 97632 72428 97684 72480
rect 101496 72564 101548 72616
rect 101864 72675 101916 72684
rect 101864 72641 101873 72675
rect 101873 72641 101907 72675
rect 101907 72641 101916 72675
rect 101864 72632 101916 72641
rect 103612 72632 103664 72684
rect 104532 72700 104584 72752
rect 103796 72675 103848 72684
rect 103796 72641 103805 72675
rect 103805 72641 103839 72675
rect 103839 72641 103848 72675
rect 103796 72632 103848 72641
rect 103336 72564 103388 72616
rect 103428 72564 103480 72616
rect 104256 72564 104308 72616
rect 101312 72496 101364 72548
rect 103520 72496 103572 72548
rect 104808 72632 104860 72684
rect 104716 72564 104768 72616
rect 105452 72675 105504 72684
rect 105452 72641 105461 72675
rect 105461 72641 105495 72675
rect 105495 72641 105504 72675
rect 105452 72632 105504 72641
rect 105912 72675 105964 72684
rect 105912 72641 105921 72675
rect 105921 72641 105955 72675
rect 105955 72641 105964 72675
rect 105912 72632 105964 72641
rect 108488 72675 108540 72684
rect 108488 72641 108497 72675
rect 108497 72641 108531 72675
rect 108531 72641 108540 72675
rect 108488 72632 108540 72641
rect 103060 72428 103112 72480
rect 103152 72428 103204 72480
rect 103704 72428 103756 72480
rect 105176 72496 105228 72548
rect 105820 72471 105872 72480
rect 105820 72437 105829 72471
rect 105829 72437 105863 72471
rect 105863 72437 105872 72471
rect 105820 72428 105872 72437
rect 106004 72471 106056 72480
rect 106004 72437 106013 72471
rect 106013 72437 106047 72471
rect 106047 72437 106056 72471
rect 106004 72428 106056 72437
rect 106096 72428 106148 72480
rect 108304 72471 108356 72480
rect 108304 72437 108313 72471
rect 108313 72437 108347 72471
rect 108347 72437 108356 72471
rect 108304 72428 108356 72437
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 34934 72326 34986 72378
rect 34998 72326 35050 72378
rect 35062 72326 35114 72378
rect 35126 72326 35178 72378
rect 35190 72326 35242 72378
rect 65654 72326 65706 72378
rect 65718 72326 65770 72378
rect 65782 72326 65834 72378
rect 65846 72326 65898 72378
rect 65910 72326 65962 72378
rect 96374 72326 96426 72378
rect 96438 72326 96490 72378
rect 96502 72326 96554 72378
rect 96566 72326 96618 72378
rect 96630 72326 96682 72378
rect 81992 72267 82044 72276
rect 81992 72233 82001 72267
rect 82001 72233 82035 72267
rect 82035 72233 82044 72267
rect 81992 72224 82044 72233
rect 85488 72267 85540 72276
rect 85488 72233 85497 72267
rect 85497 72233 85531 72267
rect 85531 72233 85540 72267
rect 85488 72224 85540 72233
rect 88156 72224 88208 72276
rect 85120 72156 85172 72208
rect 85212 72088 85264 72140
rect 85396 72063 85448 72072
rect 85396 72029 85405 72063
rect 85405 72029 85439 72063
rect 85439 72029 85448 72063
rect 85396 72020 85448 72029
rect 89720 72224 89772 72276
rect 94504 72224 94556 72276
rect 93952 72156 94004 72208
rect 96804 72131 96856 72140
rect 96804 72097 96813 72131
rect 96813 72097 96847 72131
rect 96847 72097 96856 72131
rect 96804 72088 96856 72097
rect 97632 72156 97684 72208
rect 98460 72199 98512 72208
rect 98460 72165 98469 72199
rect 98469 72165 98503 72199
rect 98503 72165 98512 72199
rect 98460 72156 98512 72165
rect 99104 72224 99156 72276
rect 101772 72224 101824 72276
rect 103244 72224 103296 72276
rect 104716 72224 104768 72276
rect 104072 72156 104124 72208
rect 93584 72063 93636 72072
rect 93584 72029 93591 72063
rect 93591 72029 93636 72063
rect 93584 72020 93636 72029
rect 94320 72020 94372 72072
rect 96712 72063 96764 72072
rect 96712 72029 96721 72063
rect 96721 72029 96755 72063
rect 96755 72029 96764 72063
rect 96712 72020 96764 72029
rect 98736 72088 98788 72140
rect 98000 72020 98052 72072
rect 98092 72063 98144 72072
rect 98092 72029 98101 72063
rect 98101 72029 98135 72063
rect 98135 72029 98144 72063
rect 98092 72020 98144 72029
rect 90088 71952 90140 72004
rect 83464 71927 83516 71936
rect 83464 71893 83473 71927
rect 83473 71893 83507 71927
rect 83507 71893 83516 71927
rect 83464 71884 83516 71893
rect 93768 71995 93820 72004
rect 93768 71961 93777 71995
rect 93777 71961 93811 71995
rect 93811 71961 93820 71995
rect 93768 71952 93820 71961
rect 98552 72063 98604 72072
rect 98552 72029 98561 72063
rect 98561 72029 98595 72063
rect 98595 72029 98604 72063
rect 98552 72020 98604 72029
rect 100852 72088 100904 72140
rect 102324 72088 102376 72140
rect 103980 72088 104032 72140
rect 100024 72063 100076 72072
rect 100024 72029 100033 72063
rect 100033 72029 100067 72063
rect 100067 72029 100076 72063
rect 100024 72020 100076 72029
rect 93860 71884 93912 71936
rect 95056 71884 95108 71936
rect 98368 71952 98420 72004
rect 99196 71995 99248 72004
rect 99196 71961 99205 71995
rect 99205 71961 99239 71995
rect 99239 71961 99248 71995
rect 99196 71952 99248 71961
rect 99564 71952 99616 72004
rect 100300 72020 100352 72072
rect 101220 72020 101272 72072
rect 102508 72020 102560 72072
rect 103060 72063 103112 72072
rect 103060 72029 103069 72063
rect 103069 72029 103103 72063
rect 103103 72029 103112 72063
rect 103060 72020 103112 72029
rect 103152 72063 103204 72072
rect 103152 72029 103161 72063
rect 103161 72029 103195 72063
rect 103195 72029 103204 72063
rect 103152 72020 103204 72029
rect 103428 72063 103480 72072
rect 103428 72029 103437 72063
rect 103437 72029 103471 72063
rect 103471 72029 103480 72063
rect 103428 72020 103480 72029
rect 103520 72063 103572 72072
rect 103520 72029 103529 72063
rect 103529 72029 103563 72063
rect 103563 72029 103572 72063
rect 103520 72020 103572 72029
rect 107292 72156 107344 72208
rect 104532 72063 104584 72072
rect 104532 72029 104541 72063
rect 104541 72029 104575 72063
rect 104575 72029 104584 72063
rect 104532 72020 104584 72029
rect 106004 72088 106056 72140
rect 105268 72063 105320 72072
rect 105268 72029 105277 72063
rect 105277 72029 105311 72063
rect 105311 72029 105320 72063
rect 105268 72020 105320 72029
rect 105360 72020 105412 72072
rect 101404 71952 101456 72004
rect 103336 71952 103388 72004
rect 104900 71952 104952 72004
rect 98644 71884 98696 71936
rect 99012 71927 99064 71936
rect 99012 71893 99039 71927
rect 99039 71893 99064 71927
rect 99012 71884 99064 71893
rect 100576 71884 100628 71936
rect 102324 71927 102376 71936
rect 102324 71893 102333 71927
rect 102333 71893 102367 71927
rect 102367 71893 102376 71927
rect 102324 71884 102376 71893
rect 102784 71884 102836 71936
rect 103520 71884 103572 71936
rect 103796 71884 103848 71936
rect 104440 71884 104492 71936
rect 104808 71884 104860 71936
rect 105636 72063 105688 72072
rect 105636 72029 105645 72063
rect 105645 72029 105679 72063
rect 105679 72029 105688 72063
rect 105636 72020 105688 72029
rect 105820 72020 105872 72072
rect 106096 71952 106148 72004
rect 105544 71884 105596 71936
rect 105820 71927 105872 71936
rect 105820 71893 105829 71927
rect 105829 71893 105863 71927
rect 105863 71893 105872 71927
rect 105820 71884 105872 71893
rect 106004 71927 106056 71936
rect 106004 71893 106013 71927
rect 106013 71893 106047 71927
rect 106047 71893 106056 71927
rect 106004 71884 106056 71893
rect 4874 71782 4926 71834
rect 4938 71782 4990 71834
rect 5002 71782 5054 71834
rect 5066 71782 5118 71834
rect 5130 71782 5182 71834
rect 35594 71782 35646 71834
rect 35658 71782 35710 71834
rect 35722 71782 35774 71834
rect 35786 71782 35838 71834
rect 35850 71782 35902 71834
rect 66314 71782 66366 71834
rect 66378 71782 66430 71834
rect 66442 71782 66494 71834
rect 66506 71782 66558 71834
rect 66570 71782 66622 71834
rect 97034 71782 97086 71834
rect 97098 71782 97150 71834
rect 97162 71782 97214 71834
rect 97226 71782 97278 71834
rect 97290 71782 97342 71834
rect 89628 71655 89680 71664
rect 89628 71621 89637 71655
rect 89637 71621 89671 71655
rect 89671 71621 89680 71655
rect 89628 71612 89680 71621
rect 90088 71612 90140 71664
rect 92480 71680 92532 71732
rect 96804 71680 96856 71732
rect 98092 71680 98144 71732
rect 98920 71680 98972 71732
rect 100300 71680 100352 71732
rect 100392 71680 100444 71732
rect 101404 71723 101456 71732
rect 101404 71689 101413 71723
rect 101413 71689 101447 71723
rect 101447 71689 101456 71723
rect 101404 71680 101456 71689
rect 96160 71655 96212 71664
rect 96160 71621 96169 71655
rect 96169 71621 96203 71655
rect 96203 71621 96212 71655
rect 96160 71612 96212 71621
rect 98552 71655 98604 71664
rect 1216 71544 1268 71596
rect 98552 71621 98561 71655
rect 98561 71621 98595 71655
rect 98595 71621 98604 71655
rect 98552 71612 98604 71621
rect 97540 71544 97592 71596
rect 97908 71544 97960 71596
rect 98368 71544 98420 71596
rect 99196 71612 99248 71664
rect 104532 71680 104584 71732
rect 98092 71476 98144 71528
rect 99012 71476 99064 71528
rect 94320 71408 94372 71460
rect 23480 71340 23532 71392
rect 36176 71340 36228 71392
rect 84844 71340 84896 71392
rect 89168 71383 89220 71392
rect 89168 71349 89177 71383
rect 89177 71349 89211 71383
rect 89211 71349 89220 71383
rect 89168 71340 89220 71349
rect 95700 71383 95752 71392
rect 95700 71349 95709 71383
rect 95709 71349 95743 71383
rect 95743 71349 95752 71383
rect 95700 71340 95752 71349
rect 97448 71408 97500 71460
rect 97632 71408 97684 71460
rect 97908 71340 97960 71392
rect 98552 71408 98604 71460
rect 99104 71408 99156 71460
rect 99748 71587 99800 71596
rect 99748 71553 99757 71587
rect 99757 71553 99791 71587
rect 99791 71553 99800 71587
rect 99748 71544 99800 71553
rect 99840 71587 99892 71596
rect 99840 71553 99849 71587
rect 99849 71553 99883 71587
rect 99883 71553 99892 71587
rect 99840 71544 99892 71553
rect 100852 71587 100904 71596
rect 100852 71553 100861 71587
rect 100861 71553 100895 71587
rect 100895 71553 100904 71587
rect 100852 71544 100904 71553
rect 101772 71587 101824 71596
rect 101772 71553 101781 71587
rect 101781 71553 101815 71587
rect 101815 71553 101824 71587
rect 101772 71544 101824 71553
rect 102140 71544 102192 71596
rect 102784 71587 102836 71596
rect 102784 71553 102793 71587
rect 102793 71553 102827 71587
rect 102827 71553 102836 71587
rect 102784 71544 102836 71553
rect 103244 71544 103296 71596
rect 104900 71612 104952 71664
rect 100300 71476 100352 71528
rect 100576 71408 100628 71460
rect 98920 71383 98972 71392
rect 98920 71349 98929 71383
rect 98929 71349 98963 71383
rect 98963 71349 98972 71383
rect 98920 71340 98972 71349
rect 99380 71340 99432 71392
rect 100668 71340 100720 71392
rect 103428 71408 103480 71460
rect 103796 71587 103848 71596
rect 103796 71553 103805 71587
rect 103805 71553 103839 71587
rect 103839 71553 103848 71587
rect 103796 71544 103848 71553
rect 104440 71587 104492 71596
rect 104440 71553 104449 71587
rect 104449 71553 104483 71587
rect 104483 71553 104492 71587
rect 104440 71544 104492 71553
rect 104624 71544 104676 71596
rect 104716 71587 104768 71596
rect 104716 71553 104725 71587
rect 104725 71553 104759 71587
rect 104759 71553 104768 71587
rect 104716 71544 104768 71553
rect 104992 71544 105044 71596
rect 105360 71587 105412 71596
rect 105360 71553 105369 71587
rect 105369 71553 105403 71587
rect 105403 71553 105412 71587
rect 105360 71544 105412 71553
rect 105728 71544 105780 71596
rect 108304 71544 108356 71596
rect 108488 71587 108540 71596
rect 108488 71553 108497 71587
rect 108497 71553 108531 71587
rect 108531 71553 108540 71587
rect 108488 71544 108540 71553
rect 106004 71476 106056 71528
rect 104992 71408 105044 71460
rect 103888 71340 103940 71392
rect 104900 71340 104952 71392
rect 105360 71340 105412 71392
rect 106280 71340 106332 71392
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 34934 71238 34986 71290
rect 34998 71238 35050 71290
rect 35062 71238 35114 71290
rect 35126 71238 35178 71290
rect 35190 71238 35242 71290
rect 65654 71238 65706 71290
rect 65718 71238 65770 71290
rect 65782 71238 65834 71290
rect 65846 71238 65898 71290
rect 65910 71238 65962 71290
rect 96374 71238 96426 71290
rect 96438 71238 96490 71290
rect 96502 71238 96554 71290
rect 96566 71238 96618 71290
rect 96630 71238 96682 71290
rect 31760 71136 31812 71188
rect 5264 70864 5316 70916
rect 55128 71136 55180 71188
rect 84016 71136 84068 71188
rect 85212 71136 85264 71188
rect 86316 71179 86368 71188
rect 86316 71145 86325 71179
rect 86325 71145 86359 71179
rect 86359 71145 86368 71179
rect 86316 71136 86368 71145
rect 93308 71136 93360 71188
rect 85396 71068 85448 71120
rect 92480 71068 92532 71120
rect 96712 71136 96764 71188
rect 72884 71043 72936 71052
rect 72884 71009 72893 71043
rect 72893 71009 72927 71043
rect 72927 71009 72936 71043
rect 72884 71000 72936 71009
rect 86040 71000 86092 71052
rect 89168 71000 89220 71052
rect 93860 71000 93912 71052
rect 94872 71000 94924 71052
rect 68652 70932 68704 70984
rect 30288 70796 30340 70848
rect 34520 70796 34572 70848
rect 79508 70932 79560 70984
rect 81164 70932 81216 70984
rect 83464 70932 83516 70984
rect 85396 70975 85448 70984
rect 85396 70941 85405 70975
rect 85405 70941 85439 70975
rect 85439 70941 85448 70975
rect 85396 70932 85448 70941
rect 87788 70907 87840 70916
rect 87788 70873 87797 70907
rect 87797 70873 87831 70907
rect 87831 70873 87840 70907
rect 87788 70864 87840 70873
rect 93308 70975 93360 70984
rect 93308 70941 93317 70975
rect 93317 70941 93351 70975
rect 93351 70941 93360 70975
rect 93308 70932 93360 70941
rect 93400 70975 93452 70984
rect 93400 70941 93409 70975
rect 93409 70941 93443 70975
rect 93443 70941 93452 70975
rect 97724 71068 97776 71120
rect 93400 70932 93452 70941
rect 96804 70932 96856 70984
rect 94044 70864 94096 70916
rect 97724 70932 97776 70984
rect 98828 71136 98880 71188
rect 99380 71136 99432 71188
rect 98552 71111 98604 71120
rect 98552 71077 98561 71111
rect 98561 71077 98595 71111
rect 98595 71077 98604 71111
rect 98552 71068 98604 71077
rect 98000 71000 98052 71052
rect 98276 71000 98328 71052
rect 99656 71000 99708 71052
rect 100024 71136 100076 71188
rect 100300 71179 100352 71188
rect 100300 71145 100309 71179
rect 100309 71145 100343 71179
rect 100343 71145 100352 71179
rect 100300 71136 100352 71145
rect 105820 71179 105872 71188
rect 105820 71145 105829 71179
rect 105829 71145 105863 71179
rect 105863 71145 105872 71179
rect 105820 71136 105872 71145
rect 107292 71136 107344 71188
rect 101864 71068 101916 71120
rect 106004 71068 106056 71120
rect 98644 70975 98696 70984
rect 98644 70941 98653 70975
rect 98653 70941 98687 70975
rect 98687 70941 98696 70975
rect 98644 70932 98696 70941
rect 98736 70932 98788 70984
rect 99472 70975 99524 70984
rect 99472 70941 99482 70975
rect 99482 70941 99524 70975
rect 99472 70932 99524 70941
rect 100024 70975 100076 70984
rect 100024 70941 100033 70975
rect 100033 70941 100067 70975
rect 100067 70941 100076 70975
rect 100024 70932 100076 70941
rect 101036 70975 101088 70984
rect 101036 70941 101045 70975
rect 101045 70941 101079 70975
rect 101079 70941 101088 70975
rect 101036 70932 101088 70941
rect 101956 70932 102008 70984
rect 102140 70975 102192 70984
rect 102140 70941 102149 70975
rect 102149 70941 102183 70975
rect 102183 70941 102192 70975
rect 102140 70932 102192 70941
rect 103612 71000 103664 71052
rect 103796 71000 103848 71052
rect 105268 71000 105320 71052
rect 105544 71043 105596 71052
rect 105544 71009 105553 71043
rect 105553 71009 105587 71043
rect 105587 71009 105596 71043
rect 105544 71000 105596 71009
rect 106188 71000 106240 71052
rect 102784 70932 102836 70984
rect 103428 70932 103480 70984
rect 105820 70932 105872 70984
rect 108488 70975 108540 70984
rect 56140 70796 56192 70848
rect 72700 70839 72752 70848
rect 72700 70805 72709 70839
rect 72709 70805 72743 70839
rect 72743 70805 72752 70839
rect 72700 70796 72752 70805
rect 89260 70796 89312 70848
rect 92940 70839 92992 70848
rect 92940 70805 92949 70839
rect 92949 70805 92983 70839
rect 92983 70805 92992 70839
rect 92940 70796 92992 70805
rect 93032 70796 93084 70848
rect 93860 70839 93912 70848
rect 93860 70805 93869 70839
rect 93869 70805 93903 70839
rect 93903 70805 93912 70839
rect 93860 70796 93912 70805
rect 96896 70839 96948 70848
rect 96896 70805 96905 70839
rect 96905 70805 96939 70839
rect 96939 70805 96948 70839
rect 96896 70796 96948 70805
rect 97540 70796 97592 70848
rect 97908 70796 97960 70848
rect 98000 70839 98052 70848
rect 98000 70805 98009 70839
rect 98009 70805 98043 70839
rect 98043 70805 98052 70839
rect 98000 70796 98052 70805
rect 103060 70864 103112 70916
rect 105084 70864 105136 70916
rect 105544 70864 105596 70916
rect 98460 70796 98512 70848
rect 98920 70796 98972 70848
rect 100024 70796 100076 70848
rect 101772 70796 101824 70848
rect 103152 70839 103204 70848
rect 103152 70805 103161 70839
rect 103161 70805 103195 70839
rect 103195 70805 103204 70839
rect 103152 70796 103204 70805
rect 105636 70839 105688 70848
rect 105636 70805 105645 70839
rect 105645 70805 105679 70839
rect 105679 70805 105688 70839
rect 105636 70796 105688 70805
rect 108488 70941 108497 70975
rect 108497 70941 108531 70975
rect 108531 70941 108540 70975
rect 108488 70932 108540 70941
rect 4874 70694 4926 70746
rect 4938 70694 4990 70746
rect 5002 70694 5054 70746
rect 5066 70694 5118 70746
rect 5130 70694 5182 70746
rect 35594 70694 35646 70746
rect 35658 70694 35710 70746
rect 35722 70694 35774 70746
rect 35786 70694 35838 70746
rect 35850 70694 35902 70746
rect 66314 70694 66366 70746
rect 66378 70694 66430 70746
rect 66442 70694 66494 70746
rect 66506 70694 66558 70746
rect 66570 70694 66622 70746
rect 97034 70694 97086 70746
rect 97098 70694 97150 70746
rect 97162 70694 97214 70746
rect 97226 70694 97278 70746
rect 97290 70694 97342 70746
rect 30564 70635 30616 70644
rect 30564 70601 30573 70635
rect 30573 70601 30607 70635
rect 30607 70601 30616 70635
rect 30564 70592 30616 70601
rect 28448 70524 28500 70576
rect 34520 70635 34572 70644
rect 34520 70601 34529 70635
rect 34529 70601 34563 70635
rect 34563 70601 34572 70635
rect 34520 70592 34572 70601
rect 87788 70592 87840 70644
rect 88156 70592 88208 70644
rect 93216 70592 93268 70644
rect 97080 70635 97132 70644
rect 97080 70601 97089 70635
rect 97089 70601 97123 70635
rect 97123 70601 97132 70635
rect 97080 70592 97132 70601
rect 31668 70499 31720 70508
rect 31668 70465 31686 70499
rect 31686 70465 31720 70499
rect 31668 70456 31720 70465
rect 31852 70456 31904 70508
rect 35532 70524 35584 70576
rect 84844 70524 84896 70576
rect 90364 70524 90416 70576
rect 34520 70388 34572 70440
rect 88800 70456 88852 70508
rect 97080 70456 97132 70508
rect 97264 70499 97316 70508
rect 97264 70465 97273 70499
rect 97273 70465 97307 70499
rect 97307 70465 97316 70499
rect 97264 70456 97316 70465
rect 41144 70388 41196 70440
rect 91008 70388 91060 70440
rect 96804 70388 96856 70440
rect 97908 70524 97960 70576
rect 97816 70456 97868 70508
rect 98184 70499 98236 70508
rect 98184 70465 98193 70499
rect 98193 70465 98227 70499
rect 98227 70465 98236 70499
rect 98184 70456 98236 70465
rect 98368 70524 98420 70576
rect 99472 70635 99524 70644
rect 99472 70601 99481 70635
rect 99481 70601 99515 70635
rect 99515 70601 99524 70635
rect 99472 70592 99524 70601
rect 99656 70524 99708 70576
rect 103612 70635 103664 70644
rect 103612 70601 103621 70635
rect 103621 70601 103655 70635
rect 103655 70601 103664 70635
rect 103612 70592 103664 70601
rect 105268 70592 105320 70644
rect 106188 70635 106240 70644
rect 106188 70601 106197 70635
rect 106197 70601 106231 70635
rect 106231 70601 106240 70635
rect 106188 70592 106240 70601
rect 108120 70592 108172 70644
rect 105544 70524 105596 70576
rect 105636 70524 105688 70576
rect 106004 70567 106056 70576
rect 106004 70533 106013 70567
rect 106013 70533 106047 70567
rect 106047 70533 106056 70567
rect 106004 70524 106056 70533
rect 97448 70388 97500 70440
rect 97632 70388 97684 70440
rect 97908 70388 97960 70440
rect 98552 70499 98604 70508
rect 98552 70465 98561 70499
rect 98561 70465 98595 70499
rect 98595 70465 98604 70499
rect 98552 70456 98604 70465
rect 98092 70363 98144 70372
rect 98092 70329 98101 70363
rect 98101 70329 98135 70363
rect 98135 70329 98144 70363
rect 98092 70320 98144 70329
rect 99196 70388 99248 70440
rect 99380 70499 99432 70508
rect 99380 70465 99389 70499
rect 99389 70465 99423 70499
rect 99423 70465 99432 70499
rect 99380 70456 99432 70465
rect 100208 70499 100260 70508
rect 100208 70465 100217 70499
rect 100217 70465 100251 70499
rect 100251 70465 100260 70499
rect 100208 70456 100260 70465
rect 101312 70456 101364 70508
rect 102140 70456 102192 70508
rect 103888 70456 103940 70508
rect 105084 70456 105136 70508
rect 106280 70499 106332 70508
rect 106280 70465 106289 70499
rect 106289 70465 106323 70499
rect 106323 70465 106332 70499
rect 106280 70456 106332 70465
rect 108488 70499 108540 70508
rect 108488 70465 108497 70499
rect 108497 70465 108531 70499
rect 108531 70465 108540 70499
rect 108488 70456 108540 70465
rect 101864 70388 101916 70440
rect 103152 70388 103204 70440
rect 104992 70388 105044 70440
rect 105360 70431 105412 70440
rect 105360 70397 105369 70431
rect 105369 70397 105403 70431
rect 105403 70397 105412 70431
rect 105360 70388 105412 70397
rect 102324 70363 102376 70372
rect 102324 70329 102333 70363
rect 102333 70329 102367 70363
rect 102367 70329 102376 70363
rect 102324 70320 102376 70329
rect 105544 70320 105596 70372
rect 107936 70388 107988 70440
rect 93308 70295 93360 70304
rect 93308 70261 93317 70295
rect 93317 70261 93351 70295
rect 93351 70261 93360 70295
rect 93308 70252 93360 70261
rect 99748 70252 99800 70304
rect 105176 70252 105228 70304
rect 105636 70295 105688 70304
rect 105636 70261 105645 70295
rect 105645 70261 105679 70295
rect 105679 70261 105688 70295
rect 105636 70252 105688 70261
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 34934 70150 34986 70202
rect 34998 70150 35050 70202
rect 35062 70150 35114 70202
rect 35126 70150 35178 70202
rect 35190 70150 35242 70202
rect 65654 70150 65706 70202
rect 65718 70150 65770 70202
rect 65782 70150 65834 70202
rect 65846 70150 65898 70202
rect 65910 70150 65962 70202
rect 96374 70150 96426 70202
rect 96438 70150 96490 70202
rect 96502 70150 96554 70202
rect 96566 70150 96618 70202
rect 96630 70150 96682 70202
rect 31852 70048 31904 70100
rect 35532 70091 35584 70100
rect 35532 70057 35541 70091
rect 35541 70057 35575 70091
rect 35575 70057 35584 70091
rect 35532 70048 35584 70057
rect 32956 69980 33008 70032
rect 72884 70048 72936 70100
rect 38660 69912 38712 69964
rect 79508 69955 79560 69964
rect 79508 69921 79517 69955
rect 79517 69921 79551 69955
rect 79551 69921 79560 69955
rect 79508 69912 79560 69921
rect 81164 70091 81216 70100
rect 81164 70057 81173 70091
rect 81173 70057 81207 70091
rect 81207 70057 81216 70091
rect 81164 70048 81216 70057
rect 89720 70091 89772 70100
rect 89720 70057 89729 70091
rect 89729 70057 89763 70091
rect 89763 70057 89772 70091
rect 89720 70048 89772 70057
rect 90640 70048 90692 70100
rect 97540 70048 97592 70100
rect 99196 70048 99248 70100
rect 99380 70048 99432 70100
rect 99840 70048 99892 70100
rect 100208 70048 100260 70100
rect 88340 69980 88392 70032
rect 90364 69980 90416 70032
rect 95240 69980 95292 70032
rect 97264 69980 97316 70032
rect 97908 69980 97960 70032
rect 98644 69980 98696 70032
rect 101956 70048 102008 70100
rect 105728 70048 105780 70100
rect 83096 69912 83148 69964
rect 85396 69912 85448 69964
rect 79324 69887 79376 69896
rect 79324 69853 79333 69887
rect 79333 69853 79367 69887
rect 79367 69853 79376 69887
rect 79324 69844 79376 69853
rect 45100 69776 45152 69828
rect 31668 69708 31720 69760
rect 66720 69751 66772 69760
rect 66720 69717 66729 69751
rect 66729 69717 66763 69751
rect 66763 69717 66772 69751
rect 66720 69708 66772 69717
rect 72424 69708 72476 69760
rect 77852 69819 77904 69828
rect 77852 69785 77886 69819
rect 77886 69785 77904 69819
rect 77852 69776 77904 69785
rect 86776 69844 86828 69896
rect 90364 69887 90416 69896
rect 90364 69853 90373 69887
rect 90373 69853 90407 69887
rect 90407 69853 90416 69887
rect 90364 69844 90416 69853
rect 90640 69955 90692 69964
rect 90640 69921 90649 69955
rect 90649 69921 90683 69955
rect 90683 69921 90692 69955
rect 90640 69912 90692 69921
rect 95700 69912 95752 69964
rect 97816 69912 97868 69964
rect 94320 69844 94372 69896
rect 94872 69844 94924 69896
rect 96160 69844 96212 69896
rect 97540 69844 97592 69896
rect 99012 69887 99064 69896
rect 79324 69708 79376 69760
rect 92480 69776 92532 69828
rect 93768 69776 93820 69828
rect 94780 69751 94832 69760
rect 94780 69717 94789 69751
rect 94789 69717 94823 69751
rect 94823 69717 94832 69751
rect 94780 69708 94832 69717
rect 96068 69708 96120 69760
rect 97448 69776 97500 69828
rect 98184 69776 98236 69828
rect 99012 69853 99021 69887
rect 99021 69853 99055 69887
rect 99055 69853 99064 69887
rect 99012 69844 99064 69853
rect 99472 69844 99524 69896
rect 99748 69887 99800 69896
rect 99748 69853 99757 69887
rect 99757 69853 99791 69887
rect 99791 69853 99800 69887
rect 99748 69844 99800 69853
rect 101404 69912 101456 69964
rect 100484 69887 100536 69896
rect 100484 69853 100493 69887
rect 100493 69853 100527 69887
rect 100527 69853 100536 69887
rect 100484 69844 100536 69853
rect 100852 69887 100904 69896
rect 100852 69853 100861 69887
rect 100861 69853 100895 69887
rect 100895 69853 100904 69887
rect 100852 69844 100904 69853
rect 100944 69887 100996 69896
rect 100944 69853 100953 69887
rect 100953 69853 100987 69887
rect 100987 69853 100996 69887
rect 100944 69844 100996 69853
rect 101312 69887 101364 69896
rect 101312 69853 101321 69887
rect 101321 69853 101355 69887
rect 101355 69853 101364 69887
rect 101312 69844 101364 69853
rect 101496 69887 101548 69896
rect 101496 69853 101505 69887
rect 101505 69853 101539 69887
rect 101539 69853 101548 69887
rect 101496 69844 101548 69853
rect 101956 69955 102008 69964
rect 101956 69921 101965 69955
rect 101965 69921 101999 69955
rect 101999 69921 102008 69955
rect 101956 69912 102008 69921
rect 103612 69912 103664 69964
rect 104992 69912 105044 69964
rect 104900 69844 104952 69896
rect 105084 69887 105136 69896
rect 105084 69853 105093 69887
rect 105093 69853 105127 69887
rect 105127 69853 105136 69887
rect 105084 69844 105136 69853
rect 105268 69887 105320 69896
rect 105268 69853 105277 69887
rect 105277 69853 105311 69887
rect 105311 69853 105320 69887
rect 105268 69844 105320 69853
rect 108488 69887 108540 69896
rect 108488 69853 108497 69887
rect 108497 69853 108531 69887
rect 108531 69853 108540 69887
rect 108488 69844 108540 69853
rect 100760 69819 100812 69828
rect 100760 69785 100769 69819
rect 100769 69785 100803 69819
rect 100803 69785 100812 69819
rect 100760 69776 100812 69785
rect 101680 69776 101732 69828
rect 105636 69776 105688 69828
rect 96804 69708 96856 69760
rect 99656 69708 99708 69760
rect 100024 69751 100076 69760
rect 100024 69717 100033 69751
rect 100033 69717 100067 69751
rect 100067 69717 100076 69751
rect 100024 69708 100076 69717
rect 100116 69751 100168 69760
rect 100116 69717 100125 69751
rect 100125 69717 100159 69751
rect 100159 69717 100168 69751
rect 100116 69708 100168 69717
rect 100944 69708 100996 69760
rect 102232 69751 102284 69760
rect 102232 69717 102241 69751
rect 102241 69717 102275 69751
rect 102275 69717 102284 69751
rect 102232 69708 102284 69717
rect 103336 69708 103388 69760
rect 104900 69751 104952 69760
rect 104900 69717 104909 69751
rect 104909 69717 104943 69751
rect 104943 69717 104952 69751
rect 104900 69708 104952 69717
rect 4874 69606 4926 69658
rect 4938 69606 4990 69658
rect 5002 69606 5054 69658
rect 5066 69606 5118 69658
rect 5130 69606 5182 69658
rect 35594 69606 35646 69658
rect 35658 69606 35710 69658
rect 35722 69606 35774 69658
rect 35786 69606 35838 69658
rect 35850 69606 35902 69658
rect 66314 69606 66366 69658
rect 66378 69606 66430 69658
rect 66442 69606 66494 69658
rect 66506 69606 66558 69658
rect 66570 69606 66622 69658
rect 97034 69606 97086 69658
rect 97098 69606 97150 69658
rect 97162 69606 97214 69658
rect 97226 69606 97278 69658
rect 97290 69606 97342 69658
rect 42432 69547 42484 69556
rect 42432 69513 42441 69547
rect 42441 69513 42475 69547
rect 42475 69513 42484 69547
rect 42432 69504 42484 69513
rect 43720 69368 43772 69420
rect 67180 69436 67232 69488
rect 66720 69368 66772 69420
rect 67364 69504 67416 69556
rect 69112 69504 69164 69556
rect 79324 69504 79376 69556
rect 88800 69547 88852 69556
rect 88800 69513 88809 69547
rect 88809 69513 88843 69547
rect 88843 69513 88852 69547
rect 88800 69504 88852 69513
rect 69020 69368 69072 69420
rect 86316 69368 86368 69420
rect 91560 69479 91612 69488
rect 91560 69445 91569 69479
rect 91569 69445 91603 69479
rect 91603 69445 91612 69479
rect 91560 69436 91612 69445
rect 89720 69368 89772 69420
rect 91836 69411 91888 69420
rect 91836 69377 91845 69411
rect 91845 69377 91879 69411
rect 91879 69377 91888 69411
rect 91836 69368 91888 69377
rect 92940 69504 92992 69556
rect 97816 69547 97868 69556
rect 97816 69513 97825 69547
rect 97825 69513 97859 69547
rect 97859 69513 97868 69547
rect 97816 69504 97868 69513
rect 99472 69504 99524 69556
rect 100944 69504 100996 69556
rect 92296 69479 92348 69488
rect 92296 69445 92305 69479
rect 92305 69445 92339 69479
rect 92339 69445 92348 69479
rect 92296 69436 92348 69445
rect 92480 69368 92532 69420
rect 93032 69368 93084 69420
rect 98276 69368 98328 69420
rect 98736 69368 98788 69420
rect 42156 69207 42208 69216
rect 42156 69173 42165 69207
rect 42165 69173 42199 69207
rect 42199 69173 42208 69207
rect 42156 69164 42208 69173
rect 66444 69343 66496 69352
rect 66444 69309 66453 69343
rect 66453 69309 66487 69343
rect 66487 69309 66496 69343
rect 66444 69300 66496 69309
rect 89076 69343 89128 69352
rect 89076 69309 89085 69343
rect 89085 69309 89119 69343
rect 89119 69309 89128 69343
rect 89076 69300 89128 69309
rect 94964 69300 95016 69352
rect 95884 69300 95936 69352
rect 98920 69411 98972 69420
rect 98920 69377 98929 69411
rect 98929 69377 98963 69411
rect 98963 69377 98972 69411
rect 98920 69368 98972 69377
rect 99104 69411 99156 69420
rect 99104 69377 99113 69411
rect 99113 69377 99147 69411
rect 99147 69377 99156 69411
rect 99104 69368 99156 69377
rect 99564 69436 99616 69488
rect 100852 69436 100904 69488
rect 99380 69368 99432 69420
rect 99656 69411 99708 69420
rect 99656 69377 99665 69411
rect 99665 69377 99699 69411
rect 99699 69377 99708 69411
rect 99656 69368 99708 69377
rect 99748 69368 99800 69420
rect 100760 69368 100812 69420
rect 101496 69368 101548 69420
rect 100852 69300 100904 69352
rect 102324 69368 102376 69420
rect 103244 69368 103296 69420
rect 103336 69411 103388 69420
rect 103336 69377 103345 69411
rect 103345 69377 103379 69411
rect 103379 69377 103388 69411
rect 103336 69368 103388 69377
rect 103520 69411 103572 69420
rect 103520 69377 103529 69411
rect 103529 69377 103563 69411
rect 103563 69377 103572 69411
rect 103520 69368 103572 69377
rect 102048 69300 102100 69352
rect 102416 69343 102468 69352
rect 102416 69309 102425 69343
rect 102425 69309 102459 69343
rect 102459 69309 102468 69343
rect 102416 69300 102468 69309
rect 102968 69343 103020 69352
rect 102968 69309 102977 69343
rect 102977 69309 103011 69343
rect 103011 69309 103020 69343
rect 102968 69300 103020 69309
rect 104624 69368 104676 69420
rect 104992 69411 105044 69420
rect 104992 69377 105001 69411
rect 105001 69377 105035 69411
rect 105035 69377 105044 69411
rect 104992 69368 105044 69377
rect 43812 69164 43864 69216
rect 61476 69164 61528 69216
rect 74540 69164 74592 69216
rect 91744 69164 91796 69216
rect 92756 69207 92808 69216
rect 92756 69173 92765 69207
rect 92765 69173 92799 69207
rect 92799 69173 92808 69207
rect 92756 69164 92808 69173
rect 98920 69164 98972 69216
rect 99656 69164 99708 69216
rect 100484 69207 100536 69216
rect 100484 69173 100493 69207
rect 100493 69173 100527 69207
rect 100527 69173 100536 69207
rect 100484 69164 100536 69173
rect 101128 69164 101180 69216
rect 101772 69207 101824 69216
rect 101772 69173 101781 69207
rect 101781 69173 101815 69207
rect 101815 69173 101824 69207
rect 101772 69164 101824 69173
rect 103428 69164 103480 69216
rect 103612 69207 103664 69216
rect 103612 69173 103621 69207
rect 103621 69173 103655 69207
rect 103655 69173 103664 69207
rect 103612 69164 103664 69173
rect 104532 69164 104584 69216
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 96374 69062 96426 69114
rect 96438 69062 96490 69114
rect 96502 69062 96554 69114
rect 96566 69062 96618 69114
rect 96630 69062 96682 69114
rect 43812 68960 43864 69012
rect 42708 68892 42760 68944
rect 58624 69003 58676 69012
rect 58624 68969 58633 69003
rect 58633 68969 58667 69003
rect 58667 68969 58676 69003
rect 58624 68960 58676 68969
rect 67364 69003 67416 69012
rect 67364 68969 67373 69003
rect 67373 68969 67407 69003
rect 67407 68969 67416 69003
rect 67364 68960 67416 68969
rect 70400 68892 70452 68944
rect 89720 68960 89772 69012
rect 68560 68756 68612 68808
rect 86868 68756 86920 68808
rect 93308 68960 93360 69012
rect 91744 68824 91796 68876
rect 43720 68688 43772 68740
rect 58716 68731 58768 68740
rect 58716 68697 58725 68731
rect 58725 68697 58759 68731
rect 58759 68697 58768 68731
rect 58716 68688 58768 68697
rect 66076 68688 66128 68740
rect 95976 68960 96028 69012
rect 98276 69003 98328 69012
rect 98276 68969 98285 69003
rect 98285 68969 98319 69003
rect 98319 68969 98328 69003
rect 98276 68960 98328 68969
rect 100852 68960 100904 69012
rect 102968 68960 103020 69012
rect 104808 68960 104860 69012
rect 104992 68960 105044 69012
rect 105268 69003 105320 69012
rect 105268 68969 105277 69003
rect 105277 68969 105311 69003
rect 105311 68969 105320 69003
rect 105268 68960 105320 68969
rect 100300 68892 100352 68944
rect 95240 68824 95292 68876
rect 95516 68867 95568 68876
rect 95516 68833 95525 68867
rect 95525 68833 95559 68867
rect 95559 68833 95568 68867
rect 95516 68824 95568 68833
rect 96160 68824 96212 68876
rect 46480 68663 46532 68672
rect 46480 68629 46489 68663
rect 46489 68629 46523 68663
rect 46523 68629 46532 68663
rect 46480 68620 46532 68629
rect 61476 68663 61528 68672
rect 61476 68629 61485 68663
rect 61485 68629 61519 68663
rect 61519 68629 61528 68663
rect 61476 68620 61528 68629
rect 86776 68663 86828 68672
rect 86776 68629 86785 68663
rect 86785 68629 86819 68663
rect 86819 68629 86828 68663
rect 86776 68620 86828 68629
rect 89260 68620 89312 68672
rect 94964 68756 95016 68808
rect 96068 68756 96120 68808
rect 97448 68799 97500 68808
rect 97448 68765 97457 68799
rect 97457 68765 97491 68799
rect 97491 68765 97500 68799
rect 97448 68756 97500 68765
rect 99748 68756 99800 68808
rect 100300 68756 100352 68808
rect 101404 68824 101456 68876
rect 101772 68824 101824 68876
rect 102232 68867 102284 68876
rect 102232 68833 102241 68867
rect 102241 68833 102275 68867
rect 102275 68833 102284 68867
rect 102232 68824 102284 68833
rect 103152 68824 103204 68876
rect 101128 68756 101180 68808
rect 101220 68756 101272 68808
rect 103060 68799 103112 68808
rect 103060 68765 103069 68799
rect 103069 68765 103103 68799
rect 103103 68765 103112 68799
rect 103060 68756 103112 68765
rect 103244 68756 103296 68808
rect 103428 68799 103480 68808
rect 103428 68765 103437 68799
rect 103437 68765 103471 68799
rect 103471 68765 103480 68799
rect 103428 68756 103480 68765
rect 98000 68688 98052 68740
rect 98736 68688 98788 68740
rect 99196 68688 99248 68740
rect 94504 68663 94556 68672
rect 94504 68629 94513 68663
rect 94513 68629 94547 68663
rect 94547 68629 94556 68663
rect 94504 68620 94556 68629
rect 95148 68663 95200 68672
rect 95148 68629 95157 68663
rect 95157 68629 95191 68663
rect 95191 68629 95200 68663
rect 95148 68620 95200 68629
rect 96896 68663 96948 68672
rect 96896 68629 96905 68663
rect 96905 68629 96939 68663
rect 96939 68629 96948 68663
rect 96896 68620 96948 68629
rect 97908 68620 97960 68672
rect 99656 68620 99708 68672
rect 100944 68688 100996 68740
rect 103612 68799 103664 68808
rect 103612 68765 103621 68799
rect 103621 68765 103655 68799
rect 103655 68765 103664 68799
rect 103612 68756 103664 68765
rect 103704 68799 103756 68808
rect 103704 68765 103713 68799
rect 103713 68765 103747 68799
rect 103747 68765 103756 68799
rect 103704 68756 103756 68765
rect 101128 68620 101180 68672
rect 101220 68620 101272 68672
rect 102048 68663 102100 68672
rect 102048 68629 102057 68663
rect 102057 68629 102091 68663
rect 102091 68629 102100 68663
rect 102048 68620 102100 68629
rect 102876 68620 102928 68672
rect 104624 68756 104676 68808
rect 104808 68799 104860 68808
rect 104808 68765 104817 68799
rect 104817 68765 104851 68799
rect 104851 68765 104860 68799
rect 104808 68756 104860 68765
rect 105360 68824 105412 68876
rect 104900 68688 104952 68740
rect 105176 68688 105228 68740
rect 105452 68731 105504 68740
rect 105452 68697 105461 68731
rect 105461 68697 105495 68731
rect 105495 68697 105504 68731
rect 105452 68688 105504 68697
rect 104440 68620 104492 68672
rect 4874 68518 4926 68570
rect 4938 68518 4990 68570
rect 5002 68518 5054 68570
rect 5066 68518 5118 68570
rect 5130 68518 5182 68570
rect 35594 68518 35646 68570
rect 35658 68518 35710 68570
rect 35722 68518 35774 68570
rect 35786 68518 35838 68570
rect 35850 68518 35902 68570
rect 66314 68518 66366 68570
rect 66378 68518 66430 68570
rect 66442 68518 66494 68570
rect 66506 68518 66558 68570
rect 66570 68518 66622 68570
rect 97034 68518 97086 68570
rect 97098 68518 97150 68570
rect 97162 68518 97214 68570
rect 97226 68518 97278 68570
rect 97290 68518 97342 68570
rect 38660 68459 38712 68468
rect 38660 68425 38669 68459
rect 38669 68425 38703 68459
rect 38703 68425 38712 68459
rect 38660 68416 38712 68425
rect 38844 68459 38896 68468
rect 38844 68425 38853 68459
rect 38853 68425 38887 68459
rect 38887 68425 38896 68459
rect 38844 68416 38896 68425
rect 91560 68459 91612 68468
rect 91560 68425 91569 68459
rect 91569 68425 91603 68459
rect 91603 68425 91612 68459
rect 91560 68416 91612 68425
rect 92940 68416 92992 68468
rect 96068 68416 96120 68468
rect 39948 68323 40000 68332
rect 42156 68348 42208 68400
rect 91008 68348 91060 68400
rect 91928 68391 91980 68400
rect 91928 68357 91937 68391
rect 91937 68357 91971 68391
rect 91971 68357 91980 68391
rect 91928 68348 91980 68357
rect 92296 68348 92348 68400
rect 94780 68348 94832 68400
rect 98184 68459 98236 68468
rect 98184 68425 98193 68459
rect 98193 68425 98227 68459
rect 98227 68425 98236 68459
rect 98184 68416 98236 68425
rect 100116 68416 100168 68468
rect 100300 68416 100352 68468
rect 39948 68289 39966 68323
rect 39966 68289 40000 68323
rect 39948 68280 40000 68289
rect 95240 68323 95292 68332
rect 95240 68289 95249 68323
rect 95249 68289 95283 68323
rect 95283 68289 95292 68323
rect 95240 68280 95292 68289
rect 96160 68323 96212 68332
rect 96160 68289 96169 68323
rect 96169 68289 96203 68323
rect 96203 68289 96212 68323
rect 96160 68280 96212 68289
rect 96252 68280 96304 68332
rect 97448 68280 97500 68332
rect 95056 68255 95108 68264
rect 95056 68221 95065 68255
rect 95065 68221 95099 68255
rect 95099 68221 95108 68255
rect 95056 68212 95108 68221
rect 98000 68348 98052 68400
rect 99932 68348 99984 68400
rect 101864 68416 101916 68468
rect 102324 68416 102376 68468
rect 102416 68416 102468 68468
rect 103612 68416 103664 68468
rect 97632 68280 97684 68332
rect 98552 68280 98604 68332
rect 99288 68323 99340 68332
rect 99288 68289 99297 68323
rect 99297 68289 99331 68323
rect 99331 68289 99340 68323
rect 99288 68280 99340 68289
rect 99564 68323 99616 68332
rect 99564 68289 99573 68323
rect 99573 68289 99607 68323
rect 99607 68289 99616 68323
rect 99564 68280 99616 68289
rect 99840 68323 99892 68332
rect 99840 68289 99849 68323
rect 99849 68289 99883 68323
rect 99883 68289 99892 68323
rect 99840 68280 99892 68289
rect 100208 68280 100260 68332
rect 95792 68144 95844 68196
rect 97908 68212 97960 68264
rect 99472 68212 99524 68264
rect 100668 68323 100720 68332
rect 100668 68289 100677 68323
rect 100677 68289 100711 68323
rect 100711 68289 100720 68323
rect 100668 68280 100720 68289
rect 100852 68280 100904 68332
rect 101220 68348 101272 68400
rect 101404 68391 101456 68400
rect 101404 68357 101413 68391
rect 101413 68357 101447 68391
rect 101447 68357 101456 68391
rect 101404 68348 101456 68357
rect 101128 68323 101180 68332
rect 101128 68289 101137 68323
rect 101137 68289 101171 68323
rect 101171 68289 101180 68323
rect 101128 68280 101180 68289
rect 93400 68076 93452 68128
rect 95148 68119 95200 68128
rect 95148 68085 95157 68119
rect 95157 68085 95191 68119
rect 95191 68085 95200 68119
rect 95148 68076 95200 68085
rect 95332 68076 95384 68128
rect 95884 68119 95936 68128
rect 95884 68085 95893 68119
rect 95893 68085 95927 68119
rect 95927 68085 95936 68119
rect 95884 68076 95936 68085
rect 96068 68076 96120 68128
rect 96712 68076 96764 68128
rect 101036 68212 101088 68264
rect 100300 68144 100352 68196
rect 102232 68280 102284 68332
rect 103336 68280 103388 68332
rect 103704 68280 103756 68332
rect 105268 68416 105320 68468
rect 104900 68323 104952 68332
rect 104900 68289 104909 68323
rect 104909 68289 104943 68323
rect 104943 68289 104952 68323
rect 104900 68280 104952 68289
rect 105176 68323 105228 68332
rect 105176 68289 105185 68323
rect 105185 68289 105219 68323
rect 105219 68289 105228 68323
rect 105176 68280 105228 68289
rect 100576 68076 100628 68128
rect 104532 68255 104584 68264
rect 104532 68221 104541 68255
rect 104541 68221 104575 68255
rect 104575 68221 104584 68255
rect 104532 68212 104584 68221
rect 105452 68212 105504 68264
rect 101956 68144 102008 68196
rect 102508 68144 102560 68196
rect 104624 68144 104676 68196
rect 103980 68119 104032 68128
rect 103980 68085 103989 68119
rect 103989 68085 104023 68119
rect 104023 68085 104032 68119
rect 103980 68076 104032 68085
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 96374 67974 96426 68026
rect 96438 67974 96490 68026
rect 96502 67974 96554 68026
rect 96566 67974 96618 68026
rect 96630 67974 96682 68026
rect 89076 67872 89128 67924
rect 89444 67872 89496 67924
rect 90824 67872 90876 67924
rect 91928 67872 91980 67924
rect 98736 67872 98788 67924
rect 99288 67872 99340 67924
rect 100024 67872 100076 67924
rect 101680 67915 101732 67924
rect 101680 67881 101689 67915
rect 101689 67881 101723 67915
rect 101723 67881 101732 67915
rect 101680 67872 101732 67881
rect 101772 67872 101824 67924
rect 102692 67872 102744 67924
rect 107936 67915 107988 67924
rect 107936 67881 107945 67915
rect 107945 67881 107979 67915
rect 107979 67881 107988 67915
rect 107936 67872 107988 67881
rect 86776 67736 86828 67788
rect 86040 67668 86092 67720
rect 87144 67668 87196 67720
rect 94412 67804 94464 67856
rect 94964 67779 95016 67788
rect 94964 67745 94973 67779
rect 94973 67745 95007 67779
rect 95007 67745 95016 67779
rect 94964 67736 95016 67745
rect 95700 67736 95752 67788
rect 95884 67779 95936 67788
rect 95884 67745 95893 67779
rect 95893 67745 95927 67779
rect 95927 67745 95936 67779
rect 95884 67736 95936 67745
rect 89260 67668 89312 67720
rect 70216 67600 70268 67652
rect 74356 67600 74408 67652
rect 89720 67643 89772 67652
rect 89720 67609 89747 67643
rect 89747 67609 89772 67643
rect 89720 67600 89772 67609
rect 95332 67711 95384 67720
rect 95332 67677 95341 67711
rect 95341 67677 95375 67711
rect 95375 67677 95384 67711
rect 95332 67668 95384 67677
rect 96252 67668 96304 67720
rect 98828 67804 98880 67856
rect 97908 67736 97960 67788
rect 98552 67779 98604 67788
rect 98552 67745 98561 67779
rect 98561 67745 98595 67779
rect 98595 67745 98604 67779
rect 98552 67736 98604 67745
rect 99196 67804 99248 67856
rect 99748 67804 99800 67856
rect 100760 67804 100812 67856
rect 99472 67736 99524 67788
rect 102876 67804 102928 67856
rect 102968 67847 103020 67856
rect 102968 67813 102977 67847
rect 102977 67813 103011 67847
rect 103011 67813 103020 67847
rect 102968 67804 103020 67813
rect 102324 67779 102376 67788
rect 102324 67745 102333 67779
rect 102333 67745 102367 67779
rect 102367 67745 102376 67779
rect 102324 67736 102376 67745
rect 89996 67600 90048 67652
rect 91008 67600 91060 67652
rect 98276 67600 98328 67652
rect 99104 67668 99156 67720
rect 101036 67668 101088 67720
rect 101680 67668 101732 67720
rect 98920 67600 98972 67652
rect 99748 67600 99800 67652
rect 100300 67600 100352 67652
rect 101956 67711 102008 67720
rect 101956 67677 101965 67711
rect 101965 67677 101999 67711
rect 101999 67677 102008 67711
rect 101956 67668 102008 67677
rect 102140 67711 102192 67720
rect 102140 67677 102149 67711
rect 102149 67677 102183 67711
rect 102183 67677 102192 67711
rect 102140 67668 102192 67677
rect 102232 67705 102284 67720
rect 102232 67671 102241 67705
rect 102241 67671 102275 67705
rect 102275 67671 102284 67705
rect 102232 67668 102284 67671
rect 102508 67711 102560 67720
rect 102508 67677 102517 67711
rect 102517 67677 102551 67711
rect 102551 67677 102560 67711
rect 102508 67668 102560 67677
rect 102692 67668 102744 67720
rect 102784 67711 102836 67720
rect 102784 67677 102793 67711
rect 102793 67677 102827 67711
rect 102827 67677 102836 67711
rect 102784 67668 102836 67677
rect 102416 67600 102468 67652
rect 103704 67668 103756 67720
rect 108488 67711 108540 67720
rect 108488 67677 108497 67711
rect 108497 67677 108531 67711
rect 108531 67677 108540 67711
rect 108488 67668 108540 67677
rect 87420 67532 87472 67584
rect 89076 67575 89128 67584
rect 89076 67541 89085 67575
rect 89085 67541 89119 67575
rect 89119 67541 89128 67575
rect 89076 67532 89128 67541
rect 89352 67532 89404 67584
rect 95332 67532 95384 67584
rect 99656 67532 99708 67584
rect 100852 67532 100904 67584
rect 103336 67600 103388 67652
rect 103152 67575 103204 67584
rect 103152 67541 103161 67575
rect 103161 67541 103195 67575
rect 103195 67541 103204 67575
rect 103152 67532 103204 67541
rect 4874 67430 4926 67482
rect 4938 67430 4990 67482
rect 5002 67430 5054 67482
rect 5066 67430 5118 67482
rect 5130 67430 5182 67482
rect 35594 67430 35646 67482
rect 35658 67430 35710 67482
rect 35722 67430 35774 67482
rect 35786 67430 35838 67482
rect 35850 67430 35902 67482
rect 66314 67430 66366 67482
rect 66378 67430 66430 67482
rect 66442 67430 66494 67482
rect 66506 67430 66558 67482
rect 66570 67430 66622 67482
rect 97034 67430 97086 67482
rect 97098 67430 97150 67482
rect 97162 67430 97214 67482
rect 97226 67430 97278 67482
rect 97290 67430 97342 67482
rect 86868 67328 86920 67380
rect 87420 67328 87472 67380
rect 89352 67328 89404 67380
rect 90180 67328 90232 67380
rect 89904 67303 89956 67312
rect 89904 67269 89913 67303
rect 89913 67269 89947 67303
rect 89947 67269 89956 67303
rect 89904 67260 89956 67269
rect 92940 67371 92992 67380
rect 92940 67337 92949 67371
rect 92949 67337 92983 67371
rect 92983 67337 92992 67371
rect 92940 67328 92992 67337
rect 93400 67371 93452 67380
rect 93400 67337 93409 67371
rect 93409 67337 93443 67371
rect 93443 67337 93452 67371
rect 93400 67328 93452 67337
rect 95240 67328 95292 67380
rect 96804 67371 96856 67380
rect 96804 67337 96831 67371
rect 96831 67337 96856 67371
rect 96804 67328 96856 67337
rect 89352 67192 89404 67244
rect 91192 67235 91244 67244
rect 91192 67201 91201 67235
rect 91201 67201 91235 67235
rect 91235 67201 91244 67235
rect 91192 67192 91244 67201
rect 91468 67260 91520 67312
rect 92572 67260 92624 67312
rect 93032 67260 93084 67312
rect 92756 67192 92808 67244
rect 95976 67192 96028 67244
rect 99104 67328 99156 67380
rect 99564 67328 99616 67380
rect 94504 67124 94556 67176
rect 92204 67056 92256 67108
rect 94780 67056 94832 67108
rect 95516 67124 95568 67176
rect 96896 67124 96948 67176
rect 99656 67235 99708 67244
rect 99656 67201 99665 67235
rect 99665 67201 99699 67235
rect 99699 67201 99708 67235
rect 99656 67192 99708 67201
rect 99840 67260 99892 67312
rect 100024 67303 100076 67312
rect 100024 67269 100033 67303
rect 100033 67269 100067 67303
rect 100067 67269 100076 67303
rect 100024 67260 100076 67269
rect 102416 67328 102468 67380
rect 102784 67328 102836 67380
rect 101312 67260 101364 67312
rect 100116 67124 100168 67176
rect 100852 67192 100904 67244
rect 101956 67260 102008 67312
rect 102876 67303 102928 67312
rect 102876 67269 102885 67303
rect 102885 67269 102919 67303
rect 102919 67269 102928 67303
rect 102876 67260 102928 67269
rect 101772 67235 101824 67244
rect 101772 67201 101781 67235
rect 101781 67201 101815 67235
rect 101815 67201 101824 67235
rect 101772 67192 101824 67201
rect 100944 67124 100996 67176
rect 100576 67056 100628 67108
rect 102232 67192 102284 67244
rect 102600 67192 102652 67244
rect 102968 67235 103020 67244
rect 102968 67201 102977 67235
rect 102977 67201 103011 67235
rect 103011 67201 103020 67235
rect 102968 67192 103020 67201
rect 103520 67260 103572 67312
rect 103980 67260 104032 67312
rect 103704 67235 103756 67244
rect 103704 67201 103713 67235
rect 103713 67201 103747 67235
rect 103747 67201 103756 67235
rect 103704 67192 103756 67201
rect 103152 67124 103204 67176
rect 86776 67031 86828 67040
rect 86776 66997 86785 67031
rect 86785 66997 86819 67031
rect 86819 66997 86828 67031
rect 86776 66988 86828 66997
rect 89812 66988 89864 67040
rect 96160 66988 96212 67040
rect 96896 66988 96948 67040
rect 97080 67031 97132 67040
rect 97080 66997 97089 67031
rect 97089 66997 97123 67031
rect 97123 66997 97132 67031
rect 97080 66988 97132 66997
rect 100668 66988 100720 67040
rect 102048 66988 102100 67040
rect 102876 66988 102928 67040
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 96374 66886 96426 66938
rect 96438 66886 96490 66938
rect 96502 66886 96554 66938
rect 96566 66886 96618 66938
rect 96630 66886 96682 66938
rect 89444 66827 89496 66836
rect 89444 66793 89453 66827
rect 89453 66793 89487 66827
rect 89487 66793 89496 66827
rect 89444 66784 89496 66793
rect 89812 66827 89864 66836
rect 89812 66793 89821 66827
rect 89821 66793 89855 66827
rect 89855 66793 89864 66827
rect 89812 66784 89864 66793
rect 90640 66784 90692 66836
rect 91192 66784 91244 66836
rect 92480 66784 92532 66836
rect 95700 66784 95752 66836
rect 95976 66827 96028 66836
rect 95976 66793 95985 66827
rect 95985 66793 96019 66827
rect 96019 66793 96028 66827
rect 95976 66784 96028 66793
rect 99932 66784 99984 66836
rect 100116 66784 100168 66836
rect 100576 66784 100628 66836
rect 102140 66784 102192 66836
rect 103152 66784 103204 66836
rect 103704 66784 103756 66836
rect 92020 66716 92072 66768
rect 97632 66759 97684 66768
rect 97632 66725 97641 66759
rect 97641 66725 97675 66759
rect 97675 66725 97684 66759
rect 97632 66716 97684 66725
rect 91468 66648 91520 66700
rect 95240 66648 95292 66700
rect 96068 66648 96120 66700
rect 96160 66691 96212 66700
rect 96160 66657 96169 66691
rect 96169 66657 96203 66691
rect 96203 66657 96212 66691
rect 96160 66648 96212 66657
rect 97448 66648 97500 66700
rect 85396 66580 85448 66632
rect 86776 66580 86828 66632
rect 89260 66623 89312 66632
rect 89260 66589 89269 66623
rect 89269 66589 89303 66623
rect 89303 66589 89312 66623
rect 89260 66580 89312 66589
rect 89352 66623 89404 66632
rect 89352 66589 89361 66623
rect 89361 66589 89395 66623
rect 89395 66589 89404 66623
rect 89352 66580 89404 66589
rect 89904 66580 89956 66632
rect 95608 66580 95660 66632
rect 97080 66580 97132 66632
rect 98276 66580 98328 66632
rect 98552 66648 98604 66700
rect 99840 66716 99892 66768
rect 101864 66759 101916 66768
rect 101864 66725 101873 66759
rect 101873 66725 101907 66759
rect 101907 66725 101916 66759
rect 101864 66716 101916 66725
rect 102784 66716 102836 66768
rect 99472 66691 99524 66700
rect 99472 66657 99481 66691
rect 99481 66657 99515 66691
rect 99515 66657 99524 66691
rect 99472 66648 99524 66657
rect 99564 66648 99616 66700
rect 98736 66623 98788 66632
rect 98736 66589 98745 66623
rect 98745 66589 98779 66623
rect 98779 66589 98788 66623
rect 98736 66580 98788 66589
rect 99656 66623 99708 66632
rect 99656 66589 99665 66623
rect 99665 66589 99699 66623
rect 99699 66589 99708 66623
rect 99656 66580 99708 66589
rect 100484 66648 100536 66700
rect 100852 66648 100904 66700
rect 102232 66648 102284 66700
rect 103244 66691 103296 66700
rect 103244 66657 103253 66691
rect 103253 66657 103287 66691
rect 103287 66657 103296 66691
rect 103244 66648 103296 66657
rect 100668 66580 100720 66632
rect 102784 66623 102836 66632
rect 102784 66589 102793 66623
rect 102793 66589 102827 66623
rect 102827 66589 102836 66623
rect 102784 66580 102836 66589
rect 102876 66623 102928 66632
rect 102876 66589 102885 66623
rect 102885 66589 102919 66623
rect 102919 66589 102928 66623
rect 102876 66580 102928 66589
rect 103336 66623 103388 66632
rect 103336 66589 103345 66623
rect 103345 66589 103379 66623
rect 103379 66589 103388 66623
rect 103336 66580 103388 66589
rect 86868 66512 86920 66564
rect 87144 66487 87196 66496
rect 87144 66453 87153 66487
rect 87153 66453 87187 66487
rect 87187 66453 87196 66487
rect 87144 66444 87196 66453
rect 88248 66444 88300 66496
rect 89996 66555 90048 66564
rect 89996 66521 90005 66555
rect 90005 66521 90039 66555
rect 90039 66521 90048 66555
rect 89996 66512 90048 66521
rect 92296 66555 92348 66564
rect 92296 66521 92305 66555
rect 92305 66521 92339 66555
rect 92339 66521 92348 66555
rect 92756 66555 92808 66564
rect 92296 66512 92348 66521
rect 92756 66521 92765 66555
rect 92765 66521 92799 66555
rect 92799 66521 92808 66555
rect 92756 66512 92808 66521
rect 94780 66512 94832 66564
rect 97632 66512 97684 66564
rect 101680 66512 101732 66564
rect 89904 66444 89956 66496
rect 92572 66487 92624 66496
rect 92572 66453 92599 66487
rect 92599 66453 92624 66487
rect 92572 66444 92624 66453
rect 95424 66444 95476 66496
rect 95884 66444 95936 66496
rect 99932 66487 99984 66496
rect 99932 66453 99941 66487
rect 99941 66453 99975 66487
rect 99975 66453 99984 66487
rect 99932 66444 99984 66453
rect 100576 66487 100628 66496
rect 100576 66453 100585 66487
rect 100585 66453 100619 66487
rect 100619 66453 100628 66487
rect 100576 66444 100628 66453
rect 101312 66444 101364 66496
rect 103704 66487 103756 66496
rect 103704 66453 103713 66487
rect 103713 66453 103747 66487
rect 103747 66453 103756 66487
rect 103704 66444 103756 66453
rect 104164 66555 104216 66564
rect 104164 66521 104173 66555
rect 104173 66521 104207 66555
rect 104207 66521 104216 66555
rect 104164 66512 104216 66521
rect 104624 66555 104676 66564
rect 104624 66521 104633 66555
rect 104633 66521 104667 66555
rect 104667 66521 104676 66555
rect 104624 66512 104676 66521
rect 4874 66342 4926 66394
rect 4938 66342 4990 66394
rect 5002 66342 5054 66394
rect 5066 66342 5118 66394
rect 5130 66342 5182 66394
rect 35594 66342 35646 66394
rect 35658 66342 35710 66394
rect 35722 66342 35774 66394
rect 35786 66342 35838 66394
rect 35850 66342 35902 66394
rect 66314 66342 66366 66394
rect 66378 66342 66430 66394
rect 66442 66342 66494 66394
rect 66506 66342 66558 66394
rect 66570 66342 66622 66394
rect 97034 66342 97086 66394
rect 97098 66342 97150 66394
rect 97162 66342 97214 66394
rect 97226 66342 97278 66394
rect 97290 66342 97342 66394
rect 106658 66342 106710 66394
rect 106722 66342 106774 66394
rect 106786 66342 106838 66394
rect 106850 66342 106902 66394
rect 106914 66342 106966 66394
rect 9496 66172 9548 66224
rect 13820 66172 13872 66224
rect 68652 66215 68704 66224
rect 68652 66181 68661 66215
rect 68661 66181 68695 66215
rect 68695 66181 68704 66215
rect 68652 66172 68704 66181
rect 73160 66215 73212 66224
rect 73160 66181 73169 66215
rect 73169 66181 73203 66215
rect 73203 66181 73212 66215
rect 73160 66172 73212 66181
rect 74356 66215 74408 66224
rect 74356 66181 74365 66215
rect 74365 66181 74399 66215
rect 74399 66181 74408 66215
rect 74356 66172 74408 66181
rect 87144 66240 87196 66292
rect 88616 66283 88668 66292
rect 88616 66249 88625 66283
rect 88625 66249 88659 66283
rect 88659 66249 88668 66283
rect 88616 66240 88668 66249
rect 89352 66240 89404 66292
rect 89904 66240 89956 66292
rect 89076 66172 89128 66224
rect 89720 66172 89772 66224
rect 90640 66215 90692 66224
rect 90640 66181 90649 66215
rect 90649 66181 90683 66215
rect 90683 66181 90692 66215
rect 92296 66283 92348 66292
rect 92296 66249 92305 66283
rect 92305 66249 92339 66283
rect 92339 66249 92348 66283
rect 92296 66240 92348 66249
rect 95424 66283 95476 66292
rect 95424 66249 95449 66283
rect 95449 66249 95476 66283
rect 95424 66240 95476 66249
rect 95608 66283 95660 66292
rect 95608 66249 95617 66283
rect 95617 66249 95651 66283
rect 95651 66249 95660 66283
rect 95608 66240 95660 66249
rect 95792 66283 95844 66292
rect 95792 66249 95801 66283
rect 95801 66249 95835 66283
rect 95835 66249 95844 66283
rect 95792 66240 95844 66249
rect 97448 66240 97500 66292
rect 97632 66240 97684 66292
rect 103980 66240 104032 66292
rect 104164 66240 104216 66292
rect 90640 66172 90692 66181
rect 86868 66104 86920 66156
rect 88248 66147 88300 66156
rect 88248 66113 88257 66147
rect 88257 66113 88291 66147
rect 88291 66113 88300 66147
rect 88248 66104 88300 66113
rect 89260 66104 89312 66156
rect 90180 66147 90232 66156
rect 90180 66113 90189 66147
rect 90189 66113 90223 66147
rect 90223 66113 90232 66147
rect 90180 66104 90232 66113
rect 90732 66147 90784 66156
rect 90732 66113 90741 66147
rect 90741 66113 90775 66147
rect 90775 66113 90784 66147
rect 90732 66104 90784 66113
rect 88616 66036 88668 66088
rect 90824 66079 90876 66088
rect 90824 66045 90833 66079
rect 90833 66045 90867 66079
rect 90867 66045 90876 66079
rect 90824 66036 90876 66045
rect 92572 66104 92624 66156
rect 94136 66147 94188 66156
rect 92388 66036 92440 66088
rect 94136 66113 94145 66147
rect 94145 66113 94179 66147
rect 94179 66113 94188 66147
rect 94136 66104 94188 66113
rect 94780 66147 94832 66156
rect 94780 66113 94789 66147
rect 94789 66113 94823 66147
rect 94823 66113 94832 66147
rect 94780 66104 94832 66113
rect 95240 66215 95292 66224
rect 95240 66181 95249 66215
rect 95249 66181 95283 66215
rect 95283 66181 95292 66215
rect 95240 66172 95292 66181
rect 95332 66104 95384 66156
rect 95884 66172 95936 66224
rect 96712 66172 96764 66224
rect 96068 66104 96120 66156
rect 100760 66172 100812 66224
rect 89260 65968 89312 66020
rect 95884 65968 95936 66020
rect 88248 65900 88300 65952
rect 90732 65900 90784 65952
rect 94412 65943 94464 65952
rect 94412 65909 94421 65943
rect 94421 65909 94455 65943
rect 94455 65909 94464 65943
rect 94412 65900 94464 65909
rect 94964 65900 95016 65952
rect 95792 65900 95844 65952
rect 95976 65943 96028 65952
rect 95976 65909 95985 65943
rect 95985 65909 96019 65943
rect 96019 65909 96028 65943
rect 95976 65900 96028 65909
rect 97540 66147 97592 66156
rect 97540 66113 97549 66147
rect 97549 66113 97583 66147
rect 97583 66113 97592 66147
rect 97540 66104 97592 66113
rect 98552 66147 98604 66156
rect 98552 66113 98561 66147
rect 98561 66113 98595 66147
rect 98595 66113 98604 66147
rect 98552 66104 98604 66113
rect 98736 66104 98788 66156
rect 99380 66104 99432 66156
rect 99656 66104 99708 66156
rect 100852 66104 100904 66156
rect 97908 66036 97960 66088
rect 99932 66036 99984 66088
rect 100300 66079 100352 66088
rect 100300 66045 100309 66079
rect 100309 66045 100343 66079
rect 100343 66045 100352 66079
rect 100300 66036 100352 66045
rect 101312 66215 101364 66224
rect 101312 66181 101321 66215
rect 101321 66181 101355 66215
rect 101355 66181 101364 66215
rect 101312 66172 101364 66181
rect 101956 66104 102008 66156
rect 102784 66172 102836 66224
rect 102876 66104 102928 66156
rect 103704 66104 103756 66156
rect 104624 66104 104676 66156
rect 103520 66036 103572 66088
rect 96896 65968 96948 66020
rect 99380 65968 99432 66020
rect 99748 65968 99800 66020
rect 103704 65968 103756 66020
rect 100576 65900 100628 65952
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 96374 65798 96426 65850
rect 96438 65798 96490 65850
rect 96502 65798 96554 65850
rect 96566 65798 96618 65850
rect 96630 65798 96682 65850
rect 105922 65798 105974 65850
rect 105986 65798 106038 65850
rect 106050 65798 106102 65850
rect 106114 65798 106166 65850
rect 106178 65798 106230 65850
rect 94136 65696 94188 65748
rect 103612 65696 103664 65748
rect 94872 65628 94924 65680
rect 102232 65628 102284 65680
rect 4874 65254 4926 65306
rect 4938 65254 4990 65306
rect 5002 65254 5054 65306
rect 5066 65254 5118 65306
rect 5130 65254 5182 65306
rect 106658 65254 106710 65306
rect 106722 65254 106774 65306
rect 106786 65254 106838 65306
rect 106850 65254 106902 65306
rect 106914 65254 106966 65306
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 105922 64710 105974 64762
rect 105986 64710 106038 64762
rect 106050 64710 106102 64762
rect 106114 64710 106166 64762
rect 106178 64710 106230 64762
rect 4874 64166 4926 64218
rect 4938 64166 4990 64218
rect 5002 64166 5054 64218
rect 5066 64166 5118 64218
rect 5130 64166 5182 64218
rect 106658 64166 106710 64218
rect 106722 64166 106774 64218
rect 106786 64166 106838 64218
rect 106850 64166 106902 64218
rect 106914 64166 106966 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 105922 63622 105974 63674
rect 105986 63622 106038 63674
rect 106050 63622 106102 63674
rect 106114 63622 106166 63674
rect 106178 63622 106230 63674
rect 4874 63078 4926 63130
rect 4938 63078 4990 63130
rect 5002 63078 5054 63130
rect 5066 63078 5118 63130
rect 5130 63078 5182 63130
rect 106658 63078 106710 63130
rect 106722 63078 106774 63130
rect 106786 63078 106838 63130
rect 106850 63078 106902 63130
rect 106914 63078 106966 63130
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 105922 62534 105974 62586
rect 105986 62534 106038 62586
rect 106050 62534 106102 62586
rect 106114 62534 106166 62586
rect 106178 62534 106230 62586
rect 4874 61990 4926 62042
rect 4938 61990 4990 62042
rect 5002 61990 5054 62042
rect 5066 61990 5118 62042
rect 5130 61990 5182 62042
rect 106658 61990 106710 62042
rect 106722 61990 106774 62042
rect 106786 61990 106838 62042
rect 106850 61990 106902 62042
rect 106914 61990 106966 62042
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 105922 61446 105974 61498
rect 105986 61446 106038 61498
rect 106050 61446 106102 61498
rect 106114 61446 106166 61498
rect 106178 61446 106230 61498
rect 4874 60902 4926 60954
rect 4938 60902 4990 60954
rect 5002 60902 5054 60954
rect 5066 60902 5118 60954
rect 5130 60902 5182 60954
rect 106658 60902 106710 60954
rect 106722 60902 106774 60954
rect 106786 60902 106838 60954
rect 106850 60902 106902 60954
rect 106914 60902 106966 60954
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 105922 60358 105974 60410
rect 105986 60358 106038 60410
rect 106050 60358 106102 60410
rect 106114 60358 106166 60410
rect 106178 60358 106230 60410
rect 104348 60095 104400 60104
rect 104348 60061 104357 60095
rect 104357 60061 104391 60095
rect 104391 60061 104400 60095
rect 104348 60052 104400 60061
rect 4874 59814 4926 59866
rect 4938 59814 4990 59866
rect 5002 59814 5054 59866
rect 5066 59814 5118 59866
rect 5130 59814 5182 59866
rect 106658 59814 106710 59866
rect 106722 59814 106774 59866
rect 106786 59814 106838 59866
rect 106850 59814 106902 59866
rect 106914 59814 106966 59866
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 105922 59270 105974 59322
rect 105986 59270 106038 59322
rect 106050 59270 106102 59322
rect 106114 59270 106166 59322
rect 106178 59270 106230 59322
rect 4874 58726 4926 58778
rect 4938 58726 4990 58778
rect 5002 58726 5054 58778
rect 5066 58726 5118 58778
rect 5130 58726 5182 58778
rect 106658 58726 106710 58778
rect 106722 58726 106774 58778
rect 106786 58726 106838 58778
rect 106850 58726 106902 58778
rect 106914 58726 106966 58778
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 105922 58182 105974 58234
rect 105986 58182 106038 58234
rect 106050 58182 106102 58234
rect 106114 58182 106166 58234
rect 106178 58182 106230 58234
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 106658 57638 106710 57690
rect 106722 57638 106774 57690
rect 106786 57638 106838 57690
rect 106850 57638 106902 57690
rect 106914 57638 106966 57690
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 105922 57094 105974 57146
rect 105986 57094 106038 57146
rect 106050 57094 106102 57146
rect 106114 57094 106166 57146
rect 106178 57094 106230 57146
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 106658 56550 106710 56602
rect 106722 56550 106774 56602
rect 106786 56550 106838 56602
rect 106850 56550 106902 56602
rect 106914 56550 106966 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 105922 56006 105974 56058
rect 105986 56006 106038 56058
rect 106050 56006 106102 56058
rect 106114 56006 106166 56058
rect 106178 56006 106230 56058
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 106658 55462 106710 55514
rect 106722 55462 106774 55514
rect 106786 55462 106838 55514
rect 106850 55462 106902 55514
rect 106914 55462 106966 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 105922 54918 105974 54970
rect 105986 54918 106038 54970
rect 106050 54918 106102 54970
rect 106114 54918 106166 54970
rect 106178 54918 106230 54970
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 106658 54374 106710 54426
rect 106722 54374 106774 54426
rect 106786 54374 106838 54426
rect 106850 54374 106902 54426
rect 106914 54374 106966 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 105922 53830 105974 53882
rect 105986 53830 106038 53882
rect 106050 53830 106102 53882
rect 106114 53830 106166 53882
rect 106178 53830 106230 53882
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 106658 53286 106710 53338
rect 106722 53286 106774 53338
rect 106786 53286 106838 53338
rect 106850 53286 106902 53338
rect 106914 53286 106966 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 105922 52742 105974 52794
rect 105986 52742 106038 52794
rect 106050 52742 106102 52794
rect 106114 52742 106166 52794
rect 106178 52742 106230 52794
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 106658 52198 106710 52250
rect 106722 52198 106774 52250
rect 106786 52198 106838 52250
rect 106850 52198 106902 52250
rect 106914 52198 106966 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 105922 51654 105974 51706
rect 105986 51654 106038 51706
rect 106050 51654 106102 51706
rect 106114 51654 106166 51706
rect 106178 51654 106230 51706
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 106658 51110 106710 51162
rect 106722 51110 106774 51162
rect 106786 51110 106838 51162
rect 106850 51110 106902 51162
rect 106914 51110 106966 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 105922 50566 105974 50618
rect 105986 50566 106038 50618
rect 106050 50566 106102 50618
rect 106114 50566 106166 50618
rect 106178 50566 106230 50618
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 106658 50022 106710 50074
rect 106722 50022 106774 50074
rect 106786 50022 106838 50074
rect 106850 50022 106902 50074
rect 106914 50022 106966 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 105922 49478 105974 49530
rect 105986 49478 106038 49530
rect 106050 49478 106102 49530
rect 106114 49478 106166 49530
rect 106178 49478 106230 49530
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 106658 48934 106710 48986
rect 106722 48934 106774 48986
rect 106786 48934 106838 48986
rect 106850 48934 106902 48986
rect 106914 48934 106966 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 105922 48390 105974 48442
rect 105986 48390 106038 48442
rect 106050 48390 106102 48442
rect 106114 48390 106166 48442
rect 106178 48390 106230 48442
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 106658 47846 106710 47898
rect 106722 47846 106774 47898
rect 106786 47846 106838 47898
rect 106850 47846 106902 47898
rect 106914 47846 106966 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 105922 47302 105974 47354
rect 105986 47302 106038 47354
rect 106050 47302 106102 47354
rect 106114 47302 106166 47354
rect 106178 47302 106230 47354
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 106658 46758 106710 46810
rect 106722 46758 106774 46810
rect 106786 46758 106838 46810
rect 106850 46758 106902 46810
rect 106914 46758 106966 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 105922 46214 105974 46266
rect 105986 46214 106038 46266
rect 106050 46214 106102 46266
rect 106114 46214 106166 46266
rect 106178 46214 106230 46266
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 106658 45670 106710 45722
rect 106722 45670 106774 45722
rect 106786 45670 106838 45722
rect 106850 45670 106902 45722
rect 106914 45670 106966 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 105922 45126 105974 45178
rect 105986 45126 106038 45178
rect 106050 45126 106102 45178
rect 106114 45126 106166 45178
rect 106178 45126 106230 45178
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 106658 44582 106710 44634
rect 106722 44582 106774 44634
rect 106786 44582 106838 44634
rect 106850 44582 106902 44634
rect 106914 44582 106966 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 105922 44038 105974 44090
rect 105986 44038 106038 44090
rect 106050 44038 106102 44090
rect 106114 44038 106166 44090
rect 106178 44038 106230 44090
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 106658 43494 106710 43546
rect 106722 43494 106774 43546
rect 106786 43494 106838 43546
rect 106850 43494 106902 43546
rect 106914 43494 106966 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 105922 42950 105974 43002
rect 105986 42950 106038 43002
rect 106050 42950 106102 43002
rect 106114 42950 106166 43002
rect 106178 42950 106230 43002
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 106658 42406 106710 42458
rect 106722 42406 106774 42458
rect 106786 42406 106838 42458
rect 106850 42406 106902 42458
rect 106914 42406 106966 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 105922 41862 105974 41914
rect 105986 41862 106038 41914
rect 106050 41862 106102 41914
rect 106114 41862 106166 41914
rect 106178 41862 106230 41914
rect 7564 41463 7616 41472
rect 7564 41429 7573 41463
rect 7573 41429 7607 41463
rect 7607 41429 7616 41463
rect 7564 41420 7616 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 106658 41318 106710 41370
rect 106722 41318 106774 41370
rect 106786 41318 106838 41370
rect 106850 41318 106902 41370
rect 106914 41318 106966 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 105922 40774 105974 40826
rect 105986 40774 106038 40826
rect 106050 40774 106102 40826
rect 106114 40774 106166 40826
rect 106178 40774 106230 40826
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 106658 40230 106710 40282
rect 106722 40230 106774 40282
rect 106786 40230 106838 40282
rect 106850 40230 106902 40282
rect 106914 40230 106966 40282
rect 3424 39992 3476 40044
rect 7564 39992 7616 40044
rect 7288 39788 7340 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 105922 39686 105974 39738
rect 105986 39686 106038 39738
rect 106050 39686 106102 39738
rect 106114 39686 106166 39738
rect 106178 39686 106230 39738
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 106658 39142 106710 39194
rect 106722 39142 106774 39194
rect 106786 39142 106838 39194
rect 106850 39142 106902 39194
rect 106914 39142 106966 39194
rect 7564 38743 7616 38752
rect 7564 38709 7573 38743
rect 7573 38709 7607 38743
rect 7607 38709 7616 38743
rect 7564 38700 7616 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 105922 38598 105974 38650
rect 105986 38598 106038 38650
rect 106050 38598 106102 38650
rect 106114 38598 106166 38650
rect 106178 38598 106230 38650
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 106658 38054 106710 38106
rect 106722 38054 106774 38106
rect 106786 38054 106838 38106
rect 106850 38054 106902 38106
rect 106914 38054 106966 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 105922 37510 105974 37562
rect 105986 37510 106038 37562
rect 106050 37510 106102 37562
rect 106114 37510 106166 37562
rect 106178 37510 106230 37562
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 106658 36966 106710 37018
rect 106722 36966 106774 37018
rect 106786 36966 106838 37018
rect 106850 36966 106902 37018
rect 106914 36966 106966 37018
rect 7564 36635 7616 36644
rect 7564 36601 7573 36635
rect 7573 36601 7607 36635
rect 7607 36601 7616 36635
rect 7564 36592 7616 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 105922 36422 105974 36474
rect 105986 36422 106038 36474
rect 106050 36422 106102 36474
rect 106114 36422 106166 36474
rect 106178 36422 106230 36474
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 106658 35878 106710 35930
rect 106722 35878 106774 35930
rect 106786 35878 106838 35930
rect 106850 35878 106902 35930
rect 106914 35878 106966 35930
rect 7472 35479 7524 35488
rect 7472 35445 7481 35479
rect 7481 35445 7515 35479
rect 7515 35445 7524 35479
rect 7472 35436 7524 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 105922 35334 105974 35386
rect 105986 35334 106038 35386
rect 106050 35334 106102 35386
rect 106114 35334 106166 35386
rect 106178 35334 106230 35386
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 106658 34790 106710 34842
rect 106722 34790 106774 34842
rect 106786 34790 106838 34842
rect 106850 34790 106902 34842
rect 106914 34790 106966 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 105922 34246 105974 34298
rect 105986 34246 106038 34298
rect 106050 34246 106102 34298
rect 106114 34246 106166 34298
rect 106178 34246 106230 34298
rect 7564 33915 7616 33924
rect 7564 33881 7573 33915
rect 7573 33881 7607 33915
rect 7607 33881 7616 33915
rect 7564 33872 7616 33881
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 106658 33702 106710 33754
rect 106722 33702 106774 33754
rect 106786 33702 106838 33754
rect 106850 33702 106902 33754
rect 106914 33702 106966 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 105922 33158 105974 33210
rect 105986 33158 106038 33210
rect 106050 33158 106102 33210
rect 106114 33158 106166 33210
rect 106178 33158 106230 33210
rect 1584 33056 1636 33108
rect 7564 33056 7616 33108
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 106658 32614 106710 32666
rect 106722 32614 106774 32666
rect 106786 32614 106838 32666
rect 106850 32614 106902 32666
rect 106914 32614 106966 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 105922 32070 105974 32122
rect 105986 32070 106038 32122
rect 106050 32070 106102 32122
rect 106114 32070 106166 32122
rect 106178 32070 106230 32122
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 106658 31526 106710 31578
rect 106722 31526 106774 31578
rect 106786 31526 106838 31578
rect 106850 31526 106902 31578
rect 106914 31526 106966 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 105922 30982 105974 31034
rect 105986 30982 106038 31034
rect 106050 30982 106102 31034
rect 106114 30982 106166 31034
rect 106178 30982 106230 31034
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 106658 30438 106710 30490
rect 106722 30438 106774 30490
rect 106786 30438 106838 30490
rect 106850 30438 106902 30490
rect 106914 30438 106966 30490
rect 1768 30268 1820 30320
rect 7472 30268 7524 30320
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 105922 29894 105974 29946
rect 105986 29894 106038 29946
rect 106050 29894 106102 29946
rect 106114 29894 106166 29946
rect 106178 29894 106230 29946
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 106658 29350 106710 29402
rect 106722 29350 106774 29402
rect 106786 29350 106838 29402
rect 106850 29350 106902 29402
rect 106914 29350 106966 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 105922 28806 105974 28858
rect 105986 28806 106038 28858
rect 106050 28806 106102 28858
rect 106114 28806 106166 28858
rect 106178 28806 106230 28858
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 106658 28262 106710 28314
rect 106722 28262 106774 28314
rect 106786 28262 106838 28314
rect 106850 28262 106902 28314
rect 106914 28262 106966 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 105922 27718 105974 27770
rect 105986 27718 106038 27770
rect 106050 27718 106102 27770
rect 106114 27718 106166 27770
rect 106178 27718 106230 27770
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 106658 27174 106710 27226
rect 106722 27174 106774 27226
rect 106786 27174 106838 27226
rect 106850 27174 106902 27226
rect 106914 27174 106966 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 105922 26630 105974 26682
rect 105986 26630 106038 26682
rect 106050 26630 106102 26682
rect 106114 26630 106166 26682
rect 106178 26630 106230 26682
rect 1860 26256 1912 26308
rect 7380 26256 7432 26308
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 106658 26086 106710 26138
rect 106722 26086 106774 26138
rect 106786 26086 106838 26138
rect 106850 26086 106902 26138
rect 106914 26086 106966 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 105922 25542 105974 25594
rect 105986 25542 106038 25594
rect 106050 25542 106102 25594
rect 106114 25542 106166 25594
rect 106178 25542 106230 25594
rect 102600 25100 102652 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 106658 24998 106710 25050
rect 106722 24998 106774 25050
rect 106786 24998 106838 25050
rect 106850 24998 106902 25050
rect 106914 24998 106966 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 105922 24454 105974 24506
rect 105986 24454 106038 24506
rect 106050 24454 106102 24506
rect 106114 24454 106166 24506
rect 106178 24454 106230 24506
rect 2044 24012 2096 24064
rect 7564 24012 7616 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 106658 23910 106710 23962
rect 106722 23910 106774 23962
rect 106786 23910 106838 23962
rect 106850 23910 106902 23962
rect 106914 23910 106966 23962
rect 102784 23468 102836 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 105922 23366 105974 23418
rect 105986 23366 106038 23418
rect 106050 23366 106102 23418
rect 106114 23366 106166 23418
rect 106178 23366 106230 23418
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 106658 22822 106710 22874
rect 106722 22822 106774 22874
rect 106786 22822 106838 22874
rect 106850 22822 106902 22874
rect 106914 22822 106966 22874
rect 102140 22720 102192 22772
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 105922 22278 105974 22330
rect 105986 22278 106038 22330
rect 106050 22278 106102 22330
rect 106114 22278 106166 22330
rect 106178 22278 106230 22330
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 106658 21734 106710 21786
rect 106722 21734 106774 21786
rect 106786 21734 106838 21786
rect 106850 21734 106902 21786
rect 106914 21734 106966 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 105922 21190 105974 21242
rect 105986 21190 106038 21242
rect 106050 21190 106102 21242
rect 106114 21190 106166 21242
rect 106178 21190 106230 21242
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 106658 20646 106710 20698
rect 106722 20646 106774 20698
rect 106786 20646 106838 20698
rect 106850 20646 106902 20698
rect 106914 20646 106966 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 105922 20102 105974 20154
rect 105986 20102 106038 20154
rect 106050 20102 106102 20154
rect 106114 20102 106166 20154
rect 106178 20102 106230 20154
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 106658 19558 106710 19610
rect 106722 19558 106774 19610
rect 106786 19558 106838 19610
rect 106850 19558 106902 19610
rect 106914 19558 106966 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 105922 19014 105974 19066
rect 105986 19014 106038 19066
rect 106050 19014 106102 19066
rect 106114 19014 106166 19066
rect 106178 19014 106230 19066
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 106658 18470 106710 18522
rect 106722 18470 106774 18522
rect 106786 18470 106838 18522
rect 106850 18470 106902 18522
rect 106914 18470 106966 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 105922 17926 105974 17978
rect 105986 17926 106038 17978
rect 106050 17926 106102 17978
rect 106114 17926 106166 17978
rect 106178 17926 106230 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 106658 17382 106710 17434
rect 106722 17382 106774 17434
rect 106786 17382 106838 17434
rect 106850 17382 106902 17434
rect 106914 17382 106966 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 105922 16838 105974 16890
rect 105986 16838 106038 16890
rect 106050 16838 106102 16890
rect 106114 16838 106166 16890
rect 106178 16838 106230 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 106658 16294 106710 16346
rect 106722 16294 106774 16346
rect 106786 16294 106838 16346
rect 106850 16294 106902 16346
rect 106914 16294 106966 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 105922 15750 105974 15802
rect 105986 15750 106038 15802
rect 106050 15750 106102 15802
rect 106114 15750 106166 15802
rect 106178 15750 106230 15802
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 106658 15206 106710 15258
rect 106722 15206 106774 15258
rect 106786 15206 106838 15258
rect 106850 15206 106902 15258
rect 106914 15206 106966 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 105922 14662 105974 14714
rect 105986 14662 106038 14714
rect 106050 14662 106102 14714
rect 106114 14662 106166 14714
rect 106178 14662 106230 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 106658 14118 106710 14170
rect 106722 14118 106774 14170
rect 106786 14118 106838 14170
rect 106850 14118 106902 14170
rect 106914 14118 106966 14170
rect 3424 14016 3476 14068
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 105922 13574 105974 13626
rect 105986 13574 106038 13626
rect 106050 13574 106102 13626
rect 106114 13574 106166 13626
rect 106178 13574 106230 13626
rect 2044 13472 2096 13524
rect 1308 13200 1360 13252
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 106658 13030 106710 13082
rect 106722 13030 106774 13082
rect 106786 13030 106838 13082
rect 106850 13030 106902 13082
rect 106914 13030 106966 13082
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 1492 12835 1544 12844
rect 1492 12801 1501 12835
rect 1501 12801 1535 12835
rect 1535 12801 1544 12835
rect 1492 12792 1544 12801
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 105922 12486 105974 12538
rect 105986 12486 106038 12538
rect 106050 12486 106102 12538
rect 106114 12486 106166 12538
rect 106178 12486 106230 12538
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 106658 11942 106710 11994
rect 106722 11942 106774 11994
rect 106786 11942 106838 11994
rect 106850 11942 106902 11994
rect 106914 11942 106966 11994
rect 1768 11883 1820 11892
rect 1768 11849 1777 11883
rect 1777 11849 1811 11883
rect 1811 11849 1820 11883
rect 1768 11840 1820 11849
rect 1216 11704 1268 11756
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 105922 11398 105974 11450
rect 105986 11398 106038 11450
rect 106050 11398 106102 11450
rect 106114 11398 106166 11450
rect 106178 11398 106230 11450
rect 7288 11296 7340 11348
rect 1492 11067 1544 11076
rect 1492 11033 1501 11067
rect 1501 11033 1535 11067
rect 1535 11033 1544 11067
rect 1492 11024 1544 11033
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 106658 10854 106710 10906
rect 106722 10854 106774 10906
rect 106786 10854 106838 10906
rect 106850 10854 106902 10906
rect 106914 10854 106966 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 1308 10616 1360 10668
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 105922 10310 105974 10362
rect 105986 10310 106038 10362
rect 106050 10310 106102 10362
rect 106114 10310 106166 10362
rect 106178 10310 106230 10362
rect 1492 9979 1544 9988
rect 1492 9945 1501 9979
rect 1501 9945 1535 9979
rect 1535 9945 1544 9979
rect 1492 9936 1544 9945
rect 29552 9868 29604 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 106658 9766 106710 9818
rect 106722 9766 106774 9818
rect 106786 9766 106838 9818
rect 106850 9766 106902 9818
rect 106914 9766 106966 9818
rect 9496 9596 9548 9648
rect 16028 9596 16080 9648
rect 9588 9528 9640 9580
rect 16120 9528 16172 9580
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 105922 9222 105974 9274
rect 105986 9222 106038 9274
rect 106050 9222 106102 9274
rect 106114 9222 106166 9274
rect 106178 9222 106230 9274
rect 90824 9052 90876 9104
rect 103980 9052 104032 9104
rect 90640 8984 90692 9036
rect 103704 8984 103756 9036
rect 90548 8916 90600 8968
rect 103612 8916 103664 8968
rect 1216 8848 1268 8900
rect 26700 8780 26752 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 106658 8678 106710 8730
rect 106722 8678 106774 8730
rect 106786 8678 106838 8730
rect 106850 8678 106902 8730
rect 106914 8678 106966 8730
rect 2044 8372 2096 8424
rect 24676 8304 24728 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 105922 8134 105974 8186
rect 105986 8134 106038 8186
rect 106050 8134 106102 8186
rect 106114 8134 106166 8186
rect 106178 8134 106230 8186
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 1308 7760 1360 7812
rect 30472 7692 30524 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 66314 7590 66366 7642
rect 66378 7590 66430 7642
rect 66442 7590 66494 7642
rect 66506 7590 66558 7642
rect 66570 7590 66622 7642
rect 97034 7590 97086 7642
rect 97098 7590 97150 7642
rect 97162 7590 97214 7642
rect 97226 7590 97278 7642
rect 97290 7590 97342 7642
rect 106658 7590 106710 7642
rect 106722 7590 106774 7642
rect 106786 7590 106838 7642
rect 106850 7590 106902 7642
rect 106914 7590 106966 7642
rect 16028 7488 16080 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 25780 7488 25832 7540
rect 26700 7488 26752 7540
rect 28172 7531 28224 7540
rect 28172 7497 28181 7531
rect 28181 7497 28215 7531
rect 28215 7497 28224 7531
rect 28172 7488 28224 7497
rect 29552 7531 29604 7540
rect 29552 7497 29561 7531
rect 29561 7497 29595 7531
rect 29595 7497 29604 7531
rect 29552 7488 29604 7497
rect 30472 7531 30524 7540
rect 30472 7497 30481 7531
rect 30481 7497 30515 7531
rect 30515 7497 30524 7531
rect 30472 7488 30524 7497
rect 90548 7531 90600 7540
rect 90548 7497 90557 7531
rect 90557 7497 90591 7531
rect 90591 7497 90600 7531
rect 90548 7488 90600 7497
rect 90640 7488 90692 7540
rect 90824 7488 90876 7540
rect 1308 7352 1360 7404
rect 28172 7216 28224 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 105922 7046 105974 7098
rect 105986 7046 106038 7098
rect 106050 7046 106102 7098
rect 106114 7046 106166 7098
rect 106178 7046 106230 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 66314 6502 66366 6554
rect 66378 6502 66430 6554
rect 66442 6502 66494 6554
rect 66506 6502 66558 6554
rect 66570 6502 66622 6554
rect 97034 6502 97086 6554
rect 97098 6502 97150 6554
rect 97162 6502 97214 6554
rect 97226 6502 97278 6554
rect 97290 6502 97342 6554
rect 1216 6264 1268 6316
rect 25872 6060 25924 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 7472 5856 7524 5908
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 66314 5414 66366 5466
rect 66378 5414 66430 5466
rect 66442 5414 66494 5466
rect 66506 5414 66558 5466
rect 66570 5414 66622 5466
rect 97034 5414 97086 5466
rect 97098 5414 97150 5466
rect 97162 5414 97214 5466
rect 97226 5414 97278 5466
rect 97290 5414 97342 5466
rect 1308 5176 1360 5228
rect 23480 4972 23532 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 66314 4326 66366 4378
rect 66378 4326 66430 4378
rect 66442 4326 66494 4378
rect 66506 4326 66558 4378
rect 66570 4326 66622 4378
rect 97034 4326 97086 4378
rect 97098 4326 97150 4378
rect 97162 4326 97214 4378
rect 97226 4326 97278 4378
rect 97290 4326 97342 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 66314 3238 66366 3290
rect 66378 3238 66430 3290
rect 66442 3238 66494 3290
rect 66506 3238 66558 3290
rect 66570 3238 66622 3290
rect 97034 3238 97086 3290
rect 97098 3238 97150 3290
rect 97162 3238 97214 3290
rect 97226 3238 97278 3290
rect 97290 3238 97342 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 31668 2635 31720 2644
rect 31668 2601 31677 2635
rect 31677 2601 31711 2635
rect 31711 2601 31720 2635
rect 31668 2592 31720 2601
rect 32956 2635 33008 2644
rect 32956 2601 32965 2635
rect 32965 2601 32999 2635
rect 32999 2601 33008 2635
rect 32956 2592 33008 2601
rect 34244 2635 34296 2644
rect 34244 2601 34253 2635
rect 34253 2601 34287 2635
rect 34287 2601 34296 2635
rect 34244 2592 34296 2601
rect 35440 2592 35492 2644
rect 36360 2635 36412 2644
rect 36360 2601 36369 2635
rect 36369 2601 36403 2635
rect 36403 2601 36412 2635
rect 36360 2592 36412 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 38752 2635 38804 2644
rect 38752 2601 38761 2635
rect 38761 2601 38795 2635
rect 38795 2601 38804 2635
rect 38752 2592 38804 2601
rect 39948 2592 40000 2644
rect 41328 2635 41380 2644
rect 41328 2601 41337 2635
rect 41337 2601 41371 2635
rect 41371 2601 41380 2635
rect 41328 2592 41380 2601
rect 42156 2635 42208 2644
rect 42156 2601 42165 2635
rect 42165 2601 42199 2635
rect 42199 2601 42208 2635
rect 42156 2592 42208 2601
rect 43444 2635 43496 2644
rect 43444 2601 43453 2635
rect 43453 2601 43487 2635
rect 43487 2601 43496 2635
rect 43444 2592 43496 2601
rect 31576 2295 31628 2304
rect 31576 2261 31585 2295
rect 31585 2261 31619 2295
rect 31619 2261 31628 2295
rect 31576 2252 31628 2261
rect 32864 2295 32916 2304
rect 32864 2261 32873 2295
rect 32873 2261 32907 2295
rect 32907 2261 32916 2295
rect 32864 2252 32916 2261
rect 34152 2295 34204 2304
rect 34152 2261 34161 2295
rect 34161 2261 34195 2295
rect 34195 2261 34204 2295
rect 34152 2252 34204 2261
rect 35440 2295 35492 2304
rect 35440 2261 35449 2295
rect 35449 2261 35483 2295
rect 35483 2261 35492 2295
rect 35440 2252 35492 2261
rect 36084 2295 36136 2304
rect 36084 2261 36093 2295
rect 36093 2261 36127 2295
rect 36127 2261 36136 2295
rect 36084 2252 36136 2261
rect 37372 2295 37424 2304
rect 37372 2261 37381 2295
rect 37381 2261 37415 2295
rect 37415 2261 37424 2295
rect 37372 2252 37424 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 39948 2295 40000 2304
rect 39948 2261 39957 2295
rect 39957 2261 39991 2295
rect 39991 2261 40000 2295
rect 39948 2252 40000 2261
rect 41236 2295 41288 2304
rect 41236 2261 41245 2295
rect 41245 2261 41279 2295
rect 41279 2261 41288 2295
rect 41236 2252 41288 2261
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 43168 2295 43220 2304
rect 43168 2261 43177 2295
rect 43177 2261 43211 2295
rect 43211 2261 43220 2295
rect 43168 2252 43220 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 66314 2150 66366 2202
rect 66378 2150 66430 2202
rect 66442 2150 66494 2202
rect 66506 2150 66558 2202
rect 66570 2150 66622 2202
rect 97034 2150 97086 2202
rect 97098 2150 97150 2202
rect 97162 2150 97214 2202
rect 97226 2150 97278 2202
rect 97290 2150 97342 2202
<< metal2 >>
rect 4214 147452 4522 147461
rect 4214 147450 4220 147452
rect 4276 147450 4300 147452
rect 4356 147450 4380 147452
rect 4436 147450 4460 147452
rect 4516 147450 4522 147452
rect 4276 147398 4278 147450
rect 4458 147398 4460 147450
rect 4214 147396 4220 147398
rect 4276 147396 4300 147398
rect 4356 147396 4380 147398
rect 4436 147396 4460 147398
rect 4516 147396 4522 147398
rect 4214 147387 4522 147396
rect 34934 147452 35242 147461
rect 34934 147450 34940 147452
rect 34996 147450 35020 147452
rect 35076 147450 35100 147452
rect 35156 147450 35180 147452
rect 35236 147450 35242 147452
rect 34996 147398 34998 147450
rect 35178 147398 35180 147450
rect 34934 147396 34940 147398
rect 34996 147396 35020 147398
rect 35076 147396 35100 147398
rect 35156 147396 35180 147398
rect 35236 147396 35242 147398
rect 34934 147387 35242 147396
rect 65654 147452 65962 147461
rect 65654 147450 65660 147452
rect 65716 147450 65740 147452
rect 65796 147450 65820 147452
rect 65876 147450 65900 147452
rect 65956 147450 65962 147452
rect 65716 147398 65718 147450
rect 65898 147398 65900 147450
rect 65654 147396 65660 147398
rect 65716 147396 65740 147398
rect 65796 147396 65820 147398
rect 65876 147396 65900 147398
rect 65956 147396 65962 147398
rect 65654 147387 65962 147396
rect 96374 147452 96682 147461
rect 96374 147450 96380 147452
rect 96436 147450 96460 147452
rect 96516 147450 96540 147452
rect 96596 147450 96620 147452
rect 96676 147450 96682 147452
rect 96436 147398 96438 147450
rect 96618 147398 96620 147450
rect 96374 147396 96380 147398
rect 96436 147396 96460 147398
rect 96516 147396 96540 147398
rect 96596 147396 96620 147398
rect 96676 147396 96682 147398
rect 96374 147387 96682 147396
rect 4874 146908 5182 146917
rect 4874 146906 4880 146908
rect 4936 146906 4960 146908
rect 5016 146906 5040 146908
rect 5096 146906 5120 146908
rect 5176 146906 5182 146908
rect 4936 146854 4938 146906
rect 5118 146854 5120 146906
rect 4874 146852 4880 146854
rect 4936 146852 4960 146854
rect 5016 146852 5040 146854
rect 5096 146852 5120 146854
rect 5176 146852 5182 146854
rect 4874 146843 5182 146852
rect 35594 146908 35902 146917
rect 35594 146906 35600 146908
rect 35656 146906 35680 146908
rect 35736 146906 35760 146908
rect 35816 146906 35840 146908
rect 35896 146906 35902 146908
rect 35656 146854 35658 146906
rect 35838 146854 35840 146906
rect 35594 146852 35600 146854
rect 35656 146852 35680 146854
rect 35736 146852 35760 146854
rect 35816 146852 35840 146854
rect 35896 146852 35902 146854
rect 35594 146843 35902 146852
rect 66314 146908 66622 146917
rect 66314 146906 66320 146908
rect 66376 146906 66400 146908
rect 66456 146906 66480 146908
rect 66536 146906 66560 146908
rect 66616 146906 66622 146908
rect 66376 146854 66378 146906
rect 66558 146854 66560 146906
rect 66314 146852 66320 146854
rect 66376 146852 66400 146854
rect 66456 146852 66480 146854
rect 66536 146852 66560 146854
rect 66616 146852 66622 146854
rect 66314 146843 66622 146852
rect 97034 146908 97342 146917
rect 97034 146906 97040 146908
rect 97096 146906 97120 146908
rect 97176 146906 97200 146908
rect 97256 146906 97280 146908
rect 97336 146906 97342 146908
rect 97096 146854 97098 146906
rect 97278 146854 97280 146906
rect 97034 146852 97040 146854
rect 97096 146852 97120 146854
rect 97176 146852 97200 146854
rect 97256 146852 97280 146854
rect 97336 146852 97342 146854
rect 97034 146843 97342 146852
rect 4214 146364 4522 146373
rect 4214 146362 4220 146364
rect 4276 146362 4300 146364
rect 4356 146362 4380 146364
rect 4436 146362 4460 146364
rect 4516 146362 4522 146364
rect 4276 146310 4278 146362
rect 4458 146310 4460 146362
rect 4214 146308 4220 146310
rect 4276 146308 4300 146310
rect 4356 146308 4380 146310
rect 4436 146308 4460 146310
rect 4516 146308 4522 146310
rect 4214 146299 4522 146308
rect 34934 146364 35242 146373
rect 34934 146362 34940 146364
rect 34996 146362 35020 146364
rect 35076 146362 35100 146364
rect 35156 146362 35180 146364
rect 35236 146362 35242 146364
rect 34996 146310 34998 146362
rect 35178 146310 35180 146362
rect 34934 146308 34940 146310
rect 34996 146308 35020 146310
rect 35076 146308 35100 146310
rect 35156 146308 35180 146310
rect 35236 146308 35242 146310
rect 34934 146299 35242 146308
rect 65654 146364 65962 146373
rect 65654 146362 65660 146364
rect 65716 146362 65740 146364
rect 65796 146362 65820 146364
rect 65876 146362 65900 146364
rect 65956 146362 65962 146364
rect 65716 146310 65718 146362
rect 65898 146310 65900 146362
rect 65654 146308 65660 146310
rect 65716 146308 65740 146310
rect 65796 146308 65820 146310
rect 65876 146308 65900 146310
rect 65956 146308 65962 146310
rect 65654 146299 65962 146308
rect 96374 146364 96682 146373
rect 96374 146362 96380 146364
rect 96436 146362 96460 146364
rect 96516 146362 96540 146364
rect 96596 146362 96620 146364
rect 96676 146362 96682 146364
rect 96436 146310 96438 146362
rect 96618 146310 96620 146362
rect 96374 146308 96380 146310
rect 96436 146308 96460 146310
rect 96516 146308 96540 146310
rect 96596 146308 96620 146310
rect 96676 146308 96682 146310
rect 96374 146299 96682 146308
rect 4874 145820 5182 145829
rect 4874 145818 4880 145820
rect 4936 145818 4960 145820
rect 5016 145818 5040 145820
rect 5096 145818 5120 145820
rect 5176 145818 5182 145820
rect 4936 145766 4938 145818
rect 5118 145766 5120 145818
rect 4874 145764 4880 145766
rect 4936 145764 4960 145766
rect 5016 145764 5040 145766
rect 5096 145764 5120 145766
rect 5176 145764 5182 145766
rect 4874 145755 5182 145764
rect 35594 145820 35902 145829
rect 35594 145818 35600 145820
rect 35656 145818 35680 145820
rect 35736 145818 35760 145820
rect 35816 145818 35840 145820
rect 35896 145818 35902 145820
rect 35656 145766 35658 145818
rect 35838 145766 35840 145818
rect 35594 145764 35600 145766
rect 35656 145764 35680 145766
rect 35736 145764 35760 145766
rect 35816 145764 35840 145766
rect 35896 145764 35902 145766
rect 35594 145755 35902 145764
rect 66314 145820 66622 145829
rect 66314 145818 66320 145820
rect 66376 145818 66400 145820
rect 66456 145818 66480 145820
rect 66536 145818 66560 145820
rect 66616 145818 66622 145820
rect 66376 145766 66378 145818
rect 66558 145766 66560 145818
rect 66314 145764 66320 145766
rect 66376 145764 66400 145766
rect 66456 145764 66480 145766
rect 66536 145764 66560 145766
rect 66616 145764 66622 145766
rect 66314 145755 66622 145764
rect 97034 145820 97342 145829
rect 97034 145818 97040 145820
rect 97096 145818 97120 145820
rect 97176 145818 97200 145820
rect 97256 145818 97280 145820
rect 97336 145818 97342 145820
rect 97096 145766 97098 145818
rect 97278 145766 97280 145818
rect 97034 145764 97040 145766
rect 97096 145764 97120 145766
rect 97176 145764 97200 145766
rect 97256 145764 97280 145766
rect 97336 145764 97342 145766
rect 97034 145755 97342 145764
rect 4214 145276 4522 145285
rect 4214 145274 4220 145276
rect 4276 145274 4300 145276
rect 4356 145274 4380 145276
rect 4436 145274 4460 145276
rect 4516 145274 4522 145276
rect 4276 145222 4278 145274
rect 4458 145222 4460 145274
rect 4214 145220 4220 145222
rect 4276 145220 4300 145222
rect 4356 145220 4380 145222
rect 4436 145220 4460 145222
rect 4516 145220 4522 145222
rect 4214 145211 4522 145220
rect 34934 145276 35242 145285
rect 34934 145274 34940 145276
rect 34996 145274 35020 145276
rect 35076 145274 35100 145276
rect 35156 145274 35180 145276
rect 35236 145274 35242 145276
rect 34996 145222 34998 145274
rect 35178 145222 35180 145274
rect 34934 145220 34940 145222
rect 34996 145220 35020 145222
rect 35076 145220 35100 145222
rect 35156 145220 35180 145222
rect 35236 145220 35242 145222
rect 34934 145211 35242 145220
rect 65654 145276 65962 145285
rect 65654 145274 65660 145276
rect 65716 145274 65740 145276
rect 65796 145274 65820 145276
rect 65876 145274 65900 145276
rect 65956 145274 65962 145276
rect 65716 145222 65718 145274
rect 65898 145222 65900 145274
rect 65654 145220 65660 145222
rect 65716 145220 65740 145222
rect 65796 145220 65820 145222
rect 65876 145220 65900 145222
rect 65956 145220 65962 145222
rect 65654 145211 65962 145220
rect 96374 145276 96682 145285
rect 96374 145274 96380 145276
rect 96436 145274 96460 145276
rect 96516 145274 96540 145276
rect 96596 145274 96620 145276
rect 96676 145274 96682 145276
rect 96436 145222 96438 145274
rect 96618 145222 96620 145274
rect 96374 145220 96380 145222
rect 96436 145220 96460 145222
rect 96516 145220 96540 145222
rect 96596 145220 96620 145222
rect 96676 145220 96682 145222
rect 96374 145211 96682 145220
rect 4874 144732 5182 144741
rect 4874 144730 4880 144732
rect 4936 144730 4960 144732
rect 5016 144730 5040 144732
rect 5096 144730 5120 144732
rect 5176 144730 5182 144732
rect 4936 144678 4938 144730
rect 5118 144678 5120 144730
rect 4874 144676 4880 144678
rect 4936 144676 4960 144678
rect 5016 144676 5040 144678
rect 5096 144676 5120 144678
rect 5176 144676 5182 144678
rect 4874 144667 5182 144676
rect 35594 144732 35902 144741
rect 35594 144730 35600 144732
rect 35656 144730 35680 144732
rect 35736 144730 35760 144732
rect 35816 144730 35840 144732
rect 35896 144730 35902 144732
rect 35656 144678 35658 144730
rect 35838 144678 35840 144730
rect 35594 144676 35600 144678
rect 35656 144676 35680 144678
rect 35736 144676 35760 144678
rect 35816 144676 35840 144678
rect 35896 144676 35902 144678
rect 35594 144667 35902 144676
rect 66314 144732 66622 144741
rect 66314 144730 66320 144732
rect 66376 144730 66400 144732
rect 66456 144730 66480 144732
rect 66536 144730 66560 144732
rect 66616 144730 66622 144732
rect 66376 144678 66378 144730
rect 66558 144678 66560 144730
rect 66314 144676 66320 144678
rect 66376 144676 66400 144678
rect 66456 144676 66480 144678
rect 66536 144676 66560 144678
rect 66616 144676 66622 144678
rect 66314 144667 66622 144676
rect 97034 144732 97342 144741
rect 97034 144730 97040 144732
rect 97096 144730 97120 144732
rect 97176 144730 97200 144732
rect 97256 144730 97280 144732
rect 97336 144730 97342 144732
rect 97096 144678 97098 144730
rect 97278 144678 97280 144730
rect 97034 144676 97040 144678
rect 97096 144676 97120 144678
rect 97176 144676 97200 144678
rect 97256 144676 97280 144678
rect 97336 144676 97342 144678
rect 97034 144667 97342 144676
rect 4214 144188 4522 144197
rect 4214 144186 4220 144188
rect 4276 144186 4300 144188
rect 4356 144186 4380 144188
rect 4436 144186 4460 144188
rect 4516 144186 4522 144188
rect 4276 144134 4278 144186
rect 4458 144134 4460 144186
rect 4214 144132 4220 144134
rect 4276 144132 4300 144134
rect 4356 144132 4380 144134
rect 4436 144132 4460 144134
rect 4516 144132 4522 144134
rect 4214 144123 4522 144132
rect 34934 144188 35242 144197
rect 34934 144186 34940 144188
rect 34996 144186 35020 144188
rect 35076 144186 35100 144188
rect 35156 144186 35180 144188
rect 35236 144186 35242 144188
rect 34996 144134 34998 144186
rect 35178 144134 35180 144186
rect 34934 144132 34940 144134
rect 34996 144132 35020 144134
rect 35076 144132 35100 144134
rect 35156 144132 35180 144134
rect 35236 144132 35242 144134
rect 34934 144123 35242 144132
rect 65654 144188 65962 144197
rect 65654 144186 65660 144188
rect 65716 144186 65740 144188
rect 65796 144186 65820 144188
rect 65876 144186 65900 144188
rect 65956 144186 65962 144188
rect 65716 144134 65718 144186
rect 65898 144134 65900 144186
rect 65654 144132 65660 144134
rect 65716 144132 65740 144134
rect 65796 144132 65820 144134
rect 65876 144132 65900 144134
rect 65956 144132 65962 144134
rect 65654 144123 65962 144132
rect 96374 144188 96682 144197
rect 96374 144186 96380 144188
rect 96436 144186 96460 144188
rect 96516 144186 96540 144188
rect 96596 144186 96620 144188
rect 96676 144186 96682 144188
rect 96436 144134 96438 144186
rect 96618 144134 96620 144186
rect 96374 144132 96380 144134
rect 96436 144132 96460 144134
rect 96516 144132 96540 144134
rect 96596 144132 96620 144134
rect 96676 144132 96682 144134
rect 96374 144123 96682 144132
rect 4874 143644 5182 143653
rect 4874 143642 4880 143644
rect 4936 143642 4960 143644
rect 5016 143642 5040 143644
rect 5096 143642 5120 143644
rect 5176 143642 5182 143644
rect 4936 143590 4938 143642
rect 5118 143590 5120 143642
rect 4874 143588 4880 143590
rect 4936 143588 4960 143590
rect 5016 143588 5040 143590
rect 5096 143588 5120 143590
rect 5176 143588 5182 143590
rect 4874 143579 5182 143588
rect 35594 143644 35902 143653
rect 35594 143642 35600 143644
rect 35656 143642 35680 143644
rect 35736 143642 35760 143644
rect 35816 143642 35840 143644
rect 35896 143642 35902 143644
rect 35656 143590 35658 143642
rect 35838 143590 35840 143642
rect 35594 143588 35600 143590
rect 35656 143588 35680 143590
rect 35736 143588 35760 143590
rect 35816 143588 35840 143590
rect 35896 143588 35902 143590
rect 35594 143579 35902 143588
rect 66314 143644 66622 143653
rect 66314 143642 66320 143644
rect 66376 143642 66400 143644
rect 66456 143642 66480 143644
rect 66536 143642 66560 143644
rect 66616 143642 66622 143644
rect 66376 143590 66378 143642
rect 66558 143590 66560 143642
rect 66314 143588 66320 143590
rect 66376 143588 66400 143590
rect 66456 143588 66480 143590
rect 66536 143588 66560 143590
rect 66616 143588 66622 143590
rect 66314 143579 66622 143588
rect 97034 143644 97342 143653
rect 97034 143642 97040 143644
rect 97096 143642 97120 143644
rect 97176 143642 97200 143644
rect 97256 143642 97280 143644
rect 97336 143642 97342 143644
rect 97096 143590 97098 143642
rect 97278 143590 97280 143642
rect 97034 143588 97040 143590
rect 97096 143588 97120 143590
rect 97176 143588 97200 143590
rect 97256 143588 97280 143590
rect 97336 143588 97342 143590
rect 97034 143579 97342 143588
rect 4214 143100 4522 143109
rect 4214 143098 4220 143100
rect 4276 143098 4300 143100
rect 4356 143098 4380 143100
rect 4436 143098 4460 143100
rect 4516 143098 4522 143100
rect 4276 143046 4278 143098
rect 4458 143046 4460 143098
rect 4214 143044 4220 143046
rect 4276 143044 4300 143046
rect 4356 143044 4380 143046
rect 4436 143044 4460 143046
rect 4516 143044 4522 143046
rect 4214 143035 4522 143044
rect 34934 143100 35242 143109
rect 34934 143098 34940 143100
rect 34996 143098 35020 143100
rect 35076 143098 35100 143100
rect 35156 143098 35180 143100
rect 35236 143098 35242 143100
rect 34996 143046 34998 143098
rect 35178 143046 35180 143098
rect 34934 143044 34940 143046
rect 34996 143044 35020 143046
rect 35076 143044 35100 143046
rect 35156 143044 35180 143046
rect 35236 143044 35242 143046
rect 34934 143035 35242 143044
rect 65654 143100 65962 143109
rect 65654 143098 65660 143100
rect 65716 143098 65740 143100
rect 65796 143098 65820 143100
rect 65876 143098 65900 143100
rect 65956 143098 65962 143100
rect 65716 143046 65718 143098
rect 65898 143046 65900 143098
rect 65654 143044 65660 143046
rect 65716 143044 65740 143046
rect 65796 143044 65820 143046
rect 65876 143044 65900 143046
rect 65956 143044 65962 143046
rect 65654 143035 65962 143044
rect 96374 143100 96682 143109
rect 96374 143098 96380 143100
rect 96436 143098 96460 143100
rect 96516 143098 96540 143100
rect 96596 143098 96620 143100
rect 96676 143098 96682 143100
rect 96436 143046 96438 143098
rect 96618 143046 96620 143098
rect 96374 143044 96380 143046
rect 96436 143044 96460 143046
rect 96516 143044 96540 143046
rect 96596 143044 96620 143046
rect 96676 143044 96682 143046
rect 96374 143035 96682 143044
rect 4874 142556 5182 142565
rect 4874 142554 4880 142556
rect 4936 142554 4960 142556
rect 5016 142554 5040 142556
rect 5096 142554 5120 142556
rect 5176 142554 5182 142556
rect 4936 142502 4938 142554
rect 5118 142502 5120 142554
rect 4874 142500 4880 142502
rect 4936 142500 4960 142502
rect 5016 142500 5040 142502
rect 5096 142500 5120 142502
rect 5176 142500 5182 142502
rect 4874 142491 5182 142500
rect 35594 142556 35902 142565
rect 35594 142554 35600 142556
rect 35656 142554 35680 142556
rect 35736 142554 35760 142556
rect 35816 142554 35840 142556
rect 35896 142554 35902 142556
rect 35656 142502 35658 142554
rect 35838 142502 35840 142554
rect 35594 142500 35600 142502
rect 35656 142500 35680 142502
rect 35736 142500 35760 142502
rect 35816 142500 35840 142502
rect 35896 142500 35902 142502
rect 35594 142491 35902 142500
rect 66314 142556 66622 142565
rect 66314 142554 66320 142556
rect 66376 142554 66400 142556
rect 66456 142554 66480 142556
rect 66536 142554 66560 142556
rect 66616 142554 66622 142556
rect 66376 142502 66378 142554
rect 66558 142502 66560 142554
rect 66314 142500 66320 142502
rect 66376 142500 66400 142502
rect 66456 142500 66480 142502
rect 66536 142500 66560 142502
rect 66616 142500 66622 142502
rect 66314 142491 66622 142500
rect 97034 142556 97342 142565
rect 97034 142554 97040 142556
rect 97096 142554 97120 142556
rect 97176 142554 97200 142556
rect 97256 142554 97280 142556
rect 97336 142554 97342 142556
rect 97096 142502 97098 142554
rect 97278 142502 97280 142554
rect 97034 142500 97040 142502
rect 97096 142500 97120 142502
rect 97176 142500 97200 142502
rect 97256 142500 97280 142502
rect 97336 142500 97342 142502
rect 97034 142491 97342 142500
rect 4214 142012 4522 142021
rect 4214 142010 4220 142012
rect 4276 142010 4300 142012
rect 4356 142010 4380 142012
rect 4436 142010 4460 142012
rect 4516 142010 4522 142012
rect 4276 141958 4278 142010
rect 4458 141958 4460 142010
rect 4214 141956 4220 141958
rect 4276 141956 4300 141958
rect 4356 141956 4380 141958
rect 4436 141956 4460 141958
rect 4516 141956 4522 141958
rect 4214 141947 4522 141956
rect 34934 142012 35242 142021
rect 34934 142010 34940 142012
rect 34996 142010 35020 142012
rect 35076 142010 35100 142012
rect 35156 142010 35180 142012
rect 35236 142010 35242 142012
rect 34996 141958 34998 142010
rect 35178 141958 35180 142010
rect 34934 141956 34940 141958
rect 34996 141956 35020 141958
rect 35076 141956 35100 141958
rect 35156 141956 35180 141958
rect 35236 141956 35242 141958
rect 34934 141947 35242 141956
rect 65654 142012 65962 142021
rect 65654 142010 65660 142012
rect 65716 142010 65740 142012
rect 65796 142010 65820 142012
rect 65876 142010 65900 142012
rect 65956 142010 65962 142012
rect 65716 141958 65718 142010
rect 65898 141958 65900 142010
rect 65654 141956 65660 141958
rect 65716 141956 65740 141958
rect 65796 141956 65820 141958
rect 65876 141956 65900 141958
rect 65956 141956 65962 141958
rect 65654 141947 65962 141956
rect 96374 142012 96682 142021
rect 96374 142010 96380 142012
rect 96436 142010 96460 142012
rect 96516 142010 96540 142012
rect 96596 142010 96620 142012
rect 96676 142010 96682 142012
rect 96436 141958 96438 142010
rect 96618 141958 96620 142010
rect 96374 141956 96380 141958
rect 96436 141956 96460 141958
rect 96516 141956 96540 141958
rect 96596 141956 96620 141958
rect 96676 141956 96682 141958
rect 96374 141947 96682 141956
rect 4874 141468 5182 141477
rect 4874 141466 4880 141468
rect 4936 141466 4960 141468
rect 5016 141466 5040 141468
rect 5096 141466 5120 141468
rect 5176 141466 5182 141468
rect 4936 141414 4938 141466
rect 5118 141414 5120 141466
rect 4874 141412 4880 141414
rect 4936 141412 4960 141414
rect 5016 141412 5040 141414
rect 5096 141412 5120 141414
rect 5176 141412 5182 141414
rect 4874 141403 5182 141412
rect 35594 141468 35902 141477
rect 35594 141466 35600 141468
rect 35656 141466 35680 141468
rect 35736 141466 35760 141468
rect 35816 141466 35840 141468
rect 35896 141466 35902 141468
rect 35656 141414 35658 141466
rect 35838 141414 35840 141466
rect 35594 141412 35600 141414
rect 35656 141412 35680 141414
rect 35736 141412 35760 141414
rect 35816 141412 35840 141414
rect 35896 141412 35902 141414
rect 35594 141403 35902 141412
rect 66314 141468 66622 141477
rect 66314 141466 66320 141468
rect 66376 141466 66400 141468
rect 66456 141466 66480 141468
rect 66536 141466 66560 141468
rect 66616 141466 66622 141468
rect 66376 141414 66378 141466
rect 66558 141414 66560 141466
rect 66314 141412 66320 141414
rect 66376 141412 66400 141414
rect 66456 141412 66480 141414
rect 66536 141412 66560 141414
rect 66616 141412 66622 141414
rect 66314 141403 66622 141412
rect 97034 141468 97342 141477
rect 97034 141466 97040 141468
rect 97096 141466 97120 141468
rect 97176 141466 97200 141468
rect 97256 141466 97280 141468
rect 97336 141466 97342 141468
rect 97096 141414 97098 141466
rect 97278 141414 97280 141466
rect 97034 141412 97040 141414
rect 97096 141412 97120 141414
rect 97176 141412 97200 141414
rect 97256 141412 97280 141414
rect 97336 141412 97342 141414
rect 97034 141403 97342 141412
rect 4214 140924 4522 140933
rect 4214 140922 4220 140924
rect 4276 140922 4300 140924
rect 4356 140922 4380 140924
rect 4436 140922 4460 140924
rect 4516 140922 4522 140924
rect 4276 140870 4278 140922
rect 4458 140870 4460 140922
rect 4214 140868 4220 140870
rect 4276 140868 4300 140870
rect 4356 140868 4380 140870
rect 4436 140868 4460 140870
rect 4516 140868 4522 140870
rect 4214 140859 4522 140868
rect 34934 140924 35242 140933
rect 34934 140922 34940 140924
rect 34996 140922 35020 140924
rect 35076 140922 35100 140924
rect 35156 140922 35180 140924
rect 35236 140922 35242 140924
rect 34996 140870 34998 140922
rect 35178 140870 35180 140922
rect 34934 140868 34940 140870
rect 34996 140868 35020 140870
rect 35076 140868 35100 140870
rect 35156 140868 35180 140870
rect 35236 140868 35242 140870
rect 34934 140859 35242 140868
rect 65654 140924 65962 140933
rect 65654 140922 65660 140924
rect 65716 140922 65740 140924
rect 65796 140922 65820 140924
rect 65876 140922 65900 140924
rect 65956 140922 65962 140924
rect 65716 140870 65718 140922
rect 65898 140870 65900 140922
rect 65654 140868 65660 140870
rect 65716 140868 65740 140870
rect 65796 140868 65820 140870
rect 65876 140868 65900 140870
rect 65956 140868 65962 140870
rect 65654 140859 65962 140868
rect 96374 140924 96682 140933
rect 96374 140922 96380 140924
rect 96436 140922 96460 140924
rect 96516 140922 96540 140924
rect 96596 140922 96620 140924
rect 96676 140922 96682 140924
rect 96436 140870 96438 140922
rect 96618 140870 96620 140922
rect 96374 140868 96380 140870
rect 96436 140868 96460 140870
rect 96516 140868 96540 140870
rect 96596 140868 96620 140870
rect 96676 140868 96682 140870
rect 96374 140859 96682 140868
rect 4874 140380 5182 140389
rect 4874 140378 4880 140380
rect 4936 140378 4960 140380
rect 5016 140378 5040 140380
rect 5096 140378 5120 140380
rect 5176 140378 5182 140380
rect 4936 140326 4938 140378
rect 5118 140326 5120 140378
rect 4874 140324 4880 140326
rect 4936 140324 4960 140326
rect 5016 140324 5040 140326
rect 5096 140324 5120 140326
rect 5176 140324 5182 140326
rect 4874 140315 5182 140324
rect 35594 140380 35902 140389
rect 35594 140378 35600 140380
rect 35656 140378 35680 140380
rect 35736 140378 35760 140380
rect 35816 140378 35840 140380
rect 35896 140378 35902 140380
rect 35656 140326 35658 140378
rect 35838 140326 35840 140378
rect 35594 140324 35600 140326
rect 35656 140324 35680 140326
rect 35736 140324 35760 140326
rect 35816 140324 35840 140326
rect 35896 140324 35902 140326
rect 35594 140315 35902 140324
rect 66314 140380 66622 140389
rect 66314 140378 66320 140380
rect 66376 140378 66400 140380
rect 66456 140378 66480 140380
rect 66536 140378 66560 140380
rect 66616 140378 66622 140380
rect 66376 140326 66378 140378
rect 66558 140326 66560 140378
rect 66314 140324 66320 140326
rect 66376 140324 66400 140326
rect 66456 140324 66480 140326
rect 66536 140324 66560 140326
rect 66616 140324 66622 140326
rect 66314 140315 66622 140324
rect 97034 140380 97342 140389
rect 97034 140378 97040 140380
rect 97096 140378 97120 140380
rect 97176 140378 97200 140380
rect 97256 140378 97280 140380
rect 97336 140378 97342 140380
rect 97096 140326 97098 140378
rect 97278 140326 97280 140378
rect 97034 140324 97040 140326
rect 97096 140324 97120 140326
rect 97176 140324 97200 140326
rect 97256 140324 97280 140326
rect 97336 140324 97342 140326
rect 97034 140315 97342 140324
rect 4214 139836 4522 139845
rect 4214 139834 4220 139836
rect 4276 139834 4300 139836
rect 4356 139834 4380 139836
rect 4436 139834 4460 139836
rect 4516 139834 4522 139836
rect 4276 139782 4278 139834
rect 4458 139782 4460 139834
rect 4214 139780 4220 139782
rect 4276 139780 4300 139782
rect 4356 139780 4380 139782
rect 4436 139780 4460 139782
rect 4516 139780 4522 139782
rect 4214 139771 4522 139780
rect 34934 139836 35242 139845
rect 34934 139834 34940 139836
rect 34996 139834 35020 139836
rect 35076 139834 35100 139836
rect 35156 139834 35180 139836
rect 35236 139834 35242 139836
rect 34996 139782 34998 139834
rect 35178 139782 35180 139834
rect 34934 139780 34940 139782
rect 34996 139780 35020 139782
rect 35076 139780 35100 139782
rect 35156 139780 35180 139782
rect 35236 139780 35242 139782
rect 34934 139771 35242 139780
rect 65654 139836 65962 139845
rect 65654 139834 65660 139836
rect 65716 139834 65740 139836
rect 65796 139834 65820 139836
rect 65876 139834 65900 139836
rect 65956 139834 65962 139836
rect 65716 139782 65718 139834
rect 65898 139782 65900 139834
rect 65654 139780 65660 139782
rect 65716 139780 65740 139782
rect 65796 139780 65820 139782
rect 65876 139780 65900 139782
rect 65956 139780 65962 139782
rect 65654 139771 65962 139780
rect 96374 139836 96682 139845
rect 96374 139834 96380 139836
rect 96436 139834 96460 139836
rect 96516 139834 96540 139836
rect 96596 139834 96620 139836
rect 96676 139834 96682 139836
rect 96436 139782 96438 139834
rect 96618 139782 96620 139834
rect 96374 139780 96380 139782
rect 96436 139780 96460 139782
rect 96516 139780 96540 139782
rect 96596 139780 96620 139782
rect 96676 139780 96682 139782
rect 96374 139771 96682 139780
rect 4874 139292 5182 139301
rect 4874 139290 4880 139292
rect 4936 139290 4960 139292
rect 5016 139290 5040 139292
rect 5096 139290 5120 139292
rect 5176 139290 5182 139292
rect 4936 139238 4938 139290
rect 5118 139238 5120 139290
rect 4874 139236 4880 139238
rect 4936 139236 4960 139238
rect 5016 139236 5040 139238
rect 5096 139236 5120 139238
rect 5176 139236 5182 139238
rect 4874 139227 5182 139236
rect 35594 139292 35902 139301
rect 35594 139290 35600 139292
rect 35656 139290 35680 139292
rect 35736 139290 35760 139292
rect 35816 139290 35840 139292
rect 35896 139290 35902 139292
rect 35656 139238 35658 139290
rect 35838 139238 35840 139290
rect 35594 139236 35600 139238
rect 35656 139236 35680 139238
rect 35736 139236 35760 139238
rect 35816 139236 35840 139238
rect 35896 139236 35902 139238
rect 35594 139227 35902 139236
rect 66314 139292 66622 139301
rect 66314 139290 66320 139292
rect 66376 139290 66400 139292
rect 66456 139290 66480 139292
rect 66536 139290 66560 139292
rect 66616 139290 66622 139292
rect 66376 139238 66378 139290
rect 66558 139238 66560 139290
rect 66314 139236 66320 139238
rect 66376 139236 66400 139238
rect 66456 139236 66480 139238
rect 66536 139236 66560 139238
rect 66616 139236 66622 139238
rect 66314 139227 66622 139236
rect 97034 139292 97342 139301
rect 97034 139290 97040 139292
rect 97096 139290 97120 139292
rect 97176 139290 97200 139292
rect 97256 139290 97280 139292
rect 97336 139290 97342 139292
rect 97096 139238 97098 139290
rect 97278 139238 97280 139290
rect 97034 139236 97040 139238
rect 97096 139236 97120 139238
rect 97176 139236 97200 139238
rect 97256 139236 97280 139238
rect 97336 139236 97342 139238
rect 97034 139227 97342 139236
rect 4214 138748 4522 138757
rect 4214 138746 4220 138748
rect 4276 138746 4300 138748
rect 4356 138746 4380 138748
rect 4436 138746 4460 138748
rect 4516 138746 4522 138748
rect 4276 138694 4278 138746
rect 4458 138694 4460 138746
rect 4214 138692 4220 138694
rect 4276 138692 4300 138694
rect 4356 138692 4380 138694
rect 4436 138692 4460 138694
rect 4516 138692 4522 138694
rect 4214 138683 4522 138692
rect 34934 138748 35242 138757
rect 34934 138746 34940 138748
rect 34996 138746 35020 138748
rect 35076 138746 35100 138748
rect 35156 138746 35180 138748
rect 35236 138746 35242 138748
rect 34996 138694 34998 138746
rect 35178 138694 35180 138746
rect 34934 138692 34940 138694
rect 34996 138692 35020 138694
rect 35076 138692 35100 138694
rect 35156 138692 35180 138694
rect 35236 138692 35242 138694
rect 34934 138683 35242 138692
rect 65654 138748 65962 138757
rect 65654 138746 65660 138748
rect 65716 138746 65740 138748
rect 65796 138746 65820 138748
rect 65876 138746 65900 138748
rect 65956 138746 65962 138748
rect 65716 138694 65718 138746
rect 65898 138694 65900 138746
rect 65654 138692 65660 138694
rect 65716 138692 65740 138694
rect 65796 138692 65820 138694
rect 65876 138692 65900 138694
rect 65956 138692 65962 138694
rect 65654 138683 65962 138692
rect 96374 138748 96682 138757
rect 96374 138746 96380 138748
rect 96436 138746 96460 138748
rect 96516 138746 96540 138748
rect 96596 138746 96620 138748
rect 96676 138746 96682 138748
rect 96436 138694 96438 138746
rect 96618 138694 96620 138746
rect 96374 138692 96380 138694
rect 96436 138692 96460 138694
rect 96516 138692 96540 138694
rect 96596 138692 96620 138694
rect 96676 138692 96682 138694
rect 96374 138683 96682 138692
rect 4874 138204 5182 138213
rect 4874 138202 4880 138204
rect 4936 138202 4960 138204
rect 5016 138202 5040 138204
rect 5096 138202 5120 138204
rect 5176 138202 5182 138204
rect 4936 138150 4938 138202
rect 5118 138150 5120 138202
rect 4874 138148 4880 138150
rect 4936 138148 4960 138150
rect 5016 138148 5040 138150
rect 5096 138148 5120 138150
rect 5176 138148 5182 138150
rect 4874 138139 5182 138148
rect 35594 138204 35902 138213
rect 35594 138202 35600 138204
rect 35656 138202 35680 138204
rect 35736 138202 35760 138204
rect 35816 138202 35840 138204
rect 35896 138202 35902 138204
rect 35656 138150 35658 138202
rect 35838 138150 35840 138202
rect 35594 138148 35600 138150
rect 35656 138148 35680 138150
rect 35736 138148 35760 138150
rect 35816 138148 35840 138150
rect 35896 138148 35902 138150
rect 35594 138139 35902 138148
rect 66314 138204 66622 138213
rect 66314 138202 66320 138204
rect 66376 138202 66400 138204
rect 66456 138202 66480 138204
rect 66536 138202 66560 138204
rect 66616 138202 66622 138204
rect 66376 138150 66378 138202
rect 66558 138150 66560 138202
rect 66314 138148 66320 138150
rect 66376 138148 66400 138150
rect 66456 138148 66480 138150
rect 66536 138148 66560 138150
rect 66616 138148 66622 138150
rect 66314 138139 66622 138148
rect 97034 138204 97342 138213
rect 97034 138202 97040 138204
rect 97096 138202 97120 138204
rect 97176 138202 97200 138204
rect 97256 138202 97280 138204
rect 97336 138202 97342 138204
rect 97096 138150 97098 138202
rect 97278 138150 97280 138202
rect 97034 138148 97040 138150
rect 97096 138148 97120 138150
rect 97176 138148 97200 138150
rect 97256 138148 97280 138150
rect 97336 138148 97342 138150
rect 97034 138139 97342 138148
rect 4214 137660 4522 137669
rect 4214 137658 4220 137660
rect 4276 137658 4300 137660
rect 4356 137658 4380 137660
rect 4436 137658 4460 137660
rect 4516 137658 4522 137660
rect 4276 137606 4278 137658
rect 4458 137606 4460 137658
rect 4214 137604 4220 137606
rect 4276 137604 4300 137606
rect 4356 137604 4380 137606
rect 4436 137604 4460 137606
rect 4516 137604 4522 137606
rect 4214 137595 4522 137604
rect 34934 137660 35242 137669
rect 34934 137658 34940 137660
rect 34996 137658 35020 137660
rect 35076 137658 35100 137660
rect 35156 137658 35180 137660
rect 35236 137658 35242 137660
rect 34996 137606 34998 137658
rect 35178 137606 35180 137658
rect 34934 137604 34940 137606
rect 34996 137604 35020 137606
rect 35076 137604 35100 137606
rect 35156 137604 35180 137606
rect 35236 137604 35242 137606
rect 34934 137595 35242 137604
rect 65654 137660 65962 137669
rect 65654 137658 65660 137660
rect 65716 137658 65740 137660
rect 65796 137658 65820 137660
rect 65876 137658 65900 137660
rect 65956 137658 65962 137660
rect 65716 137606 65718 137658
rect 65898 137606 65900 137658
rect 65654 137604 65660 137606
rect 65716 137604 65740 137606
rect 65796 137604 65820 137606
rect 65876 137604 65900 137606
rect 65956 137604 65962 137606
rect 65654 137595 65962 137604
rect 96374 137660 96682 137669
rect 96374 137658 96380 137660
rect 96436 137658 96460 137660
rect 96516 137658 96540 137660
rect 96596 137658 96620 137660
rect 96676 137658 96682 137660
rect 96436 137606 96438 137658
rect 96618 137606 96620 137658
rect 96374 137604 96380 137606
rect 96436 137604 96460 137606
rect 96516 137604 96540 137606
rect 96596 137604 96620 137606
rect 96676 137604 96682 137606
rect 96374 137595 96682 137604
rect 4874 137116 5182 137125
rect 4874 137114 4880 137116
rect 4936 137114 4960 137116
rect 5016 137114 5040 137116
rect 5096 137114 5120 137116
rect 5176 137114 5182 137116
rect 4936 137062 4938 137114
rect 5118 137062 5120 137114
rect 4874 137060 4880 137062
rect 4936 137060 4960 137062
rect 5016 137060 5040 137062
rect 5096 137060 5120 137062
rect 5176 137060 5182 137062
rect 4874 137051 5182 137060
rect 35594 137116 35902 137125
rect 35594 137114 35600 137116
rect 35656 137114 35680 137116
rect 35736 137114 35760 137116
rect 35816 137114 35840 137116
rect 35896 137114 35902 137116
rect 35656 137062 35658 137114
rect 35838 137062 35840 137114
rect 35594 137060 35600 137062
rect 35656 137060 35680 137062
rect 35736 137060 35760 137062
rect 35816 137060 35840 137062
rect 35896 137060 35902 137062
rect 35594 137051 35902 137060
rect 66314 137116 66622 137125
rect 66314 137114 66320 137116
rect 66376 137114 66400 137116
rect 66456 137114 66480 137116
rect 66536 137114 66560 137116
rect 66616 137114 66622 137116
rect 66376 137062 66378 137114
rect 66558 137062 66560 137114
rect 66314 137060 66320 137062
rect 66376 137060 66400 137062
rect 66456 137060 66480 137062
rect 66536 137060 66560 137062
rect 66616 137060 66622 137062
rect 66314 137051 66622 137060
rect 97034 137116 97342 137125
rect 97034 137114 97040 137116
rect 97096 137114 97120 137116
rect 97176 137114 97200 137116
rect 97256 137114 97280 137116
rect 97336 137114 97342 137116
rect 97096 137062 97098 137114
rect 97278 137062 97280 137114
rect 97034 137060 97040 137062
rect 97096 137060 97120 137062
rect 97176 137060 97200 137062
rect 97256 137060 97280 137062
rect 97336 137060 97342 137062
rect 97034 137051 97342 137060
rect 102140 136876 102192 136882
rect 102140 136818 102192 136824
rect 63592 136672 63644 136678
rect 63592 136614 63644 136620
rect 95976 136672 96028 136678
rect 95976 136614 96028 136620
rect 4214 136572 4522 136581
rect 4214 136570 4220 136572
rect 4276 136570 4300 136572
rect 4356 136570 4380 136572
rect 4436 136570 4460 136572
rect 4516 136570 4522 136572
rect 4276 136518 4278 136570
rect 4458 136518 4460 136570
rect 4214 136516 4220 136518
rect 4276 136516 4300 136518
rect 4356 136516 4380 136518
rect 4436 136516 4460 136518
rect 4516 136516 4522 136518
rect 4214 136507 4522 136516
rect 34934 136572 35242 136581
rect 34934 136570 34940 136572
rect 34996 136570 35020 136572
rect 35076 136570 35100 136572
rect 35156 136570 35180 136572
rect 35236 136570 35242 136572
rect 34996 136518 34998 136570
rect 35178 136518 35180 136570
rect 34934 136516 34940 136518
rect 34996 136516 35020 136518
rect 35076 136516 35100 136518
rect 35156 136516 35180 136518
rect 35236 136516 35242 136518
rect 34934 136507 35242 136516
rect 35992 136264 36044 136270
rect 35992 136206 36044 136212
rect 38568 136264 38620 136270
rect 38568 136206 38620 136212
rect 34152 136196 34204 136202
rect 34152 136138 34204 136144
rect 34980 136196 35032 136202
rect 34980 136138 35032 136144
rect 4874 136028 5182 136037
rect 4874 136026 4880 136028
rect 4936 136026 4960 136028
rect 5016 136026 5040 136028
rect 5096 136026 5120 136028
rect 5176 136026 5182 136028
rect 4936 135974 4938 136026
rect 5118 135974 5120 136026
rect 4874 135972 4880 135974
rect 4936 135972 4960 135974
rect 5016 135972 5040 135974
rect 5096 135972 5120 135974
rect 5176 135972 5182 135974
rect 4874 135963 5182 135972
rect 9588 135924 9640 135930
rect 9588 135866 9640 135872
rect 8208 135856 8260 135862
rect 8208 135798 8260 135804
rect 8024 135788 8076 135794
rect 8024 135730 8076 135736
rect 4214 135484 4522 135493
rect 4214 135482 4220 135484
rect 4276 135482 4300 135484
rect 4356 135482 4380 135484
rect 4436 135482 4460 135484
rect 4516 135482 4522 135484
rect 4276 135430 4278 135482
rect 4458 135430 4460 135482
rect 4214 135428 4220 135430
rect 4276 135428 4300 135430
rect 4356 135428 4380 135430
rect 4436 135428 4460 135430
rect 4516 135428 4522 135430
rect 4214 135419 4522 135428
rect 4874 134940 5182 134949
rect 4874 134938 4880 134940
rect 4936 134938 4960 134940
rect 5016 134938 5040 134940
rect 5096 134938 5120 134940
rect 5176 134938 5182 134940
rect 4936 134886 4938 134938
rect 5118 134886 5120 134938
rect 4874 134884 4880 134886
rect 4936 134884 4960 134886
rect 5016 134884 5040 134886
rect 5096 134884 5120 134886
rect 5176 134884 5182 134886
rect 4874 134875 5182 134884
rect 4214 134396 4522 134405
rect 4214 134394 4220 134396
rect 4276 134394 4300 134396
rect 4356 134394 4380 134396
rect 4436 134394 4460 134396
rect 4516 134394 4522 134396
rect 4276 134342 4278 134394
rect 4458 134342 4460 134394
rect 4214 134340 4220 134342
rect 4276 134340 4300 134342
rect 4356 134340 4380 134342
rect 4436 134340 4460 134342
rect 4516 134340 4522 134342
rect 4214 134331 4522 134340
rect 4874 133852 5182 133861
rect 4874 133850 4880 133852
rect 4936 133850 4960 133852
rect 5016 133850 5040 133852
rect 5096 133850 5120 133852
rect 5176 133850 5182 133852
rect 4936 133798 4938 133850
rect 5118 133798 5120 133850
rect 4874 133796 4880 133798
rect 4936 133796 4960 133798
rect 5016 133796 5040 133798
rect 5096 133796 5120 133798
rect 5176 133796 5182 133798
rect 4874 133787 5182 133796
rect 7380 133748 7432 133754
rect 7380 133690 7432 133696
rect 4214 133308 4522 133317
rect 4214 133306 4220 133308
rect 4276 133306 4300 133308
rect 4356 133306 4380 133308
rect 4436 133306 4460 133308
rect 4516 133306 4522 133308
rect 4276 133254 4278 133306
rect 4458 133254 4460 133306
rect 4214 133252 4220 133254
rect 4276 133252 4300 133254
rect 4356 133252 4380 133254
rect 4436 133252 4460 133254
rect 4516 133252 4522 133254
rect 4214 133243 4522 133252
rect 4874 132764 5182 132773
rect 4874 132762 4880 132764
rect 4936 132762 4960 132764
rect 5016 132762 5040 132764
rect 5096 132762 5120 132764
rect 5176 132762 5182 132764
rect 4936 132710 4938 132762
rect 5118 132710 5120 132762
rect 4874 132708 4880 132710
rect 4936 132708 4960 132710
rect 5016 132708 5040 132710
rect 5096 132708 5120 132710
rect 5176 132708 5182 132710
rect 4874 132699 5182 132708
rect 4214 132220 4522 132229
rect 4214 132218 4220 132220
rect 4276 132218 4300 132220
rect 4356 132218 4380 132220
rect 4436 132218 4460 132220
rect 4516 132218 4522 132220
rect 4276 132166 4278 132218
rect 4458 132166 4460 132218
rect 4214 132164 4220 132166
rect 4276 132164 4300 132166
rect 4356 132164 4380 132166
rect 4436 132164 4460 132166
rect 4516 132164 4522 132166
rect 4214 132155 4522 132164
rect 4874 131676 5182 131685
rect 4874 131674 4880 131676
rect 4936 131674 4960 131676
rect 5016 131674 5040 131676
rect 5096 131674 5120 131676
rect 5176 131674 5182 131676
rect 4936 131622 4938 131674
rect 5118 131622 5120 131674
rect 4874 131620 4880 131622
rect 4936 131620 4960 131622
rect 5016 131620 5040 131622
rect 5096 131620 5120 131622
rect 5176 131620 5182 131622
rect 4874 131611 5182 131620
rect 4214 131132 4522 131141
rect 4214 131130 4220 131132
rect 4276 131130 4300 131132
rect 4356 131130 4380 131132
rect 4436 131130 4460 131132
rect 4516 131130 4522 131132
rect 4276 131078 4278 131130
rect 4458 131078 4460 131130
rect 4214 131076 4220 131078
rect 4276 131076 4300 131078
rect 4356 131076 4380 131078
rect 4436 131076 4460 131078
rect 4516 131076 4522 131078
rect 4214 131067 4522 131076
rect 4874 130588 5182 130597
rect 4874 130586 4880 130588
rect 4936 130586 4960 130588
rect 5016 130586 5040 130588
rect 5096 130586 5120 130588
rect 5176 130586 5182 130588
rect 4936 130534 4938 130586
rect 5118 130534 5120 130586
rect 4874 130532 4880 130534
rect 4936 130532 4960 130534
rect 5016 130532 5040 130534
rect 5096 130532 5120 130534
rect 5176 130532 5182 130534
rect 4874 130523 5182 130532
rect 4214 130044 4522 130053
rect 4214 130042 4220 130044
rect 4276 130042 4300 130044
rect 4356 130042 4380 130044
rect 4436 130042 4460 130044
rect 4516 130042 4522 130044
rect 4276 129990 4278 130042
rect 4458 129990 4460 130042
rect 4214 129988 4220 129990
rect 4276 129988 4300 129990
rect 4356 129988 4380 129990
rect 4436 129988 4460 129990
rect 4516 129988 4522 129990
rect 4214 129979 4522 129988
rect 4874 129500 5182 129509
rect 4874 129498 4880 129500
rect 4936 129498 4960 129500
rect 5016 129498 5040 129500
rect 5096 129498 5120 129500
rect 5176 129498 5182 129500
rect 4936 129446 4938 129498
rect 5118 129446 5120 129498
rect 4874 129444 4880 129446
rect 4936 129444 4960 129446
rect 5016 129444 5040 129446
rect 5096 129444 5120 129446
rect 5176 129444 5182 129446
rect 4874 129435 5182 129444
rect 4214 128956 4522 128965
rect 4214 128954 4220 128956
rect 4276 128954 4300 128956
rect 4356 128954 4380 128956
rect 4436 128954 4460 128956
rect 4516 128954 4522 128956
rect 4276 128902 4278 128954
rect 4458 128902 4460 128954
rect 4214 128900 4220 128902
rect 4276 128900 4300 128902
rect 4356 128900 4380 128902
rect 4436 128900 4460 128902
rect 4516 128900 4522 128902
rect 4214 128891 4522 128900
rect 4874 128412 5182 128421
rect 4874 128410 4880 128412
rect 4936 128410 4960 128412
rect 5016 128410 5040 128412
rect 5096 128410 5120 128412
rect 5176 128410 5182 128412
rect 4936 128358 4938 128410
rect 5118 128358 5120 128410
rect 4874 128356 4880 128358
rect 4936 128356 4960 128358
rect 5016 128356 5040 128358
rect 5096 128356 5120 128358
rect 5176 128356 5182 128358
rect 4874 128347 5182 128356
rect 4214 127868 4522 127877
rect 4214 127866 4220 127868
rect 4276 127866 4300 127868
rect 4356 127866 4380 127868
rect 4436 127866 4460 127868
rect 4516 127866 4522 127868
rect 4276 127814 4278 127866
rect 4458 127814 4460 127866
rect 4214 127812 4220 127814
rect 4276 127812 4300 127814
rect 4356 127812 4380 127814
rect 4436 127812 4460 127814
rect 4516 127812 4522 127814
rect 4214 127803 4522 127812
rect 4874 127324 5182 127333
rect 4874 127322 4880 127324
rect 4936 127322 4960 127324
rect 5016 127322 5040 127324
rect 5096 127322 5120 127324
rect 5176 127322 5182 127324
rect 4936 127270 4938 127322
rect 5118 127270 5120 127322
rect 4874 127268 4880 127270
rect 4936 127268 4960 127270
rect 5016 127268 5040 127270
rect 5096 127268 5120 127270
rect 5176 127268 5182 127270
rect 4874 127259 5182 127268
rect 4214 126780 4522 126789
rect 4214 126778 4220 126780
rect 4276 126778 4300 126780
rect 4356 126778 4380 126780
rect 4436 126778 4460 126780
rect 4516 126778 4522 126780
rect 4276 126726 4278 126778
rect 4458 126726 4460 126778
rect 4214 126724 4220 126726
rect 4276 126724 4300 126726
rect 4356 126724 4380 126726
rect 4436 126724 4460 126726
rect 4516 126724 4522 126726
rect 4214 126715 4522 126724
rect 4874 126236 5182 126245
rect 4874 126234 4880 126236
rect 4936 126234 4960 126236
rect 5016 126234 5040 126236
rect 5096 126234 5120 126236
rect 5176 126234 5182 126236
rect 4936 126182 4938 126234
rect 5118 126182 5120 126234
rect 4874 126180 4880 126182
rect 4936 126180 4960 126182
rect 5016 126180 5040 126182
rect 5096 126180 5120 126182
rect 5176 126180 5182 126182
rect 4874 126171 5182 126180
rect 4214 125692 4522 125701
rect 4214 125690 4220 125692
rect 4276 125690 4300 125692
rect 4356 125690 4380 125692
rect 4436 125690 4460 125692
rect 4516 125690 4522 125692
rect 4276 125638 4278 125690
rect 4458 125638 4460 125690
rect 4214 125636 4220 125638
rect 4276 125636 4300 125638
rect 4356 125636 4380 125638
rect 4436 125636 4460 125638
rect 4516 125636 4522 125638
rect 4214 125627 4522 125636
rect 4874 125148 5182 125157
rect 4874 125146 4880 125148
rect 4936 125146 4960 125148
rect 5016 125146 5040 125148
rect 5096 125146 5120 125148
rect 5176 125146 5182 125148
rect 4936 125094 4938 125146
rect 5118 125094 5120 125146
rect 4874 125092 4880 125094
rect 4936 125092 4960 125094
rect 5016 125092 5040 125094
rect 5096 125092 5120 125094
rect 5176 125092 5182 125094
rect 4874 125083 5182 125092
rect 4214 124604 4522 124613
rect 4214 124602 4220 124604
rect 4276 124602 4300 124604
rect 4356 124602 4380 124604
rect 4436 124602 4460 124604
rect 4516 124602 4522 124604
rect 4276 124550 4278 124602
rect 4458 124550 4460 124602
rect 4214 124548 4220 124550
rect 4276 124548 4300 124550
rect 4356 124548 4380 124550
rect 4436 124548 4460 124550
rect 4516 124548 4522 124550
rect 4214 124539 4522 124548
rect 4874 124060 5182 124069
rect 4874 124058 4880 124060
rect 4936 124058 4960 124060
rect 5016 124058 5040 124060
rect 5096 124058 5120 124060
rect 5176 124058 5182 124060
rect 4936 124006 4938 124058
rect 5118 124006 5120 124058
rect 4874 124004 4880 124006
rect 4936 124004 4960 124006
rect 5016 124004 5040 124006
rect 5096 124004 5120 124006
rect 5176 124004 5182 124006
rect 4874 123995 5182 124004
rect 4214 123516 4522 123525
rect 4214 123514 4220 123516
rect 4276 123514 4300 123516
rect 4356 123514 4380 123516
rect 4436 123514 4460 123516
rect 4516 123514 4522 123516
rect 4276 123462 4278 123514
rect 4458 123462 4460 123514
rect 4214 123460 4220 123462
rect 4276 123460 4300 123462
rect 4356 123460 4380 123462
rect 4436 123460 4460 123462
rect 4516 123460 4522 123462
rect 4214 123451 4522 123460
rect 4874 122972 5182 122981
rect 4874 122970 4880 122972
rect 4936 122970 4960 122972
rect 5016 122970 5040 122972
rect 5096 122970 5120 122972
rect 5176 122970 5182 122972
rect 4936 122918 4938 122970
rect 5118 122918 5120 122970
rect 4874 122916 4880 122918
rect 4936 122916 4960 122918
rect 5016 122916 5040 122918
rect 5096 122916 5120 122918
rect 5176 122916 5182 122918
rect 4874 122907 5182 122916
rect 4214 122428 4522 122437
rect 4214 122426 4220 122428
rect 4276 122426 4300 122428
rect 4356 122426 4380 122428
rect 4436 122426 4460 122428
rect 4516 122426 4522 122428
rect 4276 122374 4278 122426
rect 4458 122374 4460 122426
rect 4214 122372 4220 122374
rect 4276 122372 4300 122374
rect 4356 122372 4380 122374
rect 4436 122372 4460 122374
rect 4516 122372 4522 122374
rect 4214 122363 4522 122372
rect 4874 121884 5182 121893
rect 4874 121882 4880 121884
rect 4936 121882 4960 121884
rect 5016 121882 5040 121884
rect 5096 121882 5120 121884
rect 5176 121882 5182 121884
rect 4936 121830 4938 121882
rect 5118 121830 5120 121882
rect 4874 121828 4880 121830
rect 4936 121828 4960 121830
rect 5016 121828 5040 121830
rect 5096 121828 5120 121830
rect 5176 121828 5182 121830
rect 4874 121819 5182 121828
rect 4214 121340 4522 121349
rect 4214 121338 4220 121340
rect 4276 121338 4300 121340
rect 4356 121338 4380 121340
rect 4436 121338 4460 121340
rect 4516 121338 4522 121340
rect 4276 121286 4278 121338
rect 4458 121286 4460 121338
rect 4214 121284 4220 121286
rect 4276 121284 4300 121286
rect 4356 121284 4380 121286
rect 4436 121284 4460 121286
rect 4516 121284 4522 121286
rect 4214 121275 4522 121284
rect 4874 120796 5182 120805
rect 4874 120794 4880 120796
rect 4936 120794 4960 120796
rect 5016 120794 5040 120796
rect 5096 120794 5120 120796
rect 5176 120794 5182 120796
rect 4936 120742 4938 120794
rect 5118 120742 5120 120794
rect 4874 120740 4880 120742
rect 4936 120740 4960 120742
rect 5016 120740 5040 120742
rect 5096 120740 5120 120742
rect 5176 120740 5182 120742
rect 4874 120731 5182 120740
rect 4214 120252 4522 120261
rect 4214 120250 4220 120252
rect 4276 120250 4300 120252
rect 4356 120250 4380 120252
rect 4436 120250 4460 120252
rect 4516 120250 4522 120252
rect 4276 120198 4278 120250
rect 4458 120198 4460 120250
rect 4214 120196 4220 120198
rect 4276 120196 4300 120198
rect 4356 120196 4380 120198
rect 4436 120196 4460 120198
rect 4516 120196 4522 120198
rect 4214 120187 4522 120196
rect 4874 119708 5182 119717
rect 4874 119706 4880 119708
rect 4936 119706 4960 119708
rect 5016 119706 5040 119708
rect 5096 119706 5120 119708
rect 5176 119706 5182 119708
rect 4936 119654 4938 119706
rect 5118 119654 5120 119706
rect 4874 119652 4880 119654
rect 4936 119652 4960 119654
rect 5016 119652 5040 119654
rect 5096 119652 5120 119654
rect 5176 119652 5182 119654
rect 4874 119643 5182 119652
rect 4214 119164 4522 119173
rect 4214 119162 4220 119164
rect 4276 119162 4300 119164
rect 4356 119162 4380 119164
rect 4436 119162 4460 119164
rect 4516 119162 4522 119164
rect 4276 119110 4278 119162
rect 4458 119110 4460 119162
rect 4214 119108 4220 119110
rect 4276 119108 4300 119110
rect 4356 119108 4380 119110
rect 4436 119108 4460 119110
rect 4516 119108 4522 119110
rect 4214 119099 4522 119108
rect 4874 118620 5182 118629
rect 4874 118618 4880 118620
rect 4936 118618 4960 118620
rect 5016 118618 5040 118620
rect 5096 118618 5120 118620
rect 5176 118618 5182 118620
rect 4936 118566 4938 118618
rect 5118 118566 5120 118618
rect 4874 118564 4880 118566
rect 4936 118564 4960 118566
rect 5016 118564 5040 118566
rect 5096 118564 5120 118566
rect 5176 118564 5182 118566
rect 4874 118555 5182 118564
rect 7392 118522 7420 133690
rect 7380 118516 7432 118522
rect 7380 118458 7432 118464
rect 4214 118076 4522 118085
rect 4214 118074 4220 118076
rect 4276 118074 4300 118076
rect 4356 118074 4380 118076
rect 4436 118074 4460 118076
rect 4516 118074 4522 118076
rect 4276 118022 4278 118074
rect 4458 118022 4460 118074
rect 4214 118020 4220 118022
rect 4276 118020 4300 118022
rect 4356 118020 4380 118022
rect 4436 118020 4460 118022
rect 4516 118020 4522 118022
rect 4214 118011 4522 118020
rect 7392 117706 7420 118458
rect 7472 117768 7524 117774
rect 7472 117710 7524 117716
rect 7380 117700 7432 117706
rect 7380 117642 7432 117648
rect 7288 117632 7340 117638
rect 7288 117574 7340 117580
rect 4874 117532 5182 117541
rect 4874 117530 4880 117532
rect 4936 117530 4960 117532
rect 5016 117530 5040 117532
rect 5096 117530 5120 117532
rect 5176 117530 5182 117532
rect 4936 117478 4938 117530
rect 5118 117478 5120 117530
rect 4874 117476 4880 117478
rect 4936 117476 4960 117478
rect 5016 117476 5040 117478
rect 5096 117476 5120 117478
rect 5176 117476 5182 117478
rect 4874 117467 5182 117476
rect 7300 117094 7328 117574
rect 7484 117094 7512 117710
rect 7288 117088 7340 117094
rect 7288 117030 7340 117036
rect 7472 117088 7524 117094
rect 7472 117030 7524 117036
rect 4214 116988 4522 116997
rect 4214 116986 4220 116988
rect 4276 116986 4300 116988
rect 4356 116986 4380 116988
rect 4436 116986 4460 116988
rect 4516 116986 4522 116988
rect 4276 116934 4278 116986
rect 4458 116934 4460 116986
rect 4214 116932 4220 116934
rect 4276 116932 4300 116934
rect 4356 116932 4380 116934
rect 4436 116932 4460 116934
rect 4516 116932 4522 116934
rect 4214 116923 4522 116932
rect 4874 116444 5182 116453
rect 4874 116442 4880 116444
rect 4936 116442 4960 116444
rect 5016 116442 5040 116444
rect 5096 116442 5120 116444
rect 5176 116442 5182 116444
rect 4936 116390 4938 116442
rect 5118 116390 5120 116442
rect 4874 116388 4880 116390
rect 4936 116388 4960 116390
rect 5016 116388 5040 116390
rect 5096 116388 5120 116390
rect 5176 116388 5182 116390
rect 4874 116379 5182 116388
rect 4214 115900 4522 115909
rect 4214 115898 4220 115900
rect 4276 115898 4300 115900
rect 4356 115898 4380 115900
rect 4436 115898 4460 115900
rect 4516 115898 4522 115900
rect 4276 115846 4278 115898
rect 4458 115846 4460 115898
rect 4214 115844 4220 115846
rect 4276 115844 4300 115846
rect 4356 115844 4380 115846
rect 4436 115844 4460 115846
rect 4516 115844 4522 115846
rect 4214 115835 4522 115844
rect 4874 115356 5182 115365
rect 4874 115354 4880 115356
rect 4936 115354 4960 115356
rect 5016 115354 5040 115356
rect 5096 115354 5120 115356
rect 5176 115354 5182 115356
rect 4936 115302 4938 115354
rect 5118 115302 5120 115354
rect 4874 115300 4880 115302
rect 4936 115300 4960 115302
rect 5016 115300 5040 115302
rect 5096 115300 5120 115302
rect 5176 115300 5182 115302
rect 4874 115291 5182 115300
rect 4214 114812 4522 114821
rect 4214 114810 4220 114812
rect 4276 114810 4300 114812
rect 4356 114810 4380 114812
rect 4436 114810 4460 114812
rect 4516 114810 4522 114812
rect 4276 114758 4278 114810
rect 4458 114758 4460 114810
rect 4214 114756 4220 114758
rect 4276 114756 4300 114758
rect 4356 114756 4380 114758
rect 4436 114756 4460 114758
rect 4516 114756 4522 114758
rect 4214 114747 4522 114756
rect 4874 114268 5182 114277
rect 4874 114266 4880 114268
rect 4936 114266 4960 114268
rect 5016 114266 5040 114268
rect 5096 114266 5120 114268
rect 5176 114266 5182 114268
rect 4936 114214 4938 114266
rect 5118 114214 5120 114266
rect 4874 114212 4880 114214
rect 4936 114212 4960 114214
rect 5016 114212 5040 114214
rect 5096 114212 5120 114214
rect 5176 114212 5182 114214
rect 4874 114203 5182 114212
rect 4214 113724 4522 113733
rect 4214 113722 4220 113724
rect 4276 113722 4300 113724
rect 4356 113722 4380 113724
rect 4436 113722 4460 113724
rect 4516 113722 4522 113724
rect 4276 113670 4278 113722
rect 4458 113670 4460 113722
rect 4214 113668 4220 113670
rect 4276 113668 4300 113670
rect 4356 113668 4380 113670
rect 4436 113668 4460 113670
rect 4516 113668 4522 113670
rect 4214 113659 4522 113668
rect 4874 113180 5182 113189
rect 4874 113178 4880 113180
rect 4936 113178 4960 113180
rect 5016 113178 5040 113180
rect 5096 113178 5120 113180
rect 5176 113178 5182 113180
rect 4936 113126 4938 113178
rect 5118 113126 5120 113178
rect 4874 113124 4880 113126
rect 4936 113124 4960 113126
rect 5016 113124 5040 113126
rect 5096 113124 5120 113126
rect 5176 113124 5182 113126
rect 4874 113115 5182 113124
rect 4214 112636 4522 112645
rect 4214 112634 4220 112636
rect 4276 112634 4300 112636
rect 4356 112634 4380 112636
rect 4436 112634 4460 112636
rect 4516 112634 4522 112636
rect 4276 112582 4278 112634
rect 4458 112582 4460 112634
rect 4214 112580 4220 112582
rect 4276 112580 4300 112582
rect 4356 112580 4380 112582
rect 4436 112580 4460 112582
rect 4516 112580 4522 112582
rect 4214 112571 4522 112580
rect 4874 112092 5182 112101
rect 4874 112090 4880 112092
rect 4936 112090 4960 112092
rect 5016 112090 5040 112092
rect 5096 112090 5120 112092
rect 5176 112090 5182 112092
rect 4936 112038 4938 112090
rect 5118 112038 5120 112090
rect 4874 112036 4880 112038
rect 4936 112036 4960 112038
rect 5016 112036 5040 112038
rect 5096 112036 5120 112038
rect 5176 112036 5182 112038
rect 4874 112027 5182 112036
rect 4214 111548 4522 111557
rect 4214 111546 4220 111548
rect 4276 111546 4300 111548
rect 4356 111546 4380 111548
rect 4436 111546 4460 111548
rect 4516 111546 4522 111548
rect 4276 111494 4278 111546
rect 4458 111494 4460 111546
rect 4214 111492 4220 111494
rect 4276 111492 4300 111494
rect 4356 111492 4380 111494
rect 4436 111492 4460 111494
rect 4516 111492 4522 111494
rect 4214 111483 4522 111492
rect 1308 111240 1360 111246
rect 1308 111182 1360 111188
rect 1320 110945 1348 111182
rect 4874 111004 5182 111013
rect 4874 111002 4880 111004
rect 4936 111002 4960 111004
rect 5016 111002 5040 111004
rect 5096 111002 5120 111004
rect 5176 111002 5182 111004
rect 4936 110950 4938 111002
rect 5118 110950 5120 111002
rect 4874 110948 4880 110950
rect 4936 110948 4960 110950
rect 5016 110948 5040 110950
rect 5096 110948 5120 110950
rect 5176 110948 5182 110950
rect 1306 110936 1362 110945
rect 4874 110939 5182 110948
rect 1306 110871 1362 110880
rect 4214 110460 4522 110469
rect 4214 110458 4220 110460
rect 4276 110458 4300 110460
rect 4356 110458 4380 110460
rect 4436 110458 4460 110460
rect 4516 110458 4522 110460
rect 4276 110406 4278 110458
rect 4458 110406 4460 110458
rect 4214 110404 4220 110406
rect 4276 110404 4300 110406
rect 4356 110404 4380 110406
rect 4436 110404 4460 110406
rect 4516 110404 4522 110406
rect 4214 110395 4522 110404
rect 4874 109916 5182 109925
rect 4874 109914 4880 109916
rect 4936 109914 4960 109916
rect 5016 109914 5040 109916
rect 5096 109914 5120 109916
rect 5176 109914 5182 109916
rect 4936 109862 4938 109914
rect 5118 109862 5120 109914
rect 4874 109860 4880 109862
rect 4936 109860 4960 109862
rect 5016 109860 5040 109862
rect 5096 109860 5120 109862
rect 5176 109860 5182 109862
rect 4874 109851 5182 109860
rect 1308 109676 1360 109682
rect 1308 109618 1360 109624
rect 1320 109585 1348 109618
rect 1306 109576 1362 109585
rect 1306 109511 1362 109520
rect 4214 109372 4522 109381
rect 4214 109370 4220 109372
rect 4276 109370 4300 109372
rect 4356 109370 4380 109372
rect 4436 109370 4460 109372
rect 4516 109370 4522 109372
rect 4276 109318 4278 109370
rect 4458 109318 4460 109370
rect 4214 109316 4220 109318
rect 4276 109316 4300 109318
rect 4356 109316 4380 109318
rect 4436 109316 4460 109318
rect 4516 109316 4522 109318
rect 4214 109307 4522 109316
rect 4874 108828 5182 108837
rect 4874 108826 4880 108828
rect 4936 108826 4960 108828
rect 5016 108826 5040 108828
rect 5096 108826 5120 108828
rect 5176 108826 5182 108828
rect 4936 108774 4938 108826
rect 5118 108774 5120 108826
rect 4874 108772 4880 108774
rect 4936 108772 4960 108774
rect 5016 108772 5040 108774
rect 5096 108772 5120 108774
rect 5176 108772 5182 108774
rect 4874 108763 5182 108772
rect 1308 108588 1360 108594
rect 1308 108530 1360 108536
rect 1320 108225 1348 108530
rect 4214 108284 4522 108293
rect 4214 108282 4220 108284
rect 4276 108282 4300 108284
rect 4356 108282 4380 108284
rect 4436 108282 4460 108284
rect 4516 108282 4522 108284
rect 4276 108230 4278 108282
rect 4458 108230 4460 108282
rect 4214 108228 4220 108230
rect 4276 108228 4300 108230
rect 4356 108228 4380 108230
rect 4436 108228 4460 108230
rect 4516 108228 4522 108230
rect 1306 108216 1362 108225
rect 4214 108219 4522 108228
rect 1306 108151 1362 108160
rect 4874 107740 5182 107749
rect 4874 107738 4880 107740
rect 4936 107738 4960 107740
rect 5016 107738 5040 107740
rect 5096 107738 5120 107740
rect 5176 107738 5182 107740
rect 4936 107686 4938 107738
rect 5118 107686 5120 107738
rect 4874 107684 4880 107686
rect 4936 107684 4960 107686
rect 5016 107684 5040 107686
rect 5096 107684 5120 107686
rect 5176 107684 5182 107686
rect 4874 107675 5182 107684
rect 4214 107196 4522 107205
rect 4214 107194 4220 107196
rect 4276 107194 4300 107196
rect 4356 107194 4380 107196
rect 4436 107194 4460 107196
rect 4516 107194 4522 107196
rect 4276 107142 4278 107194
rect 4458 107142 4460 107194
rect 4214 107140 4220 107142
rect 4276 107140 4300 107142
rect 4356 107140 4380 107142
rect 4436 107140 4460 107142
rect 4516 107140 4522 107142
rect 4214 107131 4522 107140
rect 1216 106888 1268 106894
rect 1214 106856 1216 106865
rect 1268 106856 1270 106865
rect 1214 106791 1270 106800
rect 4874 106652 5182 106661
rect 4874 106650 4880 106652
rect 4936 106650 4960 106652
rect 5016 106650 5040 106652
rect 5096 106650 5120 106652
rect 5176 106650 5182 106652
rect 4936 106598 4938 106650
rect 5118 106598 5120 106650
rect 4874 106596 4880 106598
rect 4936 106596 4960 106598
rect 5016 106596 5040 106598
rect 5096 106596 5120 106598
rect 5176 106596 5182 106598
rect 4874 106587 5182 106596
rect 4214 106108 4522 106117
rect 4214 106106 4220 106108
rect 4276 106106 4300 106108
rect 4356 106106 4380 106108
rect 4436 106106 4460 106108
rect 4516 106106 4522 106108
rect 4276 106054 4278 106106
rect 4458 106054 4460 106106
rect 4214 106052 4220 106054
rect 4276 106052 4300 106054
rect 4356 106052 4380 106054
rect 4436 106052 4460 106054
rect 4516 106052 4522 106054
rect 4214 106043 4522 106052
rect 1308 105800 1360 105806
rect 1308 105742 1360 105748
rect 1320 105505 1348 105742
rect 4874 105564 5182 105573
rect 4874 105562 4880 105564
rect 4936 105562 4960 105564
rect 5016 105562 5040 105564
rect 5096 105562 5120 105564
rect 5176 105562 5182 105564
rect 4936 105510 4938 105562
rect 5118 105510 5120 105562
rect 4874 105508 4880 105510
rect 4936 105508 4960 105510
rect 5016 105508 5040 105510
rect 5096 105508 5120 105510
rect 5176 105508 5182 105510
rect 1306 105496 1362 105505
rect 4874 105499 5182 105508
rect 1306 105431 1362 105440
rect 4214 105020 4522 105029
rect 4214 105018 4220 105020
rect 4276 105018 4300 105020
rect 4356 105018 4380 105020
rect 4436 105018 4460 105020
rect 4516 105018 4522 105020
rect 4276 104966 4278 105018
rect 4458 104966 4460 105018
rect 4214 104964 4220 104966
rect 4276 104964 4300 104966
rect 4356 104964 4380 104966
rect 4436 104964 4460 104966
rect 4516 104964 4522 104966
rect 4214 104955 4522 104964
rect 4874 104476 5182 104485
rect 4874 104474 4880 104476
rect 4936 104474 4960 104476
rect 5016 104474 5040 104476
rect 5096 104474 5120 104476
rect 5176 104474 5182 104476
rect 4936 104422 4938 104474
rect 5118 104422 5120 104474
rect 4874 104420 4880 104422
rect 4936 104420 4960 104422
rect 5016 104420 5040 104422
rect 5096 104420 5120 104422
rect 5176 104420 5182 104422
rect 4874 104411 5182 104420
rect 1308 104236 1360 104242
rect 1308 104178 1360 104184
rect 1320 104145 1348 104178
rect 1306 104136 1362 104145
rect 1306 104071 1362 104080
rect 4214 103932 4522 103941
rect 4214 103930 4220 103932
rect 4276 103930 4300 103932
rect 4356 103930 4380 103932
rect 4436 103930 4460 103932
rect 4516 103930 4522 103932
rect 4276 103878 4278 103930
rect 4458 103878 4460 103930
rect 4214 103876 4220 103878
rect 4276 103876 4300 103878
rect 4356 103876 4380 103878
rect 4436 103876 4460 103878
rect 4516 103876 4522 103878
rect 4214 103867 4522 103876
rect 4874 103388 5182 103397
rect 4874 103386 4880 103388
rect 4936 103386 4960 103388
rect 5016 103386 5040 103388
rect 5096 103386 5120 103388
rect 5176 103386 5182 103388
rect 4936 103334 4938 103386
rect 5118 103334 5120 103386
rect 4874 103332 4880 103334
rect 4936 103332 4960 103334
rect 5016 103332 5040 103334
rect 5096 103332 5120 103334
rect 5176 103332 5182 103334
rect 4874 103323 5182 103332
rect 4214 102844 4522 102853
rect 4214 102842 4220 102844
rect 4276 102842 4300 102844
rect 4356 102842 4380 102844
rect 4436 102842 4460 102844
rect 4516 102842 4522 102844
rect 4276 102790 4278 102842
rect 4458 102790 4460 102842
rect 4214 102788 4220 102790
rect 4276 102788 4300 102790
rect 4356 102788 4380 102790
rect 4436 102788 4460 102790
rect 4516 102788 4522 102790
rect 4214 102779 4522 102788
rect 4874 102300 5182 102309
rect 4874 102298 4880 102300
rect 4936 102298 4960 102300
rect 5016 102298 5040 102300
rect 5096 102298 5120 102300
rect 5176 102298 5182 102300
rect 4936 102246 4938 102298
rect 5118 102246 5120 102298
rect 4874 102244 4880 102246
rect 4936 102244 4960 102246
rect 5016 102244 5040 102246
rect 5096 102244 5120 102246
rect 5176 102244 5182 102246
rect 4874 102235 5182 102244
rect 7300 102202 7328 117030
rect 7288 102196 7340 102202
rect 7288 102138 7340 102144
rect 4214 101756 4522 101765
rect 4214 101754 4220 101756
rect 4276 101754 4300 101756
rect 4356 101754 4380 101756
rect 4436 101754 4460 101756
rect 4516 101754 4522 101756
rect 4276 101702 4278 101754
rect 4458 101702 4460 101754
rect 4214 101700 4220 101702
rect 4276 101700 4300 101702
rect 4356 101700 4380 101702
rect 4436 101700 4460 101702
rect 4516 101700 4522 101702
rect 4214 101691 4522 101700
rect 4874 101212 5182 101221
rect 4874 101210 4880 101212
rect 4936 101210 4960 101212
rect 5016 101210 5040 101212
rect 5096 101210 5120 101212
rect 5176 101210 5182 101212
rect 4936 101158 4938 101210
rect 5118 101158 5120 101210
rect 4874 101156 4880 101158
rect 4936 101156 4960 101158
rect 5016 101156 5040 101158
rect 5096 101156 5120 101158
rect 5176 101156 5182 101158
rect 4874 101147 5182 101156
rect 7380 101108 7432 101114
rect 7380 101050 7432 101056
rect 4214 100668 4522 100677
rect 4214 100666 4220 100668
rect 4276 100666 4300 100668
rect 4356 100666 4380 100668
rect 4436 100666 4460 100668
rect 4516 100666 4522 100668
rect 4276 100614 4278 100666
rect 4458 100614 4460 100666
rect 4214 100612 4220 100614
rect 4276 100612 4300 100614
rect 4356 100612 4380 100614
rect 4436 100612 4460 100614
rect 4516 100612 4522 100614
rect 4214 100603 4522 100612
rect 7392 100298 7420 101050
rect 7484 100366 7512 117030
rect 7472 100360 7524 100366
rect 7472 100302 7524 100308
rect 7380 100292 7432 100298
rect 7380 100234 7432 100240
rect 7288 100224 7340 100230
rect 7288 100166 7340 100172
rect 4874 100124 5182 100133
rect 4874 100122 4880 100124
rect 4936 100122 4960 100124
rect 5016 100122 5040 100124
rect 5096 100122 5120 100124
rect 5176 100122 5182 100124
rect 4936 100070 4938 100122
rect 5118 100070 5120 100122
rect 4874 100068 4880 100070
rect 4936 100068 4960 100070
rect 5016 100068 5040 100070
rect 5096 100068 5120 100070
rect 5176 100068 5182 100070
rect 4874 100059 5182 100068
rect 7300 99686 7328 100166
rect 7484 100026 7512 100302
rect 7472 100020 7524 100026
rect 7472 99962 7524 99968
rect 7288 99680 7340 99686
rect 7288 99622 7340 99628
rect 4214 99580 4522 99589
rect 4214 99578 4220 99580
rect 4276 99578 4300 99580
rect 4356 99578 4380 99580
rect 4436 99578 4460 99580
rect 4516 99578 4522 99580
rect 4276 99526 4278 99578
rect 4458 99526 4460 99578
rect 4214 99524 4220 99526
rect 4276 99524 4300 99526
rect 4356 99524 4380 99526
rect 4436 99524 4460 99526
rect 4516 99524 4522 99526
rect 4214 99515 4522 99524
rect 4874 99036 5182 99045
rect 4874 99034 4880 99036
rect 4936 99034 4960 99036
rect 5016 99034 5040 99036
rect 5096 99034 5120 99036
rect 5176 99034 5182 99036
rect 4936 98982 4938 99034
rect 5118 98982 5120 99034
rect 4874 98980 4880 98982
rect 4936 98980 4960 98982
rect 5016 98980 5040 98982
rect 5096 98980 5120 98982
rect 5176 98980 5182 98982
rect 4874 98971 5182 98980
rect 4214 98492 4522 98501
rect 4214 98490 4220 98492
rect 4276 98490 4300 98492
rect 4356 98490 4380 98492
rect 4436 98490 4460 98492
rect 4516 98490 4522 98492
rect 4276 98438 4278 98490
rect 4458 98438 4460 98490
rect 4214 98436 4220 98438
rect 4276 98436 4300 98438
rect 4356 98436 4380 98438
rect 4436 98436 4460 98438
rect 4516 98436 4522 98438
rect 4214 98427 4522 98436
rect 4874 97948 5182 97957
rect 4874 97946 4880 97948
rect 4936 97946 4960 97948
rect 5016 97946 5040 97948
rect 5096 97946 5120 97948
rect 5176 97946 5182 97948
rect 4936 97894 4938 97946
rect 5118 97894 5120 97946
rect 4874 97892 4880 97894
rect 4936 97892 4960 97894
rect 5016 97892 5040 97894
rect 5096 97892 5120 97894
rect 5176 97892 5182 97894
rect 4874 97883 5182 97892
rect 4214 97404 4522 97413
rect 4214 97402 4220 97404
rect 4276 97402 4300 97404
rect 4356 97402 4380 97404
rect 4436 97402 4460 97404
rect 4516 97402 4522 97404
rect 4276 97350 4278 97402
rect 4458 97350 4460 97402
rect 4214 97348 4220 97350
rect 4276 97348 4300 97350
rect 4356 97348 4380 97350
rect 4436 97348 4460 97350
rect 4516 97348 4522 97350
rect 4214 97339 4522 97348
rect 4874 96860 5182 96869
rect 4874 96858 4880 96860
rect 4936 96858 4960 96860
rect 5016 96858 5040 96860
rect 5096 96858 5120 96860
rect 5176 96858 5182 96860
rect 4936 96806 4938 96858
rect 5118 96806 5120 96858
rect 4874 96804 4880 96806
rect 4936 96804 4960 96806
rect 5016 96804 5040 96806
rect 5096 96804 5120 96806
rect 5176 96804 5182 96806
rect 4874 96795 5182 96804
rect 4214 96316 4522 96325
rect 4214 96314 4220 96316
rect 4276 96314 4300 96316
rect 4356 96314 4380 96316
rect 4436 96314 4460 96316
rect 4516 96314 4522 96316
rect 4276 96262 4278 96314
rect 4458 96262 4460 96314
rect 4214 96260 4220 96262
rect 4276 96260 4300 96262
rect 4356 96260 4380 96262
rect 4436 96260 4460 96262
rect 4516 96260 4522 96262
rect 4214 96251 4522 96260
rect 4874 95772 5182 95781
rect 4874 95770 4880 95772
rect 4936 95770 4960 95772
rect 5016 95770 5040 95772
rect 5096 95770 5120 95772
rect 5176 95770 5182 95772
rect 4936 95718 4938 95770
rect 5118 95718 5120 95770
rect 4874 95716 4880 95718
rect 4936 95716 4960 95718
rect 5016 95716 5040 95718
rect 5096 95716 5120 95718
rect 5176 95716 5182 95718
rect 4874 95707 5182 95716
rect 4214 95228 4522 95237
rect 4214 95226 4220 95228
rect 4276 95226 4300 95228
rect 4356 95226 4380 95228
rect 4436 95226 4460 95228
rect 4516 95226 4522 95228
rect 4276 95174 4278 95226
rect 4458 95174 4460 95226
rect 4214 95172 4220 95174
rect 4276 95172 4300 95174
rect 4356 95172 4380 95174
rect 4436 95172 4460 95174
rect 4516 95172 4522 95174
rect 4214 95163 4522 95172
rect 5816 94852 5868 94858
rect 5816 94794 5868 94800
rect 4874 94684 5182 94693
rect 4874 94682 4880 94684
rect 4936 94682 4960 94684
rect 5016 94682 5040 94684
rect 5096 94682 5120 94684
rect 5176 94682 5182 94684
rect 4936 94630 4938 94682
rect 5118 94630 5120 94682
rect 4874 94628 4880 94630
rect 4936 94628 4960 94630
rect 5016 94628 5040 94630
rect 5096 94628 5120 94630
rect 5176 94628 5182 94630
rect 4874 94619 5182 94628
rect 4214 94140 4522 94149
rect 4214 94138 4220 94140
rect 4276 94138 4300 94140
rect 4356 94138 4380 94140
rect 4436 94138 4460 94140
rect 4516 94138 4522 94140
rect 4276 94086 4278 94138
rect 4458 94086 4460 94138
rect 4214 94084 4220 94086
rect 4276 94084 4300 94086
rect 4356 94084 4380 94086
rect 4436 94084 4460 94086
rect 4516 94084 4522 94086
rect 4214 94075 4522 94084
rect 4874 93596 5182 93605
rect 4874 93594 4880 93596
rect 4936 93594 4960 93596
rect 5016 93594 5040 93596
rect 5096 93594 5120 93596
rect 5176 93594 5182 93596
rect 4936 93542 4938 93594
rect 5118 93542 5120 93594
rect 4874 93540 4880 93542
rect 4936 93540 4960 93542
rect 5016 93540 5040 93542
rect 5096 93540 5120 93542
rect 5176 93540 5182 93542
rect 4874 93531 5182 93540
rect 4214 93052 4522 93061
rect 4214 93050 4220 93052
rect 4276 93050 4300 93052
rect 4356 93050 4380 93052
rect 4436 93050 4460 93052
rect 4516 93050 4522 93052
rect 4276 92998 4278 93050
rect 4458 92998 4460 93050
rect 4214 92996 4220 92998
rect 4276 92996 4300 92998
rect 4356 92996 4380 92998
rect 4436 92996 4460 92998
rect 4516 92996 4522 92998
rect 4214 92987 4522 92996
rect 4874 92508 5182 92517
rect 4874 92506 4880 92508
rect 4936 92506 4960 92508
rect 5016 92506 5040 92508
rect 5096 92506 5120 92508
rect 5176 92506 5182 92508
rect 4936 92454 4938 92506
rect 5118 92454 5120 92506
rect 4874 92452 4880 92454
rect 4936 92452 4960 92454
rect 5016 92452 5040 92454
rect 5096 92452 5120 92454
rect 5176 92452 5182 92454
rect 4874 92443 5182 92452
rect 4214 91964 4522 91973
rect 4214 91962 4220 91964
rect 4276 91962 4300 91964
rect 4356 91962 4380 91964
rect 4436 91962 4460 91964
rect 4516 91962 4522 91964
rect 4276 91910 4278 91962
rect 4458 91910 4460 91962
rect 4214 91908 4220 91910
rect 4276 91908 4300 91910
rect 4356 91908 4380 91910
rect 4436 91908 4460 91910
rect 4516 91908 4522 91910
rect 4214 91899 4522 91908
rect 4874 91420 5182 91429
rect 4874 91418 4880 91420
rect 4936 91418 4960 91420
rect 5016 91418 5040 91420
rect 5096 91418 5120 91420
rect 5176 91418 5182 91420
rect 4936 91366 4938 91418
rect 5118 91366 5120 91418
rect 4874 91364 4880 91366
rect 4936 91364 4960 91366
rect 5016 91364 5040 91366
rect 5096 91364 5120 91366
rect 5176 91364 5182 91366
rect 4874 91355 5182 91364
rect 4214 90876 4522 90885
rect 4214 90874 4220 90876
rect 4276 90874 4300 90876
rect 4356 90874 4380 90876
rect 4436 90874 4460 90876
rect 4516 90874 4522 90876
rect 4276 90822 4278 90874
rect 4458 90822 4460 90874
rect 4214 90820 4220 90822
rect 4276 90820 4300 90822
rect 4356 90820 4380 90822
rect 4436 90820 4460 90822
rect 4516 90820 4522 90822
rect 4214 90811 4522 90820
rect 4874 90332 5182 90341
rect 4874 90330 4880 90332
rect 4936 90330 4960 90332
rect 5016 90330 5040 90332
rect 5096 90330 5120 90332
rect 5176 90330 5182 90332
rect 4936 90278 4938 90330
rect 5118 90278 5120 90330
rect 4874 90276 4880 90278
rect 4936 90276 4960 90278
rect 5016 90276 5040 90278
rect 5096 90276 5120 90278
rect 5176 90276 5182 90278
rect 4874 90267 5182 90276
rect 4214 89788 4522 89797
rect 4214 89786 4220 89788
rect 4276 89786 4300 89788
rect 4356 89786 4380 89788
rect 4436 89786 4460 89788
rect 4516 89786 4522 89788
rect 4276 89734 4278 89786
rect 4458 89734 4460 89786
rect 4214 89732 4220 89734
rect 4276 89732 4300 89734
rect 4356 89732 4380 89734
rect 4436 89732 4460 89734
rect 4516 89732 4522 89734
rect 4214 89723 4522 89732
rect 4874 89244 5182 89253
rect 4874 89242 4880 89244
rect 4936 89242 4960 89244
rect 5016 89242 5040 89244
rect 5096 89242 5120 89244
rect 5176 89242 5182 89244
rect 4936 89190 4938 89242
rect 5118 89190 5120 89242
rect 4874 89188 4880 89190
rect 4936 89188 4960 89190
rect 5016 89188 5040 89190
rect 5096 89188 5120 89190
rect 5176 89188 5182 89190
rect 4874 89179 5182 89188
rect 1308 89004 1360 89010
rect 1308 88946 1360 88952
rect 1320 88505 1348 88946
rect 4214 88700 4522 88709
rect 4214 88698 4220 88700
rect 4276 88698 4300 88700
rect 4356 88698 4380 88700
rect 4436 88698 4460 88700
rect 4516 88698 4522 88700
rect 4276 88646 4278 88698
rect 4458 88646 4460 88698
rect 4214 88644 4220 88646
rect 4276 88644 4300 88646
rect 4356 88644 4380 88646
rect 4436 88644 4460 88646
rect 4516 88644 4522 88646
rect 4214 88635 4522 88644
rect 1306 88496 1362 88505
rect 1306 88431 1362 88440
rect 4874 88156 5182 88165
rect 4874 88154 4880 88156
rect 4936 88154 4960 88156
rect 5016 88154 5040 88156
rect 5096 88154 5120 88156
rect 5176 88154 5182 88156
rect 4936 88102 4938 88154
rect 5118 88102 5120 88154
rect 4874 88100 4880 88102
rect 4936 88100 4960 88102
rect 5016 88100 5040 88102
rect 5096 88100 5120 88102
rect 5176 88100 5182 88102
rect 4874 88091 5182 88100
rect 1216 87916 1268 87922
rect 1216 87858 1268 87864
rect 1228 87825 1256 87858
rect 1214 87816 1270 87825
rect 1214 87751 1270 87760
rect 4214 87612 4522 87621
rect 4214 87610 4220 87612
rect 4276 87610 4300 87612
rect 4356 87610 4380 87612
rect 4436 87610 4460 87612
rect 4516 87610 4522 87612
rect 4276 87558 4278 87610
rect 4458 87558 4460 87610
rect 4214 87556 4220 87558
rect 4276 87556 4300 87558
rect 4356 87556 4380 87558
rect 4436 87556 4460 87558
rect 4516 87556 4522 87558
rect 4214 87547 4522 87556
rect 1216 87236 1268 87242
rect 1216 87178 1268 87184
rect 1228 87145 1256 87178
rect 1860 87168 1912 87174
rect 1214 87136 1270 87145
rect 1860 87110 1912 87116
rect 1214 87071 1270 87080
rect 1308 86828 1360 86834
rect 1308 86770 1360 86776
rect 1320 86465 1348 86770
rect 1306 86456 1362 86465
rect 1306 86391 1362 86400
rect 1308 86216 1360 86222
rect 1308 86158 1360 86164
rect 1320 85785 1348 86158
rect 1306 85776 1362 85785
rect 1306 85711 1362 85720
rect 1872 85610 1900 87110
rect 4874 87068 5182 87077
rect 4874 87066 4880 87068
rect 4936 87066 4960 87068
rect 5016 87066 5040 87068
rect 5096 87066 5120 87068
rect 5176 87066 5182 87068
rect 4936 87014 4938 87066
rect 5118 87014 5120 87066
rect 4874 87012 4880 87014
rect 4936 87012 4960 87014
rect 5016 87012 5040 87014
rect 5096 87012 5120 87014
rect 5176 87012 5182 87014
rect 4874 87003 5182 87012
rect 4214 86524 4522 86533
rect 4214 86522 4220 86524
rect 4276 86522 4300 86524
rect 4356 86522 4380 86524
rect 4436 86522 4460 86524
rect 4516 86522 4522 86524
rect 4276 86470 4278 86522
rect 4458 86470 4460 86522
rect 4214 86468 4220 86470
rect 4276 86468 4300 86470
rect 4356 86468 4380 86470
rect 4436 86468 4460 86470
rect 4516 86468 4522 86470
rect 4214 86459 4522 86468
rect 5540 86080 5592 86086
rect 5540 86022 5592 86028
rect 4874 85980 5182 85989
rect 4874 85978 4880 85980
rect 4936 85978 4960 85980
rect 5016 85978 5040 85980
rect 5096 85978 5120 85980
rect 5176 85978 5182 85980
rect 4936 85926 4938 85978
rect 5118 85926 5120 85978
rect 4874 85924 4880 85926
rect 4936 85924 4960 85926
rect 5016 85924 5040 85926
rect 5096 85924 5120 85926
rect 5176 85924 5182 85926
rect 4874 85915 5182 85924
rect 1860 85604 1912 85610
rect 1860 85546 1912 85552
rect 5552 85513 5580 86022
rect 5538 85504 5594 85513
rect 4214 85436 4522 85445
rect 5538 85439 5594 85448
rect 4214 85434 4220 85436
rect 4276 85434 4300 85436
rect 4356 85434 4380 85436
rect 4436 85434 4460 85436
rect 4516 85434 4522 85436
rect 4276 85382 4278 85434
rect 4458 85382 4460 85434
rect 4214 85380 4220 85382
rect 4276 85380 4300 85382
rect 4356 85380 4380 85382
rect 4436 85380 4460 85382
rect 4516 85380 4522 85382
rect 4214 85371 4522 85380
rect 1214 85096 1270 85105
rect 1214 85031 1216 85040
rect 1268 85031 1270 85040
rect 1216 85002 1268 85008
rect 2044 84992 2096 84998
rect 2044 84934 2096 84940
rect 1308 84652 1360 84658
rect 1308 84594 1360 84600
rect 1320 84425 1348 84594
rect 1860 84516 1912 84522
rect 1860 84458 1912 84464
rect 1306 84416 1362 84425
rect 1306 84351 1362 84360
rect 1872 84182 1900 84458
rect 1860 84176 1912 84182
rect 1860 84118 1912 84124
rect 1308 84040 1360 84046
rect 1308 83982 1360 83988
rect 1320 83745 1348 83982
rect 1306 83736 1362 83745
rect 1306 83671 1362 83680
rect 1308 83564 1360 83570
rect 1308 83506 1360 83512
rect 1320 83065 1348 83506
rect 2056 83502 2084 84934
rect 4874 84892 5182 84901
rect 4874 84890 4880 84892
rect 4936 84890 4960 84892
rect 5016 84890 5040 84892
rect 5096 84890 5120 84892
rect 5176 84890 5182 84892
rect 4936 84838 4938 84890
rect 5118 84838 5120 84890
rect 4874 84836 4880 84838
rect 4936 84836 4960 84838
rect 5016 84836 5040 84838
rect 5096 84836 5120 84838
rect 5176 84836 5182 84838
rect 4874 84827 5182 84836
rect 4214 84348 4522 84357
rect 4214 84346 4220 84348
rect 4276 84346 4300 84348
rect 4356 84346 4380 84348
rect 4436 84346 4460 84348
rect 4516 84346 4522 84348
rect 4276 84294 4278 84346
rect 4458 84294 4460 84346
rect 4214 84292 4220 84294
rect 4276 84292 4300 84294
rect 4356 84292 4380 84294
rect 4436 84292 4460 84294
rect 4516 84292 4522 84294
rect 4214 84283 4522 84292
rect 2504 83904 2556 83910
rect 2504 83846 2556 83852
rect 2044 83496 2096 83502
rect 2044 83438 2096 83444
rect 2044 83360 2096 83366
rect 2044 83302 2096 83308
rect 1306 83056 1362 83065
rect 1306 82991 1362 83000
rect 1216 82476 1268 82482
rect 1216 82418 1268 82424
rect 1228 82385 1256 82418
rect 1214 82376 1270 82385
rect 1214 82311 1270 82320
rect 1216 81796 1268 81802
rect 1216 81738 1268 81744
rect 1228 81705 1256 81738
rect 1860 81728 1912 81734
rect 1214 81696 1270 81705
rect 1860 81670 1912 81676
rect 1214 81631 1270 81640
rect 1308 81388 1360 81394
rect 1308 81330 1360 81336
rect 1320 81025 1348 81330
rect 1306 81016 1362 81025
rect 1306 80951 1362 80960
rect 1872 80850 1900 81670
rect 2056 81326 2084 83302
rect 2044 81320 2096 81326
rect 2044 81262 2096 81268
rect 1860 80844 1912 80850
rect 1860 80786 1912 80792
rect 1308 80776 1360 80782
rect 1308 80718 1360 80724
rect 1320 80374 1348 80718
rect 2516 80714 2544 83846
rect 4874 83804 5182 83813
rect 4874 83802 4880 83804
rect 4936 83802 4960 83804
rect 5016 83802 5040 83804
rect 5096 83802 5120 83804
rect 5176 83802 5182 83804
rect 4936 83750 4938 83802
rect 5118 83750 5120 83802
rect 4874 83748 4880 83750
rect 4936 83748 4960 83750
rect 5016 83748 5040 83750
rect 5096 83748 5120 83750
rect 5176 83748 5182 83750
rect 4874 83739 5182 83748
rect 4214 83260 4522 83269
rect 4214 83258 4220 83260
rect 4276 83258 4300 83260
rect 4356 83258 4380 83260
rect 4436 83258 4460 83260
rect 4516 83258 4522 83260
rect 4276 83206 4278 83258
rect 4458 83206 4460 83258
rect 4214 83204 4220 83206
rect 4276 83204 4300 83206
rect 4356 83204 4380 83206
rect 4436 83204 4460 83206
rect 4516 83204 4522 83206
rect 4214 83195 4522 83204
rect 4874 82716 5182 82725
rect 4874 82714 4880 82716
rect 4936 82714 4960 82716
rect 5016 82714 5040 82716
rect 5096 82714 5120 82716
rect 5176 82714 5182 82716
rect 4936 82662 4938 82714
rect 5118 82662 5120 82714
rect 4874 82660 4880 82662
rect 4936 82660 4960 82662
rect 5016 82660 5040 82662
rect 5096 82660 5120 82662
rect 5176 82660 5182 82662
rect 4874 82651 5182 82660
rect 5264 82408 5316 82414
rect 5264 82350 5316 82356
rect 2688 82272 2740 82278
rect 2688 82214 2740 82220
rect 2700 80782 2728 82214
rect 4214 82172 4522 82181
rect 4214 82170 4220 82172
rect 4276 82170 4300 82172
rect 4356 82170 4380 82172
rect 4436 82170 4460 82172
rect 4516 82170 4522 82172
rect 4276 82118 4278 82170
rect 4458 82118 4460 82170
rect 4214 82116 4220 82118
rect 4276 82116 4300 82118
rect 4356 82116 4380 82118
rect 4436 82116 4460 82118
rect 4516 82116 4522 82118
rect 4214 82107 4522 82116
rect 4874 81628 5182 81637
rect 4874 81626 4880 81628
rect 4936 81626 4960 81628
rect 5016 81626 5040 81628
rect 5096 81626 5120 81628
rect 5176 81626 5182 81628
rect 4936 81574 4938 81626
rect 5118 81574 5120 81626
rect 4874 81572 4880 81574
rect 4936 81572 4960 81574
rect 5016 81572 5040 81574
rect 5096 81572 5120 81574
rect 5176 81572 5182 81574
rect 4874 81563 5182 81572
rect 4214 81084 4522 81093
rect 4214 81082 4220 81084
rect 4276 81082 4300 81084
rect 4356 81082 4380 81084
rect 4436 81082 4460 81084
rect 4516 81082 4522 81084
rect 4276 81030 4278 81082
rect 4458 81030 4460 81082
rect 4214 81028 4220 81030
rect 4276 81028 4300 81030
rect 4356 81028 4380 81030
rect 4436 81028 4460 81030
rect 4516 81028 4522 81030
rect 4214 81019 4522 81028
rect 2688 80776 2740 80782
rect 2688 80718 2740 80724
rect 2504 80708 2556 80714
rect 2504 80650 2556 80656
rect 4874 80540 5182 80549
rect 4874 80538 4880 80540
rect 4936 80538 4960 80540
rect 5016 80538 5040 80540
rect 5096 80538 5120 80540
rect 5176 80538 5182 80540
rect 4936 80486 4938 80538
rect 5118 80486 5120 80538
rect 4874 80484 4880 80486
rect 4936 80484 4960 80486
rect 5016 80484 5040 80486
rect 5096 80484 5120 80486
rect 5176 80484 5182 80486
rect 4874 80475 5182 80484
rect 1308 80368 1360 80374
rect 1306 80336 1308 80345
rect 1360 80336 1362 80345
rect 1306 80271 1362 80280
rect 4214 79996 4522 80005
rect 4214 79994 4220 79996
rect 4276 79994 4300 79996
rect 4356 79994 4380 79996
rect 4436 79994 4460 79996
rect 4516 79994 4522 79996
rect 4276 79942 4278 79994
rect 4458 79942 4460 79994
rect 4214 79940 4220 79942
rect 4276 79940 4300 79942
rect 4356 79940 4380 79942
rect 4436 79940 4460 79942
rect 4516 79940 4522 79942
rect 4214 79931 4522 79940
rect 1214 79656 1270 79665
rect 1214 79591 1216 79600
rect 1268 79591 1270 79600
rect 1216 79562 1268 79568
rect 4874 79452 5182 79461
rect 4874 79450 4880 79452
rect 4936 79450 4960 79452
rect 5016 79450 5040 79452
rect 5096 79450 5120 79452
rect 5176 79450 5182 79452
rect 4936 79398 4938 79450
rect 5118 79398 5120 79450
rect 4874 79396 4880 79398
rect 4936 79396 4960 79398
rect 5016 79396 5040 79398
rect 5096 79396 5120 79398
rect 5176 79396 5182 79398
rect 4874 79387 5182 79396
rect 1308 79212 1360 79218
rect 1308 79154 1360 79160
rect 1320 78985 1348 79154
rect 1306 78976 1362 78985
rect 1306 78911 1362 78920
rect 4214 78908 4522 78917
rect 4214 78906 4220 78908
rect 4276 78906 4300 78908
rect 4356 78906 4380 78908
rect 4436 78906 4460 78908
rect 4516 78906 4522 78908
rect 4276 78854 4278 78906
rect 4458 78854 4460 78906
rect 4214 78852 4220 78854
rect 4276 78852 4300 78854
rect 4356 78852 4380 78854
rect 4436 78852 4460 78854
rect 4516 78852 4522 78854
rect 4214 78843 4522 78852
rect 1308 78532 1360 78538
rect 1308 78474 1360 78480
rect 1320 78305 1348 78474
rect 4874 78364 5182 78373
rect 4874 78362 4880 78364
rect 4936 78362 4960 78364
rect 5016 78362 5040 78364
rect 5096 78362 5120 78364
rect 5176 78362 5182 78364
rect 4936 78310 4938 78362
rect 5118 78310 5120 78362
rect 4874 78308 4880 78310
rect 4936 78308 4960 78310
rect 5016 78308 5040 78310
rect 5096 78308 5120 78310
rect 5176 78308 5182 78310
rect 1306 78296 1362 78305
rect 4874 78299 5182 78308
rect 1306 78231 1362 78240
rect 1308 78124 1360 78130
rect 1308 78066 1360 78072
rect 2044 78124 2096 78130
rect 2044 78066 2096 78072
rect 1320 77625 1348 78066
rect 1306 77616 1362 77625
rect 1306 77551 1362 77560
rect 2056 77178 2084 78066
rect 4214 77820 4522 77829
rect 4214 77818 4220 77820
rect 4276 77818 4300 77820
rect 4356 77818 4380 77820
rect 4436 77818 4460 77820
rect 4516 77818 4522 77820
rect 4276 77766 4278 77818
rect 4458 77766 4460 77818
rect 4214 77764 4220 77766
rect 4276 77764 4300 77766
rect 4356 77764 4380 77766
rect 4436 77764 4460 77766
rect 4516 77764 4522 77766
rect 4214 77755 4522 77764
rect 4874 77276 5182 77285
rect 4874 77274 4880 77276
rect 4936 77274 4960 77276
rect 5016 77274 5040 77276
rect 5096 77274 5120 77276
rect 5176 77274 5182 77276
rect 4936 77222 4938 77274
rect 5118 77222 5120 77274
rect 4874 77220 4880 77222
rect 4936 77220 4960 77222
rect 5016 77220 5040 77222
rect 5096 77220 5120 77222
rect 5176 77220 5182 77222
rect 4874 77211 5182 77220
rect 2044 77172 2096 77178
rect 2044 77114 2096 77120
rect 1216 77036 1268 77042
rect 1216 76978 1268 76984
rect 1228 76945 1256 76978
rect 1214 76936 1270 76945
rect 1214 76871 1270 76880
rect 4214 76732 4522 76741
rect 4214 76730 4220 76732
rect 4276 76730 4300 76732
rect 4356 76730 4380 76732
rect 4436 76730 4460 76732
rect 4516 76730 4522 76732
rect 4276 76678 4278 76730
rect 4458 76678 4460 76730
rect 4214 76676 4220 76678
rect 4276 76676 4300 76678
rect 4356 76676 4380 76678
rect 4436 76676 4460 76678
rect 4516 76676 4522 76678
rect 4214 76667 4522 76676
rect 846 76392 902 76401
rect 846 76327 902 76336
rect 860 76294 888 76327
rect 848 76288 900 76294
rect 848 76230 900 76236
rect 4874 76188 5182 76197
rect 4874 76186 4880 76188
rect 4936 76186 4960 76188
rect 5016 76186 5040 76188
rect 5096 76186 5120 76188
rect 5176 76186 5182 76188
rect 4936 76134 4938 76186
rect 5118 76134 5120 76186
rect 4874 76132 4880 76134
rect 4936 76132 4960 76134
rect 5016 76132 5040 76134
rect 5096 76132 5120 76134
rect 5176 76132 5182 76134
rect 4874 76123 5182 76132
rect 1492 75744 1544 75750
rect 1492 75686 1544 75692
rect 1504 75585 1532 75686
rect 4214 75644 4522 75653
rect 4214 75642 4220 75644
rect 4276 75642 4300 75644
rect 4356 75642 4380 75644
rect 4436 75642 4460 75644
rect 4516 75642 4522 75644
rect 4276 75590 4278 75642
rect 4458 75590 4460 75642
rect 4214 75588 4220 75590
rect 4276 75588 4300 75590
rect 4356 75588 4380 75590
rect 4436 75588 4460 75590
rect 4516 75588 4522 75590
rect 1490 75576 1546 75585
rect 4214 75579 4522 75588
rect 1490 75511 1546 75520
rect 848 75200 900 75206
rect 848 75142 900 75148
rect 860 75041 888 75142
rect 4874 75100 5182 75109
rect 4874 75098 4880 75100
rect 4936 75098 4960 75100
rect 5016 75098 5040 75100
rect 5096 75098 5120 75100
rect 5176 75098 5182 75100
rect 4936 75046 4938 75098
rect 5118 75046 5120 75098
rect 4874 75044 4880 75046
rect 4936 75044 4960 75046
rect 5016 75044 5040 75046
rect 5096 75044 5120 75046
rect 5176 75044 5182 75046
rect 846 75032 902 75041
rect 4874 75035 5182 75044
rect 846 74967 902 74976
rect 4214 74556 4522 74565
rect 4214 74554 4220 74556
rect 4276 74554 4300 74556
rect 4356 74554 4380 74556
rect 4436 74554 4460 74556
rect 4516 74554 4522 74556
rect 4276 74502 4278 74554
rect 4458 74502 4460 74554
rect 4214 74500 4220 74502
rect 4276 74500 4300 74502
rect 4356 74500 4380 74502
rect 4436 74500 4460 74502
rect 4516 74500 4522 74502
rect 4214 74491 4522 74500
rect 848 74384 900 74390
rect 846 74352 848 74361
rect 900 74352 902 74361
rect 846 74287 902 74296
rect 4874 74012 5182 74021
rect 4874 74010 4880 74012
rect 4936 74010 4960 74012
rect 5016 74010 5040 74012
rect 5096 74010 5120 74012
rect 5176 74010 5182 74012
rect 4936 73958 4938 74010
rect 5118 73958 5120 74010
rect 4874 73956 4880 73958
rect 4936 73956 4960 73958
rect 5016 73956 5040 73958
rect 5096 73956 5120 73958
rect 5176 73956 5182 73958
rect 4874 73947 5182 73956
rect 846 73672 902 73681
rect 846 73607 848 73616
rect 900 73607 902 73616
rect 848 73578 900 73584
rect 1860 73568 1912 73574
rect 1860 73510 1912 73516
rect 1872 73370 1900 73510
rect 4214 73468 4522 73477
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73403 4522 73412
rect 1860 73364 1912 73370
rect 1860 73306 1912 73312
rect 848 73024 900 73030
rect 846 72992 848 73001
rect 900 72992 902 73001
rect 846 72927 902 72936
rect 4874 72924 5182 72933
rect 4874 72922 4880 72924
rect 4936 72922 4960 72924
rect 5016 72922 5040 72924
rect 5096 72922 5120 72924
rect 5176 72922 5182 72924
rect 4936 72870 4938 72922
rect 5118 72870 5120 72922
rect 4874 72868 4880 72870
rect 4936 72868 4960 72870
rect 5016 72868 5040 72870
rect 5096 72868 5120 72870
rect 5176 72868 5182 72870
rect 4874 72859 5182 72868
rect 848 72480 900 72486
rect 848 72422 900 72428
rect 860 72321 888 72422
rect 4214 72380 4522 72389
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 846 72312 902 72321
rect 4214 72315 4522 72324
rect 846 72247 902 72256
rect 4874 71836 5182 71845
rect 4874 71834 4880 71836
rect 4936 71834 4960 71836
rect 5016 71834 5040 71836
rect 5096 71834 5120 71836
rect 5176 71834 5182 71836
rect 4936 71782 4938 71834
rect 5118 71782 5120 71834
rect 4874 71780 4880 71782
rect 4936 71780 4960 71782
rect 5016 71780 5040 71782
rect 5096 71780 5120 71782
rect 5176 71780 5182 71782
rect 4874 71771 5182 71780
rect 1216 71596 1268 71602
rect 1216 71538 1268 71544
rect 1228 71505 1256 71538
rect 1214 71496 1270 71505
rect 1214 71431 1270 71440
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 5276 70922 5304 82350
rect 5828 82278 5856 94794
rect 7104 93696 7156 93702
rect 7104 93638 7156 93644
rect 7116 93158 7144 93638
rect 7104 93152 7156 93158
rect 7104 93094 7156 93100
rect 5816 82272 5868 82278
rect 5816 82214 5868 82220
rect 6184 82272 6236 82278
rect 6184 82214 6236 82220
rect 5540 80640 5592 80646
rect 5540 80582 5592 80588
rect 5552 79529 5580 80582
rect 5538 79520 5594 79529
rect 5538 79455 5594 79464
rect 6196 73574 6224 82214
rect 7116 77994 7144 93094
rect 7300 78674 7328 99622
rect 7484 95674 7512 99962
rect 7472 95668 7524 95674
rect 7472 95610 7524 95616
rect 7484 94994 7512 95610
rect 7472 94988 7524 94994
rect 7472 94930 7524 94936
rect 7484 94450 7512 94930
rect 7472 94444 7524 94450
rect 7472 94386 7524 94392
rect 7484 93838 7512 94386
rect 7472 93832 7524 93838
rect 7472 93774 7524 93780
rect 7484 93158 7512 93774
rect 7472 93152 7524 93158
rect 7472 93094 7524 93100
rect 7484 79937 7512 93094
rect 7564 88868 7616 88874
rect 7564 88810 7616 88816
rect 7470 79928 7526 79937
rect 7470 79863 7526 79872
rect 7576 79830 7604 88810
rect 7564 79824 7616 79830
rect 7564 79766 7616 79772
rect 7288 78668 7340 78674
rect 7288 78610 7340 78616
rect 7104 77988 7156 77994
rect 7104 77930 7156 77936
rect 8036 77722 8064 135730
rect 8116 135584 8168 135590
rect 8116 135526 8168 135532
rect 8024 77716 8076 77722
rect 8024 77658 8076 77664
rect 8128 77178 8156 135526
rect 8116 77172 8168 77178
rect 8116 77114 8168 77120
rect 8220 76974 8248 135798
rect 8944 134632 8996 134638
rect 8944 134574 8996 134580
rect 8956 93770 8984 134574
rect 9036 134564 9088 134570
rect 9036 134506 9088 134512
rect 9048 101114 9076 134506
rect 9496 111376 9548 111382
rect 9496 111318 9548 111324
rect 9508 111261 9536 111318
rect 9494 111252 9550 111261
rect 9494 111187 9550 111196
rect 9494 109552 9550 109561
rect 9494 109488 9496 109496
rect 9548 109488 9550 109496
rect 9494 109487 9550 109488
rect 9496 109482 9548 109487
rect 9496 108452 9548 108458
rect 9494 108424 9496 108433
rect 9548 108424 9550 108433
rect 9494 108359 9550 108368
rect 9496 107024 9548 107030
rect 9496 106966 9548 106972
rect 9508 106733 9536 106966
rect 9494 106724 9550 106733
rect 9494 106659 9550 106668
rect 9496 105936 9548 105942
rect 9496 105878 9548 105884
rect 9508 105650 9536 105878
rect 9494 105641 9550 105650
rect 9494 105576 9550 105585
rect 9496 104100 9548 104106
rect 9496 104042 9548 104048
rect 9508 103970 9536 104042
rect 9494 103961 9550 103970
rect 9494 103896 9550 103905
rect 9128 102196 9180 102202
rect 9128 102138 9180 102144
rect 9036 101108 9088 101114
rect 9036 101050 9088 101056
rect 8944 93764 8996 93770
rect 8944 93706 8996 93712
rect 8944 87780 8996 87786
rect 8944 87722 8996 87728
rect 8392 86692 8444 86698
rect 8392 86634 8444 86640
rect 8404 79665 8432 86634
rect 8576 85604 8628 85610
rect 8576 85546 8628 85552
rect 8390 79656 8446 79665
rect 8588 79626 8616 85546
rect 8956 79694 8984 87722
rect 8944 79688 8996 79694
rect 8944 79630 8996 79636
rect 8390 79591 8446 79600
rect 8576 79620 8628 79626
rect 8576 79562 8628 79568
rect 8208 76968 8260 76974
rect 8208 76910 8260 76916
rect 9140 76906 9168 102138
rect 9600 84194 9628 135866
rect 34164 134638 34192 136138
rect 34152 134632 34204 134638
rect 34152 134574 34204 134580
rect 34992 134570 35020 136138
rect 35594 136028 35902 136037
rect 35594 136026 35600 136028
rect 35656 136026 35680 136028
rect 35736 136026 35760 136028
rect 35816 136026 35840 136028
rect 35896 136026 35902 136028
rect 35656 135974 35658 136026
rect 35838 135974 35840 136026
rect 35594 135972 35600 135974
rect 35656 135972 35680 135974
rect 35736 135972 35760 135974
rect 35816 135972 35840 135974
rect 35896 135972 35902 135974
rect 35594 135963 35902 135972
rect 34980 134564 35032 134570
rect 34980 134506 35032 134512
rect 36004 133906 36032 136206
rect 36084 136128 36136 136134
rect 36084 136070 36136 136076
rect 36096 135794 36124 136070
rect 36084 135788 36136 135794
rect 36084 135730 36136 135736
rect 38580 133929 38608 136206
rect 38752 136196 38804 136202
rect 38752 136138 38804 136144
rect 43168 136196 43220 136202
rect 43168 136138 43220 136144
rect 48504 136196 48556 136202
rect 48504 136138 48556 136144
rect 51080 136196 51132 136202
rect 51080 136138 51132 136144
rect 55404 136196 55456 136202
rect 55404 136138 55456 136144
rect 57980 136196 58032 136202
rect 57980 136138 58032 136144
rect 60556 136196 60608 136202
rect 60556 136138 60608 136144
rect 63132 136196 63184 136202
rect 63132 136138 63184 136144
rect 38764 134201 38792 136138
rect 43076 136128 43128 136134
rect 43076 136070 43128 136076
rect 43088 135862 43116 136070
rect 43076 135856 43128 135862
rect 43076 135798 43128 135804
rect 43180 134201 43208 136138
rect 46112 136128 46164 136134
rect 46112 136070 46164 136076
rect 47676 136128 47728 136134
rect 47676 136070 47728 136076
rect 38750 134192 38806 134201
rect 38750 134127 38806 134136
rect 43166 134192 43222 134201
rect 43166 134127 43222 134136
rect 46124 133929 46152 136070
rect 47688 135930 47716 136070
rect 47676 135924 47728 135930
rect 47676 135866 47728 135872
rect 48516 133929 48544 136138
rect 50252 136128 50304 136134
rect 50252 136070 50304 136076
rect 50264 135590 50292 136070
rect 50252 135584 50304 135590
rect 50252 135526 50304 135532
rect 51092 133929 51120 136138
rect 55416 134201 55444 136138
rect 55772 136128 55824 136134
rect 55772 136070 55824 136076
rect 55784 135930 55812 136070
rect 55772 135924 55824 135930
rect 55772 135866 55824 135872
rect 57992 134201 58020 136138
rect 58348 136128 58400 136134
rect 58348 136070 58400 136076
rect 58360 135862 58388 136070
rect 58348 135856 58400 135862
rect 58348 135798 58400 135804
rect 60568 135289 60596 136138
rect 60924 136128 60976 136134
rect 60924 136070 60976 136076
rect 60936 135794 60964 136070
rect 60924 135788 60976 135794
rect 60924 135730 60976 135736
rect 63144 135289 63172 136138
rect 63604 136134 63632 136614
rect 65654 136572 65962 136581
rect 65654 136570 65660 136572
rect 65716 136570 65740 136572
rect 65796 136570 65820 136572
rect 65876 136570 65900 136572
rect 65956 136570 65962 136572
rect 65716 136518 65718 136570
rect 65898 136518 65900 136570
rect 65654 136516 65660 136518
rect 65716 136516 65740 136518
rect 65796 136516 65820 136518
rect 65876 136516 65900 136518
rect 65956 136516 65962 136518
rect 65654 136507 65962 136516
rect 72516 136196 72568 136202
rect 72516 136138 72568 136144
rect 72700 136196 72752 136202
rect 72700 136138 72752 136144
rect 77392 136196 77444 136202
rect 77392 136138 77444 136144
rect 63500 136128 63552 136134
rect 63500 136070 63552 136076
rect 63592 136128 63644 136134
rect 63592 136070 63644 136076
rect 68560 136128 68612 136134
rect 68560 136070 68612 136076
rect 63512 135726 63540 136070
rect 63500 135720 63552 135726
rect 63500 135662 63552 135668
rect 60554 135280 60610 135289
rect 60554 135215 60610 135224
rect 63130 135280 63186 135289
rect 63130 135215 63186 135224
rect 63604 135153 63632 136070
rect 66314 136028 66622 136037
rect 66314 136026 66320 136028
rect 66376 136026 66400 136028
rect 66456 136026 66480 136028
rect 66536 136026 66560 136028
rect 66616 136026 66622 136028
rect 66376 135974 66378 136026
rect 66558 135974 66560 136026
rect 66314 135972 66320 135974
rect 66376 135972 66400 135974
rect 66456 135972 66480 135974
rect 66536 135972 66560 135974
rect 66616 135972 66622 135974
rect 66314 135963 66622 135972
rect 63590 135144 63646 135153
rect 63590 135079 63646 135088
rect 55402 134192 55458 134201
rect 55402 134127 55458 134136
rect 57978 134192 58034 134201
rect 57978 134127 58034 134136
rect 68572 133929 68600 136070
rect 72528 134201 72556 136138
rect 72712 135289 72740 136138
rect 72884 136128 72936 136134
rect 72884 136070 72936 136076
rect 73804 136128 73856 136134
rect 73804 136070 73856 136076
rect 72896 135658 72924 136070
rect 72884 135652 72936 135658
rect 72884 135594 72936 135600
rect 73816 135590 73844 136070
rect 73804 135584 73856 135590
rect 73804 135526 73856 135532
rect 72698 135280 72754 135289
rect 72698 135215 72754 135224
rect 77404 134473 77432 136138
rect 95988 136134 96016 136614
rect 96374 136572 96682 136581
rect 96374 136570 96380 136572
rect 96436 136570 96460 136572
rect 96516 136570 96540 136572
rect 96596 136570 96620 136572
rect 96676 136570 96682 136572
rect 96436 136518 96438 136570
rect 96618 136518 96620 136570
rect 96374 136516 96380 136518
rect 96436 136516 96460 136518
rect 96516 136516 96540 136518
rect 96596 136516 96620 136518
rect 96676 136516 96682 136518
rect 96374 136507 96682 136516
rect 77760 136128 77812 136134
rect 77760 136070 77812 136076
rect 86316 136128 86368 136134
rect 86316 136070 86368 136076
rect 87328 136128 87380 136134
rect 87328 136070 87380 136076
rect 95976 136128 96028 136134
rect 95976 136070 96028 136076
rect 77772 135522 77800 136070
rect 77760 135516 77812 135522
rect 77760 135458 77812 135464
rect 86328 135454 86356 136070
rect 86316 135448 86368 135454
rect 86316 135390 86368 135396
rect 77390 134464 77446 134473
rect 77390 134399 77446 134408
rect 72514 134192 72570 134201
rect 72514 134127 72570 134136
rect 86328 133929 86356 135390
rect 87340 133958 87368 136070
rect 95988 135697 96016 136070
rect 97034 136028 97342 136037
rect 97034 136026 97040 136028
rect 97096 136026 97120 136028
rect 97176 136026 97200 136028
rect 97256 136026 97280 136028
rect 97336 136026 97342 136028
rect 97096 135974 97098 136026
rect 97278 135974 97280 136026
rect 97034 135972 97040 135974
rect 97096 135972 97120 135974
rect 97176 135972 97200 135974
rect 97256 135972 97280 135974
rect 97336 135972 97342 135974
rect 97034 135963 97342 135972
rect 95974 135688 96030 135697
rect 95974 135623 96030 135632
rect 87328 133952 87380 133958
rect 36082 133920 36138 133929
rect 36004 133878 36082 133906
rect 36082 133855 36138 133864
rect 38566 133920 38622 133929
rect 38566 133855 38622 133864
rect 46110 133920 46166 133929
rect 46110 133855 46166 133864
rect 48502 133920 48558 133929
rect 48502 133855 48558 133864
rect 51078 133920 51134 133929
rect 51078 133855 51134 133864
rect 68558 133920 68614 133929
rect 68558 133855 68614 133864
rect 86314 133920 86370 133929
rect 86314 133855 86370 133864
rect 87326 133920 87328 133929
rect 87380 133920 87382 133929
rect 87326 133855 87382 133864
rect 46124 133754 46152 133855
rect 68572 133754 68600 133855
rect 46112 133748 46164 133754
rect 46112 133690 46164 133696
rect 68560 133748 68612 133754
rect 68560 133690 68612 133696
rect 102046 92260 102102 92269
rect 102046 92195 102102 92204
rect 9312 84176 9364 84182
rect 9312 84118 9364 84124
rect 9416 84166 9628 84194
rect 9220 83496 9272 83502
rect 9220 83438 9272 83444
rect 9232 79121 9260 83438
rect 9324 79257 9352 84118
rect 9310 79248 9366 79257
rect 9310 79183 9366 79192
rect 9218 79112 9274 79121
rect 9218 79047 9274 79056
rect 9128 76900 9180 76906
rect 9128 76842 9180 76848
rect 9416 76634 9444 84166
rect 9772 81320 9824 81326
rect 9772 81262 9824 81268
rect 9588 81252 9640 81258
rect 9588 81194 9640 81200
rect 9600 79801 9628 81194
rect 9680 80844 9732 80850
rect 9680 80786 9732 80792
rect 9586 79792 9642 79801
rect 9692 79762 9720 80786
rect 9784 79966 9812 81262
rect 9864 80776 9916 80782
rect 9864 80718 9916 80724
rect 9772 79960 9824 79966
rect 9772 79902 9824 79908
rect 9876 79898 9904 80718
rect 9956 80708 10008 80714
rect 9956 80650 10008 80656
rect 9968 80034 9996 80650
rect 101956 80096 102008 80102
rect 101956 80038 102008 80044
rect 9956 80028 10008 80034
rect 9956 79970 10008 79976
rect 43260 80028 43312 80034
rect 43260 79970 43312 79976
rect 40960 79960 41012 79966
rect 16118 79928 16174 79937
rect 9864 79892 9916 79898
rect 16118 79863 16174 79872
rect 23478 79928 23534 79937
rect 23478 79863 23534 79872
rect 36266 79928 36322 79937
rect 36266 79863 36322 79872
rect 39762 79928 39818 79937
rect 39762 79863 39764 79872
rect 9864 79834 9916 79840
rect 9586 79727 9642 79736
rect 9680 79756 9732 79762
rect 9680 79698 9732 79704
rect 14004 78668 14056 78674
rect 14004 78610 14056 78616
rect 11060 77648 11112 77654
rect 11060 77590 11112 77596
rect 9404 76628 9456 76634
rect 9404 76570 9456 76576
rect 11072 75954 11100 77590
rect 14016 76498 14044 78610
rect 16132 77722 16160 79863
rect 16212 78056 16264 78062
rect 16212 77998 16264 78004
rect 16120 77716 16172 77722
rect 16120 77658 16172 77664
rect 16224 77450 16252 77998
rect 17132 77988 17184 77994
rect 17132 77930 17184 77936
rect 16212 77444 16264 77450
rect 16212 77386 16264 77392
rect 14648 77376 14700 77382
rect 14648 77318 14700 77324
rect 14004 76492 14056 76498
rect 14004 76434 14056 76440
rect 14556 76424 14608 76430
rect 14556 76366 14608 76372
rect 14568 75954 14596 76366
rect 14660 76090 14688 77318
rect 17144 76430 17172 77930
rect 19892 77512 19944 77518
rect 19892 77454 19944 77460
rect 19340 76560 19392 76566
rect 19340 76502 19392 76508
rect 17132 76424 17184 76430
rect 17132 76366 17184 76372
rect 16316 76090 16620 76106
rect 14648 76084 14700 76090
rect 14648 76026 14700 76032
rect 16316 76084 16632 76090
rect 16316 76078 16580 76084
rect 16316 76022 16344 76078
rect 16580 76026 16632 76032
rect 16304 76016 16356 76022
rect 16304 75958 16356 75964
rect 11060 75948 11112 75954
rect 11060 75890 11112 75896
rect 14556 75948 14608 75954
rect 14556 75890 14608 75896
rect 18052 75880 18104 75886
rect 18052 75822 18104 75828
rect 18064 75002 18092 75822
rect 19352 75818 19380 76502
rect 19340 75812 19392 75818
rect 19340 75754 19392 75760
rect 18144 75336 18196 75342
rect 18144 75278 18196 75284
rect 18052 74996 18104 75002
rect 18052 74938 18104 74944
rect 18156 74798 18184 75278
rect 19156 75268 19208 75274
rect 19156 75210 19208 75216
rect 18972 74996 19024 75002
rect 18972 74938 19024 74944
rect 18144 74792 18196 74798
rect 18144 74734 18196 74740
rect 9588 73908 9640 73914
rect 9588 73850 9640 73856
rect 6184 73568 6236 73574
rect 6184 73510 6236 73516
rect 5264 70916 5316 70922
rect 5264 70858 5316 70864
rect 4874 70748 5182 70757
rect 4874 70746 4880 70748
rect 4936 70746 4960 70748
rect 5016 70746 5040 70748
rect 5096 70746 5120 70748
rect 5176 70746 5182 70748
rect 4936 70694 4938 70746
rect 5118 70694 5120 70746
rect 4874 70692 4880 70694
rect 4936 70692 4960 70694
rect 5016 70692 5040 70694
rect 5096 70692 5120 70694
rect 5176 70692 5182 70694
rect 4874 70683 5182 70692
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70139 4522 70148
rect 4874 69660 5182 69669
rect 4874 69658 4880 69660
rect 4936 69658 4960 69660
rect 5016 69658 5040 69660
rect 5096 69658 5120 69660
rect 5176 69658 5182 69660
rect 4936 69606 4938 69658
rect 5118 69606 5120 69658
rect 4874 69604 4880 69606
rect 4936 69604 4960 69606
rect 5016 69604 5040 69606
rect 5096 69604 5120 69606
rect 5176 69604 5182 69606
rect 4874 69595 5182 69604
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 4874 68572 5182 68581
rect 4874 68570 4880 68572
rect 4936 68570 4960 68572
rect 5016 68570 5040 68572
rect 5096 68570 5120 68572
rect 5176 68570 5182 68572
rect 4936 68518 4938 68570
rect 5118 68518 5120 68570
rect 4874 68516 4880 68518
rect 4936 68516 4960 68518
rect 5016 68516 5040 68518
rect 5096 68516 5120 68518
rect 5176 68516 5182 68518
rect 4874 68507 5182 68516
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 4874 67484 5182 67493
rect 4874 67482 4880 67484
rect 4936 67482 4960 67484
rect 5016 67482 5040 67484
rect 5096 67482 5120 67484
rect 5176 67482 5182 67484
rect 4936 67430 4938 67482
rect 5118 67430 5120 67482
rect 4874 67428 4880 67430
rect 4936 67428 4960 67430
rect 5016 67428 5040 67430
rect 5096 67428 5120 67430
rect 5176 67428 5182 67430
rect 4874 67419 5182 67428
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 4874 66396 5182 66405
rect 4874 66394 4880 66396
rect 4936 66394 4960 66396
rect 5016 66394 5040 66396
rect 5096 66394 5120 66396
rect 5176 66394 5182 66396
rect 4936 66342 4938 66394
rect 5118 66342 5120 66394
rect 4874 66340 4880 66342
rect 4936 66340 4960 66342
rect 5016 66340 5040 66342
rect 5096 66340 5120 66342
rect 5176 66340 5182 66342
rect 4874 66331 5182 66340
rect 9496 66224 9548 66230
rect 9496 66166 9548 66172
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 4874 65308 5182 65317
rect 4874 65306 4880 65308
rect 4936 65306 4960 65308
rect 5016 65306 5040 65308
rect 5096 65306 5120 65308
rect 5176 65306 5182 65308
rect 4936 65254 4938 65306
rect 5118 65254 5120 65306
rect 4874 65252 4880 65254
rect 4936 65252 4960 65254
rect 5016 65252 5040 65254
rect 5096 65252 5120 65254
rect 5176 65252 5182 65254
rect 4874 65243 5182 65252
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 4874 64220 5182 64229
rect 4874 64218 4880 64220
rect 4936 64218 4960 64220
rect 5016 64218 5040 64220
rect 5096 64218 5120 64220
rect 5176 64218 5182 64220
rect 4936 64166 4938 64218
rect 5118 64166 5120 64218
rect 4874 64164 4880 64166
rect 4936 64164 4960 64166
rect 5016 64164 5040 64166
rect 5096 64164 5120 64166
rect 5176 64164 5182 64166
rect 4874 64155 5182 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 4874 63132 5182 63141
rect 4874 63130 4880 63132
rect 4936 63130 4960 63132
rect 5016 63130 5040 63132
rect 5096 63130 5120 63132
rect 5176 63130 5182 63132
rect 4936 63078 4938 63130
rect 5118 63078 5120 63130
rect 4874 63076 4880 63078
rect 4936 63076 4960 63078
rect 5016 63076 5040 63078
rect 5096 63076 5120 63078
rect 5176 63076 5182 63078
rect 4874 63067 5182 63076
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 4874 62044 5182 62053
rect 4874 62042 4880 62044
rect 4936 62042 4960 62044
rect 5016 62042 5040 62044
rect 5096 62042 5120 62044
rect 5176 62042 5182 62044
rect 4936 61990 4938 62042
rect 5118 61990 5120 62042
rect 4874 61988 4880 61990
rect 4936 61988 4960 61990
rect 5016 61988 5040 61990
rect 5096 61988 5120 61990
rect 5176 61988 5182 61990
rect 4874 61979 5182 61988
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4874 60956 5182 60965
rect 4874 60954 4880 60956
rect 4936 60954 4960 60956
rect 5016 60954 5040 60956
rect 5096 60954 5120 60956
rect 5176 60954 5182 60956
rect 4936 60902 4938 60954
rect 5118 60902 5120 60954
rect 4874 60900 4880 60902
rect 4936 60900 4960 60902
rect 5016 60900 5040 60902
rect 5096 60900 5120 60902
rect 5176 60900 5182 60902
rect 4874 60891 5182 60900
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 4874 59868 5182 59877
rect 4874 59866 4880 59868
rect 4936 59866 4960 59868
rect 5016 59866 5040 59868
rect 5096 59866 5120 59868
rect 5176 59866 5182 59868
rect 4936 59814 4938 59866
rect 5118 59814 5120 59866
rect 4874 59812 4880 59814
rect 4936 59812 4960 59814
rect 5016 59812 5040 59814
rect 5096 59812 5120 59814
rect 5176 59812 5182 59814
rect 4874 59803 5182 59812
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4874 58780 5182 58789
rect 4874 58778 4880 58780
rect 4936 58778 4960 58780
rect 5016 58778 5040 58780
rect 5096 58778 5120 58780
rect 5176 58778 5182 58780
rect 4936 58726 4938 58778
rect 5118 58726 5120 58778
rect 4874 58724 4880 58726
rect 4936 58724 4960 58726
rect 5016 58724 5040 58726
rect 5096 58724 5120 58726
rect 5176 58724 5182 58726
rect 4874 58715 5182 58724
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 7564 41472 7616 41478
rect 7564 41414 7616 41420
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 7576 41313 7604 41414
rect 7562 41304 7618 41313
rect 7562 41239 7618 41248
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 7576 40050 7604 41239
rect 3424 40044 3476 40050
rect 3424 39986 3476 39992
rect 7564 40044 7616 40050
rect 7564 39986 7616 39992
rect 1584 33108 1636 33114
rect 1584 33050 1636 33056
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1504 13705 1532 13874
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1308 13252 1360 13258
rect 1308 13194 1360 13200
rect 1320 13025 1348 13194
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1504 12345 1532 12786
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1216 11756 1268 11762
rect 1216 11698 1268 11704
rect 1228 11665 1256 11698
rect 1214 11656 1270 11665
rect 1214 11591 1270 11600
rect 1492 11076 1544 11082
rect 1492 11018 1544 11024
rect 1504 10985 1532 11018
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1596 10810 1624 33050
rect 1768 30320 1820 30326
rect 1768 30262 1820 30268
rect 1780 11898 1808 30262
rect 1860 26308 1912 26314
rect 1860 26250 1912 26256
rect 1872 12986 1900 26250
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 2056 13530 2084 24006
rect 3436 14074 3464 39986
rect 7288 39840 7340 39846
rect 7288 39782 7340 39788
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 7300 39545 7328 39782
rect 7286 39536 7342 39545
rect 7286 39471 7342 39480
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 7300 11354 7328 39471
rect 7564 38752 7616 38758
rect 7564 38694 7616 38700
rect 7576 38457 7604 38694
rect 7562 38448 7618 38457
rect 7618 38406 7696 38434
rect 7562 38383 7618 38392
rect 7562 36680 7618 36689
rect 7562 36615 7564 36624
rect 7616 36615 7618 36624
rect 7564 36586 7616 36592
rect 7576 36394 7604 36586
rect 7392 36366 7604 36394
rect 7392 26314 7420 36366
rect 7470 35592 7526 35601
rect 7470 35527 7526 35536
rect 7484 35494 7512 35527
rect 7472 35488 7524 35494
rect 7472 35430 7524 35436
rect 7484 30326 7512 35430
rect 7562 33960 7618 33969
rect 7562 33895 7564 33904
rect 7616 33895 7618 33904
rect 7564 33866 7616 33872
rect 7576 33114 7604 33866
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7472 30320 7524 30326
rect 7472 30262 7524 30268
rect 7380 26308 7432 26314
rect 7380 26250 7432 26256
rect 7668 26234 7696 38406
rect 7576 26206 7696 26234
rect 7576 24070 7604 26206
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7470 15464 7526 15473
rect 7470 15399 7526 15408
rect 7484 15366 7512 15399
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10305 1348 10610
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 1306 10296 1362 10305
rect 4214 10299 4522 10308
rect 1306 10231 1362 10240
rect 1492 9988 1544 9994
rect 1492 9930 1544 9936
rect 1504 9625 1532 9930
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 1214 8936 1270 8945
rect 1214 8871 1216 8880
rect 1268 8871 1270 8880
rect 1216 8842 1268 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1950 8256 2006 8265
rect 2056 8242 2084 8366
rect 2006 8214 2084 8242
rect 1950 8191 2006 8200
rect 1964 8090 1992 8191
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 1320 7585 1348 7754
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 1306 7576 1362 7585
rect 4874 7579 5182 7588
rect 1306 7511 1362 7520
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1320 6905 1348 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1306 6896 1362 6905
rect 1306 6831 1362 6840
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 1216 6316 1268 6322
rect 1216 6258 1268 6264
rect 1228 6225 1256 6258
rect 1214 6216 1270 6225
rect 1214 6151 1270 6160
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 7484 5914 7512 15302
rect 9508 9654 9536 66166
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9600 9586 9628 73850
rect 18984 73778 19012 74938
rect 19168 74934 19196 75210
rect 19904 75002 19932 77454
rect 23492 77382 23520 79863
rect 36280 79830 36308 79863
rect 39816 79863 39818 79872
rect 40958 79928 40960 79937
rect 43272 79937 43300 79970
rect 41012 79928 41014 79937
rect 40958 79863 41014 79872
rect 43258 79928 43314 79937
rect 43258 79863 43314 79872
rect 39764 79834 39816 79840
rect 36268 79824 36320 79830
rect 36268 79766 36320 79772
rect 38658 79792 38714 79801
rect 33968 79688 34020 79694
rect 30470 79656 30526 79665
rect 30470 79591 30526 79600
rect 31666 79656 31722 79665
rect 33968 79630 34020 79636
rect 31666 79591 31668 79600
rect 24674 79520 24730 79529
rect 24674 79455 24730 79464
rect 26054 79520 26110 79529
rect 26054 79455 26110 79464
rect 26974 79520 27030 79529
rect 26974 79455 27030 79464
rect 28170 79520 28226 79529
rect 28170 79455 28226 79464
rect 29550 79520 29606 79529
rect 29550 79455 29606 79464
rect 20720 77376 20772 77382
rect 20720 77318 20772 77324
rect 23480 77376 23532 77382
rect 23480 77318 23532 77324
rect 20732 77110 20760 77318
rect 20720 77104 20772 77110
rect 20720 77046 20772 77052
rect 22468 77036 22520 77042
rect 22468 76978 22520 76984
rect 22480 76922 22508 76978
rect 22388 76894 22508 76922
rect 22388 76838 22416 76894
rect 22376 76832 22428 76838
rect 22376 76774 22428 76780
rect 22284 76084 22336 76090
rect 22284 76026 22336 76032
rect 22296 75546 22324 76026
rect 22284 75540 22336 75546
rect 22284 75482 22336 75488
rect 22388 75342 22416 76774
rect 22376 75336 22428 75342
rect 22376 75278 22428 75284
rect 22388 75206 22416 75278
rect 22376 75200 22428 75206
rect 22376 75142 22428 75148
rect 19892 74996 19944 75002
rect 19892 74938 19944 74944
rect 19156 74928 19208 74934
rect 19156 74870 19208 74876
rect 19904 74866 19932 74938
rect 19892 74860 19944 74866
rect 19892 74802 19944 74808
rect 23388 74180 23440 74186
rect 23388 74122 23440 74128
rect 23400 73846 23428 74122
rect 23388 73840 23440 73846
rect 23388 73782 23440 73788
rect 18972 73772 19024 73778
rect 18972 73714 19024 73720
rect 11704 73704 11756 73710
rect 11704 73646 11756 73652
rect 11716 72690 11744 73646
rect 13820 73636 13872 73642
rect 13820 73578 13872 73584
rect 11704 72684 11756 72690
rect 11704 72626 11756 72632
rect 13832 66230 13860 73578
rect 18984 73574 19012 73714
rect 18972 73568 19024 73574
rect 18972 73510 19024 73516
rect 22928 73568 22980 73574
rect 22928 73510 22980 73516
rect 22940 73234 22968 73510
rect 22928 73228 22980 73234
rect 22928 73170 22980 73176
rect 23492 71398 23520 77318
rect 24688 77110 24716 79455
rect 25412 78056 25464 78062
rect 25412 77998 25464 78004
rect 24676 77104 24728 77110
rect 24676 77046 24728 77052
rect 25228 77104 25280 77110
rect 25228 77046 25280 77052
rect 25240 76906 25268 77046
rect 25228 76900 25280 76906
rect 25228 76842 25280 76848
rect 25424 76838 25452 77998
rect 26068 77926 26096 79455
rect 26988 79257 27016 79455
rect 26974 79248 27030 79257
rect 26974 79183 27030 79192
rect 26056 77920 26108 77926
rect 26056 77862 26108 77868
rect 26068 77722 26096 77862
rect 26988 77722 27016 79183
rect 28184 79121 28212 79455
rect 28170 79112 28226 79121
rect 28170 79047 28226 79056
rect 28184 77722 28212 79047
rect 29564 78470 29592 79455
rect 29552 78464 29604 78470
rect 29552 78406 29604 78412
rect 29564 77722 29592 78406
rect 30484 77722 30512 79591
rect 31720 79591 31722 79600
rect 31668 79562 31720 79568
rect 31680 78962 31708 79562
rect 33980 79529 34008 79630
rect 33966 79520 34022 79529
rect 33966 79455 34022 79464
rect 35346 79520 35402 79529
rect 35346 79455 35402 79464
rect 32862 79112 32918 79121
rect 32862 79047 32918 79056
rect 31680 78934 31800 78962
rect 31772 77722 31800 78934
rect 32876 77722 32904 79047
rect 33980 77722 34008 79455
rect 35360 78130 35388 79455
rect 35348 78124 35400 78130
rect 35348 78066 35400 78072
rect 34934 77820 35242 77829
rect 34934 77818 34940 77820
rect 34996 77818 35020 77820
rect 35076 77818 35100 77820
rect 35156 77818 35180 77820
rect 35236 77818 35242 77820
rect 34996 77766 34998 77818
rect 35178 77766 35180 77818
rect 34934 77764 34940 77766
rect 34996 77764 35020 77766
rect 35076 77764 35100 77766
rect 35156 77764 35180 77766
rect 35236 77764 35242 77766
rect 34934 77755 35242 77764
rect 35360 77722 35388 78066
rect 36280 77722 36308 79766
rect 38658 79727 38660 79736
rect 38712 79727 38714 79736
rect 38660 79698 38712 79704
rect 37462 79656 37518 79665
rect 37462 79591 37518 79600
rect 37476 79558 37504 79591
rect 37464 79552 37516 79558
rect 37464 79494 37516 79500
rect 37476 77722 37504 79494
rect 38672 77722 38700 79698
rect 39776 77722 39804 79834
rect 40972 77722 41000 79863
rect 42154 79520 42210 79529
rect 42154 79455 42210 79464
rect 42168 79014 42196 79455
rect 42156 79008 42208 79014
rect 42156 78950 42208 78956
rect 42168 77722 42196 78950
rect 43272 77722 43300 79863
rect 98000 79688 98052 79694
rect 98000 79630 98052 79636
rect 92112 79484 92164 79490
rect 92112 79426 92164 79432
rect 90272 79416 90324 79422
rect 90272 79358 90324 79364
rect 73804 79348 73856 79354
rect 73804 79290 73856 79296
rect 65654 77820 65962 77829
rect 65654 77818 65660 77820
rect 65716 77818 65740 77820
rect 65796 77818 65820 77820
rect 65876 77818 65900 77820
rect 65956 77818 65962 77820
rect 65716 77766 65718 77818
rect 65898 77766 65900 77818
rect 65654 77764 65660 77766
rect 65716 77764 65740 77766
rect 65796 77764 65820 77766
rect 65876 77764 65900 77766
rect 65956 77764 65962 77766
rect 65654 77755 65962 77764
rect 26056 77716 26108 77722
rect 26056 77658 26108 77664
rect 26976 77716 27028 77722
rect 26976 77658 27028 77664
rect 28172 77716 28224 77722
rect 28172 77658 28224 77664
rect 29552 77716 29604 77722
rect 29552 77658 29604 77664
rect 30472 77716 30524 77722
rect 30472 77658 30524 77664
rect 31760 77716 31812 77722
rect 31760 77658 31812 77664
rect 32864 77716 32916 77722
rect 32864 77658 32916 77664
rect 33968 77716 34020 77722
rect 33968 77658 34020 77664
rect 35348 77716 35400 77722
rect 35348 77658 35400 77664
rect 36268 77716 36320 77722
rect 36268 77658 36320 77664
rect 37464 77716 37516 77722
rect 37464 77658 37516 77664
rect 38660 77716 38712 77722
rect 38660 77658 38712 77664
rect 39764 77716 39816 77722
rect 39764 77658 39816 77664
rect 40960 77716 41012 77722
rect 40960 77658 41012 77664
rect 42156 77716 42208 77722
rect 42156 77658 42208 77664
rect 43260 77716 43312 77722
rect 43260 77658 43312 77664
rect 27528 77648 27580 77654
rect 27528 77590 27580 77596
rect 26332 76968 26384 76974
rect 26332 76910 26384 76916
rect 26344 76838 26372 76910
rect 25412 76832 25464 76838
rect 25412 76774 25464 76780
rect 26332 76832 26384 76838
rect 26332 76774 26384 76780
rect 26344 76498 26372 76774
rect 27540 76498 27568 77590
rect 55036 77512 55088 77518
rect 55036 77454 55088 77460
rect 55048 77382 55076 77454
rect 55128 77444 55180 77450
rect 55128 77386 55180 77392
rect 55036 77376 55088 77382
rect 55036 77318 55088 77324
rect 35594 77276 35902 77285
rect 35594 77274 35600 77276
rect 35656 77274 35680 77276
rect 35736 77274 35760 77276
rect 35816 77274 35840 77276
rect 35896 77274 35902 77276
rect 35656 77222 35658 77274
rect 35838 77222 35840 77274
rect 35594 77220 35600 77222
rect 35656 77220 35680 77222
rect 35736 77220 35760 77222
rect 35816 77220 35840 77222
rect 35896 77220 35902 77222
rect 35594 77211 35902 77220
rect 46940 77172 46992 77178
rect 46940 77114 46992 77120
rect 32956 77036 33008 77042
rect 32956 76978 33008 76984
rect 26332 76492 26384 76498
rect 26332 76434 26384 76440
rect 27528 76492 27580 76498
rect 27528 76434 27580 76440
rect 30288 76356 30340 76362
rect 30288 76298 30340 76304
rect 23572 76288 23624 76294
rect 23572 76230 23624 76236
rect 24860 76288 24912 76294
rect 24860 76230 24912 76236
rect 28448 76288 28500 76294
rect 28448 76230 28500 76236
rect 28540 76288 28592 76294
rect 28540 76230 28592 76236
rect 23584 76090 23612 76230
rect 23572 76084 23624 76090
rect 23572 76026 23624 76032
rect 24768 75200 24820 75206
rect 24768 75142 24820 75148
rect 24780 74254 24808 75142
rect 24768 74248 24820 74254
rect 24768 74190 24820 74196
rect 24872 73794 24900 76230
rect 28264 74248 28316 74254
rect 28264 74190 28316 74196
rect 25044 74180 25096 74186
rect 25044 74122 25096 74128
rect 24688 73766 24900 73794
rect 24688 73710 24716 73766
rect 25056 73710 25084 74122
rect 28276 73778 28304 74190
rect 28264 73772 28316 73778
rect 28264 73714 28316 73720
rect 24676 73704 24728 73710
rect 24676 73646 24728 73652
rect 24768 73704 24820 73710
rect 24768 73646 24820 73652
rect 25044 73704 25096 73710
rect 25044 73646 25096 73652
rect 24780 73166 24808 73646
rect 25056 73370 25084 73646
rect 27896 73568 27948 73574
rect 27896 73510 27948 73516
rect 25044 73364 25096 73370
rect 25044 73306 25096 73312
rect 24768 73160 24820 73166
rect 24768 73102 24820 73108
rect 27908 73030 27936 73510
rect 27896 73024 27948 73030
rect 27896 72966 27948 72972
rect 23480 71392 23532 71398
rect 23480 71334 23532 71340
rect 28460 70582 28488 76230
rect 28552 74798 28580 76230
rect 28540 74792 28592 74798
rect 28540 74734 28592 74740
rect 29644 74112 29696 74118
rect 29644 74054 29696 74060
rect 29656 73846 29684 74054
rect 29644 73840 29696 73846
rect 29644 73782 29696 73788
rect 29368 73568 29420 73574
rect 29368 73510 29420 73516
rect 29380 73234 29408 73510
rect 29368 73228 29420 73234
rect 29368 73170 29420 73176
rect 30300 70854 30328 76298
rect 30564 76084 30616 76090
rect 30564 76026 30616 76032
rect 30288 70848 30340 70854
rect 30288 70790 30340 70796
rect 30576 70650 30604 76026
rect 31760 73704 31812 73710
rect 31760 73646 31812 73652
rect 31772 71194 31800 73646
rect 31760 71188 31812 71194
rect 31760 71130 31812 71136
rect 30564 70644 30616 70650
rect 30564 70586 30616 70592
rect 28448 70576 28500 70582
rect 28448 70518 28500 70524
rect 31668 70508 31720 70514
rect 31668 70450 31720 70456
rect 31680 69766 31708 70450
rect 31772 70394 31800 71130
rect 31852 70508 31904 70514
rect 31852 70450 31904 70456
rect 31864 70394 31892 70450
rect 31772 70366 31892 70394
rect 31864 70106 31892 70366
rect 31852 70100 31904 70106
rect 31852 70042 31904 70048
rect 32968 70038 32996 76978
rect 41328 76900 41380 76906
rect 41328 76842 41380 76848
rect 34934 76732 35242 76741
rect 34934 76730 34940 76732
rect 34996 76730 35020 76732
rect 35076 76730 35100 76732
rect 35156 76730 35180 76732
rect 35236 76730 35242 76732
rect 34996 76678 34998 76730
rect 35178 76678 35180 76730
rect 34934 76676 34940 76678
rect 34996 76676 35020 76678
rect 35076 76676 35100 76678
rect 35156 76676 35180 76678
rect 35236 76676 35242 76678
rect 34934 76667 35242 76676
rect 41340 76634 41368 76842
rect 46952 76634 46980 77114
rect 55048 76838 55076 77318
rect 55036 76832 55088 76838
rect 55036 76774 55088 76780
rect 41328 76628 41380 76634
rect 41328 76570 41380 76576
rect 46940 76628 46992 76634
rect 46940 76570 46992 76576
rect 41340 76294 41368 76570
rect 46952 76362 46980 76570
rect 55048 76430 55076 76774
rect 55036 76424 55088 76430
rect 55036 76366 55088 76372
rect 46940 76356 46992 76362
rect 46940 76298 46992 76304
rect 33048 76288 33100 76294
rect 33048 76230 33100 76236
rect 39856 76288 39908 76294
rect 39856 76230 39908 76236
rect 41328 76288 41380 76294
rect 41328 76230 41380 76236
rect 42892 76288 42944 76294
rect 42892 76230 42944 76236
rect 45468 76288 45520 76294
rect 45468 76230 45520 76236
rect 33060 73710 33088 76230
rect 35594 76188 35902 76197
rect 35594 76186 35600 76188
rect 35656 76186 35680 76188
rect 35736 76186 35760 76188
rect 35816 76186 35840 76188
rect 35896 76186 35902 76188
rect 35656 76134 35658 76186
rect 35838 76134 35840 76186
rect 35594 76132 35600 76134
rect 35656 76132 35680 76134
rect 35736 76132 35760 76134
rect 35816 76132 35840 76134
rect 35896 76132 35902 76134
rect 35594 76123 35902 76132
rect 34934 75644 35242 75653
rect 34934 75642 34940 75644
rect 34996 75642 35020 75644
rect 35076 75642 35100 75644
rect 35156 75642 35180 75644
rect 35236 75642 35242 75644
rect 34996 75590 34998 75642
rect 35178 75590 35180 75642
rect 34934 75588 34940 75590
rect 34996 75588 35020 75590
rect 35076 75588 35100 75590
rect 35156 75588 35180 75590
rect 35236 75588 35242 75590
rect 34934 75579 35242 75588
rect 35594 75100 35902 75109
rect 35594 75098 35600 75100
rect 35656 75098 35680 75100
rect 35736 75098 35760 75100
rect 35816 75098 35840 75100
rect 35896 75098 35902 75100
rect 35656 75046 35658 75098
rect 35838 75046 35840 75098
rect 35594 75044 35600 75046
rect 35656 75044 35680 75046
rect 35736 75044 35760 75046
rect 35816 75044 35840 75046
rect 35896 75044 35902 75046
rect 35594 75035 35902 75044
rect 34934 74556 35242 74565
rect 34934 74554 34940 74556
rect 34996 74554 35020 74556
rect 35076 74554 35100 74556
rect 35156 74554 35180 74556
rect 35236 74554 35242 74556
rect 34996 74502 34998 74554
rect 35178 74502 35180 74554
rect 34934 74500 34940 74502
rect 34996 74500 35020 74502
rect 35076 74500 35100 74502
rect 35156 74500 35180 74502
rect 35236 74500 35242 74502
rect 34934 74491 35242 74500
rect 35440 74452 35492 74458
rect 35440 74394 35492 74400
rect 33048 73704 33100 73710
rect 33048 73646 33100 73652
rect 34934 73468 35242 73477
rect 34934 73466 34940 73468
rect 34996 73466 35020 73468
rect 35076 73466 35100 73468
rect 35156 73466 35180 73468
rect 35236 73466 35242 73468
rect 34996 73414 34998 73466
rect 35178 73414 35180 73466
rect 34934 73412 34940 73414
rect 34996 73412 35020 73414
rect 35076 73412 35100 73414
rect 35156 73412 35180 73414
rect 35236 73412 35242 73414
rect 34934 73403 35242 73412
rect 35452 73030 35480 74394
rect 36176 74112 36228 74118
rect 36176 74054 36228 74060
rect 35594 74012 35902 74021
rect 35594 74010 35600 74012
rect 35656 74010 35680 74012
rect 35736 74010 35760 74012
rect 35816 74010 35840 74012
rect 35896 74010 35902 74012
rect 35656 73958 35658 74010
rect 35838 73958 35840 74010
rect 35594 73956 35600 73958
rect 35656 73956 35680 73958
rect 35736 73956 35760 73958
rect 35816 73956 35840 73958
rect 35896 73956 35902 73958
rect 35594 73947 35902 73956
rect 35440 73024 35492 73030
rect 35440 72966 35492 72972
rect 35594 72924 35902 72933
rect 35594 72922 35600 72924
rect 35656 72922 35680 72924
rect 35736 72922 35760 72924
rect 35816 72922 35840 72924
rect 35896 72922 35902 72924
rect 35656 72870 35658 72922
rect 35838 72870 35840 72922
rect 35594 72868 35600 72870
rect 35656 72868 35680 72870
rect 35736 72868 35760 72870
rect 35816 72868 35840 72870
rect 35896 72868 35902 72870
rect 35594 72859 35902 72868
rect 34934 72380 35242 72389
rect 34934 72378 34940 72380
rect 34996 72378 35020 72380
rect 35076 72378 35100 72380
rect 35156 72378 35180 72380
rect 35236 72378 35242 72380
rect 34996 72326 34998 72378
rect 35178 72326 35180 72378
rect 34934 72324 34940 72326
rect 34996 72324 35020 72326
rect 35076 72324 35100 72326
rect 35156 72324 35180 72326
rect 35236 72324 35242 72326
rect 34934 72315 35242 72324
rect 35594 71836 35902 71845
rect 35594 71834 35600 71836
rect 35656 71834 35680 71836
rect 35736 71834 35760 71836
rect 35816 71834 35840 71836
rect 35896 71834 35902 71836
rect 35656 71782 35658 71834
rect 35838 71782 35840 71834
rect 35594 71780 35600 71782
rect 35656 71780 35680 71782
rect 35736 71780 35760 71782
rect 35816 71780 35840 71782
rect 35896 71780 35902 71782
rect 35594 71771 35902 71780
rect 36188 71398 36216 74054
rect 39868 73914 39896 76230
rect 39856 73908 39908 73914
rect 39856 73850 39908 73856
rect 38844 73772 38896 73778
rect 38844 73714 38896 73720
rect 37924 73704 37976 73710
rect 37924 73646 37976 73652
rect 37936 73234 37964 73646
rect 37924 73228 37976 73234
rect 37924 73170 37976 73176
rect 37740 73024 37792 73030
rect 37740 72966 37792 72972
rect 37832 73024 37884 73030
rect 37832 72966 37884 72972
rect 37752 72758 37780 72966
rect 37844 72826 37872 72966
rect 37832 72820 37884 72826
rect 37832 72762 37884 72768
rect 37740 72752 37792 72758
rect 37740 72694 37792 72700
rect 36176 71392 36228 71398
rect 36176 71334 36228 71340
rect 34934 71292 35242 71301
rect 34934 71290 34940 71292
rect 34996 71290 35020 71292
rect 35076 71290 35100 71292
rect 35156 71290 35180 71292
rect 35236 71290 35242 71292
rect 34996 71238 34998 71290
rect 35178 71238 35180 71290
rect 34934 71236 34940 71238
rect 34996 71236 35020 71238
rect 35076 71236 35100 71238
rect 35156 71236 35180 71238
rect 35236 71236 35242 71238
rect 34934 71227 35242 71236
rect 34520 70848 34572 70854
rect 34520 70790 34572 70796
rect 34532 70650 34560 70790
rect 35594 70748 35902 70757
rect 35594 70746 35600 70748
rect 35656 70746 35680 70748
rect 35736 70746 35760 70748
rect 35816 70746 35840 70748
rect 35896 70746 35902 70748
rect 35656 70694 35658 70746
rect 35838 70694 35840 70746
rect 35594 70692 35600 70694
rect 35656 70692 35680 70694
rect 35736 70692 35760 70694
rect 35816 70692 35840 70694
rect 35896 70692 35902 70694
rect 35594 70683 35902 70692
rect 34520 70644 34572 70650
rect 34520 70586 34572 70592
rect 35532 70576 35584 70582
rect 35532 70518 35584 70524
rect 34520 70440 34572 70446
rect 34520 70382 34572 70388
rect 32956 70032 33008 70038
rect 32956 69974 33008 69980
rect 31668 69760 31720 69766
rect 31668 69702 31720 69708
rect 13820 66224 13872 66230
rect 13820 66166 13872 66172
rect 31680 65521 31708 69702
rect 34532 65657 34560 70382
rect 34934 70204 35242 70213
rect 34934 70202 34940 70204
rect 34996 70202 35020 70204
rect 35076 70202 35100 70204
rect 35156 70202 35180 70204
rect 35236 70202 35242 70204
rect 34996 70150 34998 70202
rect 35178 70150 35180 70202
rect 34934 70148 34940 70150
rect 34996 70148 35020 70150
rect 35076 70148 35100 70150
rect 35156 70148 35180 70150
rect 35236 70148 35242 70150
rect 34934 70139 35242 70148
rect 35544 70106 35572 70518
rect 35532 70100 35584 70106
rect 35532 70042 35584 70048
rect 38660 69964 38712 69970
rect 38660 69906 38712 69912
rect 35594 69660 35902 69669
rect 35594 69658 35600 69660
rect 35656 69658 35680 69660
rect 35736 69658 35760 69660
rect 35816 69658 35840 69660
rect 35896 69658 35902 69660
rect 35656 69606 35658 69658
rect 35838 69606 35840 69658
rect 35594 69604 35600 69606
rect 35656 69604 35680 69606
rect 35736 69604 35760 69606
rect 35816 69604 35840 69606
rect 35896 69604 35902 69606
rect 35594 69595 35902 69604
rect 34934 69116 35242 69125
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69051 35242 69060
rect 35594 68572 35902 68581
rect 35594 68570 35600 68572
rect 35656 68570 35680 68572
rect 35736 68570 35760 68572
rect 35816 68570 35840 68572
rect 35896 68570 35902 68572
rect 35656 68518 35658 68570
rect 35838 68518 35840 68570
rect 35594 68516 35600 68518
rect 35656 68516 35680 68518
rect 35736 68516 35760 68518
rect 35816 68516 35840 68518
rect 35896 68516 35902 68518
rect 35594 68507 35902 68516
rect 38672 68474 38700 69906
rect 38856 68474 38884 73714
rect 42708 73024 42760 73030
rect 42708 72966 42760 72972
rect 42432 72752 42484 72758
rect 42432 72694 42484 72700
rect 41144 70440 41196 70446
rect 41144 70382 41196 70388
rect 38660 68468 38712 68474
rect 38660 68410 38712 68416
rect 38844 68468 38896 68474
rect 38844 68410 38896 68416
rect 39948 68332 40000 68338
rect 39948 68274 40000 68280
rect 34934 68028 35242 68037
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67963 35242 67972
rect 35594 67484 35902 67493
rect 35594 67482 35600 67484
rect 35656 67482 35680 67484
rect 35736 67482 35760 67484
rect 35816 67482 35840 67484
rect 35896 67482 35902 67484
rect 35656 67430 35658 67482
rect 35838 67430 35840 67482
rect 35594 67428 35600 67430
rect 35656 67428 35680 67430
rect 35736 67428 35760 67430
rect 35816 67428 35840 67430
rect 35896 67428 35902 67430
rect 35594 67419 35902 67428
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 35594 66396 35902 66405
rect 35594 66394 35600 66396
rect 35656 66394 35680 66396
rect 35736 66394 35760 66396
rect 35816 66394 35840 66396
rect 35896 66394 35902 66396
rect 35656 66342 35658 66394
rect 35838 66342 35840 66394
rect 35594 66340 35600 66342
rect 35656 66340 35680 66342
rect 35736 66340 35760 66342
rect 35816 66340 35840 66342
rect 35896 66340 35902 66342
rect 35594 66331 35902 66340
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 34518 65648 34574 65657
rect 34518 65583 34574 65592
rect 31666 65512 31722 65521
rect 31666 65447 31722 65456
rect 39960 64161 39988 68274
rect 41156 64297 41184 70382
rect 42444 69562 42472 72694
rect 42432 69556 42484 69562
rect 42432 69498 42484 69504
rect 42156 69216 42208 69222
rect 42156 69158 42208 69164
rect 42168 68406 42196 69158
rect 42720 68950 42748 72966
rect 42904 72826 42932 76230
rect 45480 73166 45508 76230
rect 45468 73160 45520 73166
rect 45468 73102 45520 73108
rect 42892 72820 42944 72826
rect 42892 72762 42944 72768
rect 55140 71194 55168 77386
rect 59268 77376 59320 77382
rect 59268 77318 59320 77324
rect 59280 76634 59308 77318
rect 66314 77276 66622 77285
rect 66314 77274 66320 77276
rect 66376 77274 66400 77276
rect 66456 77274 66480 77276
rect 66536 77274 66560 77276
rect 66616 77274 66622 77276
rect 66376 77222 66378 77274
rect 66558 77222 66560 77274
rect 66314 77220 66320 77222
rect 66376 77220 66400 77222
rect 66456 77220 66480 77222
rect 66536 77220 66560 77222
rect 66616 77220 66622 77222
rect 66314 77211 66622 77220
rect 67914 77072 67970 77081
rect 67914 77007 67970 77016
rect 65982 76936 66038 76945
rect 65982 76871 66038 76880
rect 65654 76732 65962 76741
rect 65654 76730 65660 76732
rect 65716 76730 65740 76732
rect 65796 76730 65820 76732
rect 65876 76730 65900 76732
rect 65956 76730 65962 76732
rect 65716 76678 65718 76730
rect 65898 76678 65900 76730
rect 65654 76676 65660 76678
rect 65716 76676 65740 76678
rect 65796 76676 65820 76678
rect 65876 76676 65900 76678
rect 65956 76676 65962 76678
rect 65654 76667 65962 76676
rect 58624 76628 58676 76634
rect 58624 76570 58676 76576
rect 59268 76628 59320 76634
rect 59268 76570 59320 76576
rect 56140 73568 56192 73574
rect 56140 73510 56192 73516
rect 55128 71188 55180 71194
rect 55128 71130 55180 71136
rect 56152 70854 56180 73510
rect 56140 70848 56192 70854
rect 56140 70790 56192 70796
rect 45100 69828 45152 69834
rect 45100 69770 45152 69776
rect 43720 69420 43772 69426
rect 43720 69362 43772 69368
rect 42708 68944 42760 68950
rect 42708 68886 42760 68892
rect 43732 68746 43760 69362
rect 43812 69216 43864 69222
rect 43812 69158 43864 69164
rect 43824 69018 43852 69158
rect 43812 69012 43864 69018
rect 43812 68954 43864 68960
rect 43720 68740 43772 68746
rect 43720 68682 43772 68688
rect 42156 68400 42208 68406
rect 42156 68342 42208 68348
rect 43732 68241 43760 68682
rect 43718 68232 43774 68241
rect 43718 68167 43774 68176
rect 45112 65657 45140 69770
rect 58636 69018 58664 76570
rect 63130 76528 63186 76537
rect 63130 76463 63186 76472
rect 61014 76392 61070 76401
rect 63144 76362 63172 76463
rect 65996 76362 66024 76871
rect 67928 76362 67956 77007
rect 68928 76628 68980 76634
rect 68928 76570 68980 76576
rect 61014 76327 61016 76336
rect 61068 76327 61070 76336
rect 63132 76356 63184 76362
rect 61016 76298 61068 76304
rect 63132 76298 63184 76304
rect 65984 76356 66036 76362
rect 65984 76298 66036 76304
rect 67916 76356 67968 76362
rect 67916 76298 67968 76304
rect 62120 76288 62172 76294
rect 62120 76230 62172 76236
rect 64236 76288 64288 76294
rect 64236 76230 64288 76236
rect 62132 76090 62160 76230
rect 62120 76084 62172 76090
rect 62120 76026 62172 76032
rect 64248 76022 64276 76230
rect 66314 76188 66622 76197
rect 66314 76186 66320 76188
rect 66376 76186 66400 76188
rect 66456 76186 66480 76188
rect 66536 76186 66560 76188
rect 66616 76186 66622 76188
rect 66376 76134 66378 76186
rect 66558 76134 66560 76186
rect 66314 76132 66320 76134
rect 66376 76132 66400 76134
rect 66456 76132 66480 76134
rect 66536 76132 66560 76134
rect 66616 76132 66622 76134
rect 66314 76123 66622 76132
rect 68468 76084 68520 76090
rect 68468 76026 68520 76032
rect 64236 76016 64288 76022
rect 64236 75958 64288 75964
rect 65654 75644 65962 75653
rect 65654 75642 65660 75644
rect 65716 75642 65740 75644
rect 65796 75642 65820 75644
rect 65876 75642 65900 75644
rect 65956 75642 65962 75644
rect 65716 75590 65718 75642
rect 65898 75590 65900 75642
rect 65654 75588 65660 75590
rect 65716 75588 65740 75590
rect 65796 75588 65820 75590
rect 65876 75588 65900 75590
rect 65956 75588 65962 75590
rect 65654 75579 65962 75588
rect 66314 75100 66622 75109
rect 66314 75098 66320 75100
rect 66376 75098 66400 75100
rect 66456 75098 66480 75100
rect 66536 75098 66560 75100
rect 66616 75098 66622 75100
rect 66376 75046 66378 75098
rect 66558 75046 66560 75098
rect 66314 75044 66320 75046
rect 66376 75044 66400 75046
rect 66456 75044 66480 75046
rect 66536 75044 66560 75046
rect 66616 75044 66622 75046
rect 66314 75035 66622 75044
rect 65654 74556 65962 74565
rect 65654 74554 65660 74556
rect 65716 74554 65740 74556
rect 65796 74554 65820 74556
rect 65876 74554 65900 74556
rect 65956 74554 65962 74556
rect 65716 74502 65718 74554
rect 65898 74502 65900 74554
rect 65654 74500 65660 74502
rect 65716 74500 65740 74502
rect 65796 74500 65820 74502
rect 65876 74500 65900 74502
rect 65956 74500 65962 74502
rect 65654 74491 65962 74500
rect 66314 74012 66622 74021
rect 66314 74010 66320 74012
rect 66376 74010 66400 74012
rect 66456 74010 66480 74012
rect 66536 74010 66560 74012
rect 66616 74010 66622 74012
rect 66376 73958 66378 74010
rect 66558 73958 66560 74010
rect 66314 73956 66320 73958
rect 66376 73956 66400 73958
rect 66456 73956 66480 73958
rect 66536 73956 66560 73958
rect 66616 73956 66622 73958
rect 66314 73947 66622 73956
rect 68480 73914 68508 76026
rect 68468 73908 68520 73914
rect 68468 73850 68520 73856
rect 68560 73772 68612 73778
rect 68560 73714 68612 73720
rect 68284 73704 68336 73710
rect 68284 73646 68336 73652
rect 65654 73468 65962 73477
rect 65654 73466 65660 73468
rect 65716 73466 65740 73468
rect 65796 73466 65820 73468
rect 65876 73466 65900 73468
rect 65956 73466 65962 73468
rect 65716 73414 65718 73466
rect 65898 73414 65900 73466
rect 65654 73412 65660 73414
rect 65716 73412 65740 73414
rect 65796 73412 65820 73414
rect 65876 73412 65900 73414
rect 65956 73412 65962 73414
rect 65654 73403 65962 73412
rect 68296 73234 68324 73646
rect 68284 73228 68336 73234
rect 68284 73170 68336 73176
rect 66314 72924 66622 72933
rect 66314 72922 66320 72924
rect 66376 72922 66400 72924
rect 66456 72922 66480 72924
rect 66536 72922 66560 72924
rect 66616 72922 66622 72924
rect 66376 72870 66378 72922
rect 66558 72870 66560 72922
rect 66314 72868 66320 72870
rect 66376 72868 66400 72870
rect 66456 72868 66480 72870
rect 66536 72868 66560 72870
rect 66616 72868 66622 72870
rect 66314 72859 66622 72868
rect 65654 72380 65962 72389
rect 65654 72378 65660 72380
rect 65716 72378 65740 72380
rect 65796 72378 65820 72380
rect 65876 72378 65900 72380
rect 65956 72378 65962 72380
rect 65716 72326 65718 72378
rect 65898 72326 65900 72378
rect 65654 72324 65660 72326
rect 65716 72324 65740 72326
rect 65796 72324 65820 72326
rect 65876 72324 65900 72326
rect 65956 72324 65962 72326
rect 65654 72315 65962 72324
rect 66314 71836 66622 71845
rect 66314 71834 66320 71836
rect 66376 71834 66400 71836
rect 66456 71834 66480 71836
rect 66536 71834 66560 71836
rect 66616 71834 66622 71836
rect 66376 71782 66378 71834
rect 66558 71782 66560 71834
rect 66314 71780 66320 71782
rect 66376 71780 66400 71782
rect 66456 71780 66480 71782
rect 66536 71780 66560 71782
rect 66616 71780 66622 71782
rect 66314 71771 66622 71780
rect 65654 71292 65962 71301
rect 65654 71290 65660 71292
rect 65716 71290 65740 71292
rect 65796 71290 65820 71292
rect 65876 71290 65900 71292
rect 65956 71290 65962 71292
rect 65716 71238 65718 71290
rect 65898 71238 65900 71290
rect 65654 71236 65660 71238
rect 65716 71236 65740 71238
rect 65796 71236 65820 71238
rect 65876 71236 65900 71238
rect 65956 71236 65962 71238
rect 65654 71227 65962 71236
rect 66314 70748 66622 70757
rect 66314 70746 66320 70748
rect 66376 70746 66400 70748
rect 66456 70746 66480 70748
rect 66536 70746 66560 70748
rect 66616 70746 66622 70748
rect 66376 70694 66378 70746
rect 66558 70694 66560 70746
rect 66314 70692 66320 70694
rect 66376 70692 66400 70694
rect 66456 70692 66480 70694
rect 66536 70692 66560 70694
rect 66616 70692 66622 70694
rect 66314 70683 66622 70692
rect 65654 70204 65962 70213
rect 65654 70202 65660 70204
rect 65716 70202 65740 70204
rect 65796 70202 65820 70204
rect 65876 70202 65900 70204
rect 65956 70202 65962 70204
rect 65716 70150 65718 70202
rect 65898 70150 65900 70202
rect 65654 70148 65660 70150
rect 65716 70148 65740 70150
rect 65796 70148 65820 70150
rect 65876 70148 65900 70150
rect 65956 70148 65962 70150
rect 65654 70139 65962 70148
rect 66720 69760 66772 69766
rect 66720 69702 66772 69708
rect 66314 69660 66622 69669
rect 66314 69658 66320 69660
rect 66376 69658 66400 69660
rect 66456 69658 66480 69660
rect 66536 69658 66560 69660
rect 66616 69658 66622 69660
rect 66376 69606 66378 69658
rect 66558 69606 66560 69658
rect 66314 69604 66320 69606
rect 66376 69604 66400 69606
rect 66456 69604 66480 69606
rect 66536 69604 66560 69606
rect 66616 69604 66622 69606
rect 66314 69595 66622 69604
rect 66732 69426 66760 69702
rect 67364 69556 67416 69562
rect 67364 69498 67416 69504
rect 67180 69488 67232 69494
rect 67376 69442 67404 69498
rect 67232 69436 67404 69442
rect 67180 69430 67404 69436
rect 66720 69420 66772 69426
rect 67192 69414 67404 69430
rect 66720 69362 66772 69368
rect 66444 69352 66496 69358
rect 66442 69320 66444 69329
rect 66496 69320 66498 69329
rect 66442 69255 66498 69264
rect 61476 69216 61528 69222
rect 61476 69158 61528 69164
rect 58624 69012 58676 69018
rect 58624 68954 58676 68960
rect 58714 68776 58770 68785
rect 58714 68711 58716 68720
rect 58768 68711 58770 68720
rect 58716 68682 58768 68688
rect 61488 68678 61516 69158
rect 65654 69116 65962 69125
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69051 65962 69060
rect 67376 69018 67404 69414
rect 67364 69012 67416 69018
rect 67364 68954 67416 68960
rect 68572 68814 68600 73714
rect 68940 73166 68968 76570
rect 69112 76356 69164 76362
rect 69112 76298 69164 76304
rect 69020 73772 69072 73778
rect 69020 73714 69072 73720
rect 68928 73160 68980 73166
rect 68928 73102 68980 73108
rect 68652 70984 68704 70990
rect 68652 70926 68704 70932
rect 68560 68808 68612 68814
rect 68560 68750 68612 68756
rect 66076 68740 66128 68746
rect 66076 68682 66128 68688
rect 46480 68672 46532 68678
rect 61476 68672 61528 68678
rect 46480 68614 46532 68620
rect 61474 68640 61476 68649
rect 61528 68640 61530 68649
rect 45098 65648 45154 65657
rect 45098 65583 45154 65592
rect 41142 64288 41198 64297
rect 41142 64223 41198 64232
rect 46492 64161 46520 68614
rect 61474 68575 61530 68584
rect 65654 68028 65962 68037
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67963 65962 67972
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 66088 64161 66116 68682
rect 66314 68572 66622 68581
rect 66314 68570 66320 68572
rect 66376 68570 66400 68572
rect 66456 68570 66480 68572
rect 66536 68570 66560 68572
rect 66616 68570 66622 68572
rect 66376 68518 66378 68570
rect 66558 68518 66560 68570
rect 66314 68516 66320 68518
rect 66376 68516 66400 68518
rect 66456 68516 66480 68518
rect 66536 68516 66560 68518
rect 66616 68516 66622 68518
rect 66314 68507 66622 68516
rect 66314 67484 66622 67493
rect 66314 67482 66320 67484
rect 66376 67482 66400 67484
rect 66456 67482 66480 67484
rect 66536 67482 66560 67484
rect 66616 67482 66622 67484
rect 66376 67430 66378 67482
rect 66558 67430 66560 67482
rect 66314 67428 66320 67430
rect 66376 67428 66400 67430
rect 66456 67428 66480 67430
rect 66536 67428 66560 67430
rect 66616 67428 66622 67430
rect 66314 67419 66622 67428
rect 66314 66396 66622 66405
rect 66314 66394 66320 66396
rect 66376 66394 66400 66396
rect 66456 66394 66480 66396
rect 66536 66394 66560 66396
rect 66616 66394 66622 66396
rect 66376 66342 66378 66394
rect 66558 66342 66560 66394
rect 66314 66340 66320 66342
rect 66376 66340 66400 66342
rect 66456 66340 66480 66342
rect 66536 66340 66560 66342
rect 66616 66340 66622 66342
rect 66314 66331 66622 66340
rect 68664 66230 68692 70926
rect 69032 69426 69060 73714
rect 69124 73302 69152 76298
rect 70124 76016 70176 76022
rect 70124 75958 70176 75964
rect 70136 73914 70164 75958
rect 70124 73908 70176 73914
rect 70124 73850 70176 73856
rect 72424 73704 72476 73710
rect 72424 73646 72476 73652
rect 70584 73568 70636 73574
rect 70584 73510 70636 73516
rect 70596 73370 70624 73510
rect 70584 73364 70636 73370
rect 70584 73306 70636 73312
rect 69112 73296 69164 73302
rect 69112 73238 69164 73244
rect 69124 73030 69152 73238
rect 72436 73234 72464 73646
rect 73816 73642 73844 79290
rect 89904 77988 89956 77994
rect 89904 77930 89956 77936
rect 87236 77920 87288 77926
rect 87236 77862 87288 77868
rect 87248 77654 87276 77862
rect 87236 77648 87288 77654
rect 87236 77590 87288 77596
rect 89628 77648 89680 77654
rect 89628 77590 89680 77596
rect 89720 77648 89772 77654
rect 89720 77590 89772 77596
rect 89812 77648 89864 77654
rect 89812 77590 89864 77596
rect 86408 77580 86460 77586
rect 86408 77522 86460 77528
rect 82820 77376 82872 77382
rect 82740 77336 82820 77364
rect 82740 76498 82768 77336
rect 82820 77318 82872 77324
rect 84016 77376 84068 77382
rect 84016 77318 84068 77324
rect 85856 77376 85908 77382
rect 85856 77318 85908 77324
rect 82544 76492 82596 76498
rect 82544 76434 82596 76440
rect 82728 76492 82780 76498
rect 82728 76434 82780 76440
rect 82556 76294 82584 76434
rect 74540 76288 74592 76294
rect 74540 76230 74592 76236
rect 82544 76288 82596 76294
rect 82544 76230 82596 76236
rect 83096 76288 83148 76294
rect 83096 76230 83148 76236
rect 83464 76288 83516 76294
rect 83464 76230 83516 76236
rect 83648 76288 83700 76294
rect 83648 76230 83700 76236
rect 74172 74248 74224 74254
rect 74172 74190 74224 74196
rect 74184 73778 74212 74190
rect 74552 73914 74580 76230
rect 82556 74458 82584 76230
rect 75092 74452 75144 74458
rect 75092 74394 75144 74400
rect 82544 74452 82596 74458
rect 82544 74394 82596 74400
rect 75104 73914 75132 74394
rect 78772 74248 78824 74254
rect 78772 74190 78824 74196
rect 74540 73908 74592 73914
rect 74540 73850 74592 73856
rect 75092 73908 75144 73914
rect 75092 73850 75144 73856
rect 74724 73840 74776 73846
rect 74908 73840 74960 73846
rect 74776 73788 74908 73794
rect 74724 73782 74960 73788
rect 74172 73772 74224 73778
rect 74172 73714 74224 73720
rect 74540 73772 74592 73778
rect 74736 73766 74948 73782
rect 74540 73714 74592 73720
rect 73160 73636 73212 73642
rect 73160 73578 73212 73584
rect 73804 73636 73856 73642
rect 73804 73578 73856 73584
rect 72424 73228 72476 73234
rect 72424 73170 72476 73176
rect 72884 73228 72936 73234
rect 72884 73170 72936 73176
rect 70216 73092 70268 73098
rect 70216 73034 70268 73040
rect 70400 73092 70452 73098
rect 70400 73034 70452 73040
rect 69112 73024 69164 73030
rect 69112 72966 69164 72972
rect 69124 72826 69152 72966
rect 69112 72820 69164 72826
rect 69112 72762 69164 72768
rect 69124 69562 69152 72762
rect 69112 69556 69164 69562
rect 69112 69498 69164 69504
rect 69020 69420 69072 69426
rect 69020 69362 69072 69368
rect 70228 67658 70256 73034
rect 70412 68950 70440 73034
rect 72896 71058 72924 73170
rect 73068 73024 73120 73030
rect 73068 72966 73120 72972
rect 73080 72826 73108 72966
rect 73068 72820 73120 72826
rect 73068 72762 73120 72768
rect 72884 71052 72936 71058
rect 72884 70994 72936 71000
rect 72700 70848 72752 70854
rect 72700 70790 72752 70796
rect 72712 69873 72740 70790
rect 72896 70106 72924 70994
rect 72884 70100 72936 70106
rect 72884 70042 72936 70048
rect 72698 69864 72754 69873
rect 72698 69799 72754 69808
rect 72424 69760 72476 69766
rect 72424 69702 72476 69708
rect 70400 68944 70452 68950
rect 70400 68886 70452 68892
rect 70216 67652 70268 67658
rect 70216 67594 70268 67600
rect 68652 66224 68704 66230
rect 68650 66192 68652 66201
rect 68704 66192 68706 66201
rect 68650 66127 68706 66136
rect 39946 64152 40002 64161
rect 39946 64087 40002 64096
rect 46478 64152 46534 64161
rect 46478 64087 46534 64096
rect 66074 64152 66130 64161
rect 66074 64087 66130 64096
rect 72436 64025 72464 69702
rect 73172 66230 73200 73578
rect 74552 69222 74580 73714
rect 78588 73704 78640 73710
rect 78588 73646 78640 73652
rect 78600 73370 78628 73646
rect 78588 73364 78640 73370
rect 78588 73306 78640 73312
rect 78784 73302 78812 74190
rect 78772 73296 78824 73302
rect 78772 73238 78824 73244
rect 81992 73092 82044 73098
rect 81992 73034 82044 73040
rect 82004 72282 82032 73034
rect 81992 72276 82044 72282
rect 81992 72218 82044 72224
rect 79508 70984 79560 70990
rect 79508 70926 79560 70932
rect 81164 70984 81216 70990
rect 81164 70926 81216 70932
rect 79520 69970 79548 70926
rect 81176 70106 81204 70926
rect 81164 70100 81216 70106
rect 81164 70042 81216 70048
rect 83108 69970 83136 76230
rect 83476 75954 83504 76230
rect 83660 76090 83688 76230
rect 83648 76084 83700 76090
rect 83648 76026 83700 76032
rect 83464 75948 83516 75954
rect 83464 75890 83516 75896
rect 83464 71936 83516 71942
rect 83464 71878 83516 71884
rect 83476 70990 83504 71878
rect 84028 71194 84056 77318
rect 85868 76498 85896 77318
rect 86420 77178 86448 77522
rect 89640 77450 89668 77590
rect 89628 77444 89680 77450
rect 89628 77386 89680 77392
rect 86776 77376 86828 77382
rect 86776 77318 86828 77324
rect 86408 77172 86460 77178
rect 86408 77114 86460 77120
rect 85856 76492 85908 76498
rect 85856 76434 85908 76440
rect 84844 76356 84896 76362
rect 84844 76298 84896 76304
rect 84856 76090 84884 76298
rect 84844 76084 84896 76090
rect 84844 76026 84896 76032
rect 84856 75993 84884 76026
rect 84842 75984 84898 75993
rect 84842 75919 84898 75928
rect 85672 74928 85724 74934
rect 85672 74870 85724 74876
rect 85684 74458 85712 74870
rect 85948 74656 86000 74662
rect 85948 74598 86000 74604
rect 85960 74458 85988 74598
rect 85672 74452 85724 74458
rect 85672 74394 85724 74400
rect 85948 74452 86000 74458
rect 85948 74394 86000 74400
rect 84292 74384 84344 74390
rect 84292 74326 84344 74332
rect 84304 73778 84332 74326
rect 85960 74254 85988 74394
rect 85120 74248 85172 74254
rect 85120 74190 85172 74196
rect 85948 74248 86000 74254
rect 85948 74190 86000 74196
rect 85132 73778 85160 74190
rect 84292 73772 84344 73778
rect 84292 73714 84344 73720
rect 85120 73772 85172 73778
rect 85120 73714 85172 73720
rect 85132 72214 85160 73714
rect 85580 73704 85632 73710
rect 85580 73646 85632 73652
rect 85592 72826 85620 73646
rect 86040 73568 86092 73574
rect 86040 73510 86092 73516
rect 85580 72820 85632 72826
rect 85580 72762 85632 72768
rect 85488 72752 85540 72758
rect 85488 72694 85540 72700
rect 85500 72282 85528 72694
rect 86052 72570 86080 73510
rect 86684 72820 86736 72826
rect 86684 72762 86736 72768
rect 86696 72622 86724 72762
rect 86224 72616 86276 72622
rect 86052 72564 86224 72570
rect 86052 72558 86276 72564
rect 86684 72616 86736 72622
rect 86684 72558 86736 72564
rect 86052 72542 86264 72558
rect 86052 72486 86080 72542
rect 86040 72480 86092 72486
rect 86040 72422 86092 72428
rect 85488 72276 85540 72282
rect 85488 72218 85540 72224
rect 85120 72208 85172 72214
rect 85120 72150 85172 72156
rect 85212 72140 85264 72146
rect 85212 72082 85264 72088
rect 84844 71392 84896 71398
rect 84844 71334 84896 71340
rect 84016 71188 84068 71194
rect 84016 71130 84068 71136
rect 83464 70984 83516 70990
rect 83464 70926 83516 70932
rect 84856 70582 84884 71334
rect 85224 71194 85252 72082
rect 85396 72072 85448 72078
rect 85396 72014 85448 72020
rect 85212 71188 85264 71194
rect 85212 71130 85264 71136
rect 85408 71126 85436 72014
rect 85396 71120 85448 71126
rect 85396 71062 85448 71068
rect 85408 70990 85436 71062
rect 86052 71058 86080 72422
rect 86316 71188 86368 71194
rect 86316 71130 86368 71136
rect 86040 71052 86092 71058
rect 86040 70994 86092 71000
rect 85396 70984 85448 70990
rect 85396 70926 85448 70932
rect 84844 70576 84896 70582
rect 84844 70518 84896 70524
rect 85408 69970 85436 70926
rect 79508 69964 79560 69970
rect 79508 69906 79560 69912
rect 83096 69964 83148 69970
rect 83096 69906 83148 69912
rect 85396 69964 85448 69970
rect 85396 69906 85448 69912
rect 79324 69896 79376 69902
rect 79322 69864 79324 69873
rect 79376 69864 79378 69873
rect 77852 69828 77904 69834
rect 79322 69799 79378 69808
rect 77852 69770 77904 69776
rect 74540 69216 74592 69222
rect 74540 69158 74592 69164
rect 74356 67652 74408 67658
rect 74356 67594 74408 67600
rect 74368 66230 74396 67594
rect 73160 66224 73212 66230
rect 73160 66166 73212 66172
rect 74356 66224 74408 66230
rect 74356 66166 74408 66172
rect 72422 64016 72478 64025
rect 72422 63951 72478 63960
rect 77864 63889 77892 69770
rect 79336 69766 79364 69799
rect 79324 69760 79376 69766
rect 79324 69702 79376 69708
rect 79336 69562 79364 69702
rect 79324 69556 79376 69562
rect 79324 69498 79376 69504
rect 85408 66638 85436 69906
rect 86052 67726 86080 70994
rect 86328 69426 86356 71130
rect 86788 69902 86816 77318
rect 89732 77178 89760 77590
rect 89824 77382 89852 77590
rect 89916 77586 89944 77930
rect 89904 77580 89956 77586
rect 89904 77522 89956 77528
rect 89812 77376 89864 77382
rect 89812 77318 89864 77324
rect 90088 77376 90140 77382
rect 90088 77318 90140 77324
rect 89720 77172 89772 77178
rect 89720 77114 89772 77120
rect 88432 77036 88484 77042
rect 88432 76978 88484 76984
rect 86868 76424 86920 76430
rect 86868 76366 86920 76372
rect 86880 75342 86908 76366
rect 88248 75812 88300 75818
rect 88248 75754 88300 75760
rect 88064 75744 88116 75750
rect 88116 75704 88196 75732
rect 88064 75686 88116 75692
rect 86868 75336 86920 75342
rect 86868 75278 86920 75284
rect 86880 75002 86908 75278
rect 88168 75274 88196 75704
rect 88260 75478 88288 75754
rect 88248 75472 88300 75478
rect 88248 75414 88300 75420
rect 88156 75268 88208 75274
rect 88156 75210 88208 75216
rect 87788 75200 87840 75206
rect 87788 75142 87840 75148
rect 86868 74996 86920 75002
rect 86868 74938 86920 74944
rect 87800 74934 87828 75142
rect 88168 75002 88196 75210
rect 88156 74996 88208 75002
rect 88156 74938 88208 74944
rect 87788 74928 87840 74934
rect 87788 74870 87840 74876
rect 88168 74798 88196 74938
rect 88340 74928 88392 74934
rect 88340 74870 88392 74876
rect 88156 74792 88208 74798
rect 88156 74734 88208 74740
rect 87144 74452 87196 74458
rect 87144 74394 87196 74400
rect 88156 74452 88208 74458
rect 88156 74394 88208 74400
rect 87156 74254 87184 74394
rect 87144 74248 87196 74254
rect 87144 74190 87196 74196
rect 88168 73370 88196 74394
rect 88352 74322 88380 74870
rect 88340 74316 88392 74322
rect 88340 74258 88392 74264
rect 88156 73364 88208 73370
rect 88156 73306 88208 73312
rect 88168 72282 88196 73306
rect 88156 72276 88208 72282
rect 88156 72218 88208 72224
rect 87788 70916 87840 70922
rect 87788 70858 87840 70864
rect 87800 70650 87828 70858
rect 87788 70644 87840 70650
rect 87788 70586 87840 70592
rect 88156 70644 88208 70650
rect 88156 70586 88208 70592
rect 86776 69896 86828 69902
rect 86776 69838 86828 69844
rect 86316 69420 86368 69426
rect 86316 69362 86368 69368
rect 86868 68808 86920 68814
rect 86868 68750 86920 68756
rect 86776 68672 86828 68678
rect 86776 68614 86828 68620
rect 86788 67794 86816 68614
rect 86776 67788 86828 67794
rect 86776 67730 86828 67736
rect 86040 67720 86092 67726
rect 86040 67662 86092 67668
rect 86880 67386 86908 68750
rect 87144 67720 87196 67726
rect 87144 67662 87196 67668
rect 86868 67380 86920 67386
rect 86868 67322 86920 67328
rect 86776 67040 86828 67046
rect 86776 66982 86828 66988
rect 86788 66638 86816 66982
rect 85396 66632 85448 66638
rect 85396 66574 85448 66580
rect 86776 66632 86828 66638
rect 86776 66574 86828 66580
rect 86868 66564 86920 66570
rect 86868 66506 86920 66512
rect 86880 66162 86908 66506
rect 87156 66502 87184 67662
rect 87420 67584 87472 67590
rect 87420 67526 87472 67532
rect 87432 67386 87460 67526
rect 87420 67380 87472 67386
rect 87420 67322 87472 67328
rect 87144 66496 87196 66502
rect 87144 66438 87196 66444
rect 87156 66298 87184 66438
rect 87144 66292 87196 66298
rect 87144 66234 87196 66240
rect 86868 66156 86920 66162
rect 86868 66098 86920 66104
rect 88168 66042 88196 70586
rect 88444 70394 88472 76978
rect 89260 76968 89312 76974
rect 89260 76910 89312 76916
rect 88708 74996 88760 75002
rect 88708 74938 88760 74944
rect 88720 74730 88748 74938
rect 88708 74724 88760 74730
rect 88708 74666 88760 74672
rect 88984 74656 89036 74662
rect 88984 74598 89036 74604
rect 88800 74112 88852 74118
rect 88800 74054 88852 74060
rect 88812 73930 88840 74054
rect 88720 73914 88840 73930
rect 88708 73908 88840 73914
rect 88760 73902 88840 73908
rect 88708 73850 88760 73856
rect 88996 72593 89024 74598
rect 89076 73704 89128 73710
rect 89076 73646 89128 73652
rect 88982 72584 89038 72593
rect 88982 72519 89038 72528
rect 89088 72486 89116 73646
rect 89076 72480 89128 72486
rect 89076 72422 89128 72428
rect 89168 71392 89220 71398
rect 89168 71334 89220 71340
rect 89180 71058 89208 71334
rect 89168 71052 89220 71058
rect 89168 70994 89220 71000
rect 89272 70854 89300 76910
rect 89732 75818 89760 77114
rect 89720 75812 89772 75818
rect 89720 75754 89772 75760
rect 89628 75268 89680 75274
rect 89628 75210 89680 75216
rect 89640 75002 89668 75210
rect 89732 75002 89760 75754
rect 89628 74996 89680 75002
rect 89628 74938 89680 74944
rect 89720 74996 89772 75002
rect 89720 74938 89772 74944
rect 89824 74780 89852 77318
rect 90100 75750 90128 77318
rect 90284 77042 90312 79358
rect 91928 78192 91980 78198
rect 91928 78134 91980 78140
rect 91466 77752 91522 77761
rect 91192 77716 91244 77722
rect 91466 77687 91522 77696
rect 91192 77658 91244 77664
rect 90548 77648 90600 77654
rect 90548 77590 90600 77596
rect 90364 77172 90416 77178
rect 90364 77114 90416 77120
rect 90376 77042 90404 77114
rect 90560 77042 90588 77590
rect 90272 77036 90324 77042
rect 90272 76978 90324 76984
rect 90364 77036 90416 77042
rect 90364 76978 90416 76984
rect 90548 77036 90600 77042
rect 90548 76978 90600 76984
rect 90456 76832 90508 76838
rect 90456 76774 90508 76780
rect 90468 76090 90496 76774
rect 90456 76084 90508 76090
rect 90456 76026 90508 76032
rect 90272 76016 90324 76022
rect 90272 75958 90324 75964
rect 89904 75744 89956 75750
rect 89904 75686 89956 75692
rect 90088 75744 90140 75750
rect 90088 75686 90140 75692
rect 89916 75206 89944 75686
rect 90284 75546 90312 75958
rect 91204 75954 91232 77658
rect 91480 77450 91508 77687
rect 91940 77654 91968 78134
rect 91928 77648 91980 77654
rect 91928 77590 91980 77596
rect 91558 77480 91614 77489
rect 91468 77444 91520 77450
rect 91558 77415 91614 77424
rect 91468 77386 91520 77392
rect 91572 77382 91600 77415
rect 91560 77376 91612 77382
rect 91560 77318 91612 77324
rect 91192 75948 91244 75954
rect 91192 75890 91244 75896
rect 90272 75540 90324 75546
rect 90272 75482 90324 75488
rect 91008 75540 91060 75546
rect 91008 75482 91060 75488
rect 90732 75268 90784 75274
rect 90732 75210 90784 75216
rect 89904 75200 89956 75206
rect 89904 75142 89956 75148
rect 90744 74798 90772 75210
rect 89904 74792 89956 74798
rect 89824 74752 89904 74780
rect 89904 74734 89956 74740
rect 90732 74792 90784 74798
rect 90732 74734 90784 74740
rect 91020 73846 91048 75482
rect 91204 74458 91232 75890
rect 91468 75268 91520 75274
rect 91468 75210 91520 75216
rect 91376 75200 91428 75206
rect 91376 75142 91428 75148
rect 91284 74656 91336 74662
rect 91284 74598 91336 74604
rect 91192 74452 91244 74458
rect 91192 74394 91244 74400
rect 91204 74254 91232 74394
rect 91192 74248 91244 74254
rect 91192 74190 91244 74196
rect 89536 73840 89588 73846
rect 89536 73782 89588 73788
rect 91008 73840 91060 73846
rect 91008 73782 91060 73788
rect 89548 73166 89576 73782
rect 89628 73568 89680 73574
rect 89628 73510 89680 73516
rect 89536 73160 89588 73166
rect 89536 73102 89588 73108
rect 89640 71670 89668 73510
rect 89720 72276 89772 72282
rect 89720 72218 89772 72224
rect 89628 71664 89680 71670
rect 89628 71606 89680 71612
rect 89260 70848 89312 70854
rect 89260 70790 89312 70796
rect 88800 70508 88852 70514
rect 88800 70450 88852 70456
rect 88352 70366 88472 70394
rect 88352 70038 88380 70366
rect 88340 70032 88392 70038
rect 88340 69974 88392 69980
rect 88812 69562 88840 70450
rect 89732 70106 89760 72218
rect 90088 72004 90140 72010
rect 90088 71946 90140 71952
rect 90100 71670 90128 71946
rect 90088 71664 90140 71670
rect 90088 71606 90140 71612
rect 90364 70576 90416 70582
rect 90364 70518 90416 70524
rect 89720 70100 89772 70106
rect 89720 70042 89772 70048
rect 88800 69556 88852 69562
rect 88800 69498 88852 69504
rect 89732 69426 89760 70042
rect 90376 70038 90404 70518
rect 91020 70446 91048 73782
rect 91296 73778 91324 74598
rect 91388 74118 91416 75142
rect 91480 74866 91508 75210
rect 91468 74860 91520 74866
rect 91468 74802 91520 74808
rect 91468 74656 91520 74662
rect 91468 74598 91520 74604
rect 91376 74112 91428 74118
rect 91376 74054 91428 74060
rect 91388 73914 91416 74054
rect 91376 73908 91428 73914
rect 91376 73850 91428 73856
rect 91284 73772 91336 73778
rect 91284 73714 91336 73720
rect 91388 73574 91416 73850
rect 91480 73642 91508 74598
rect 91468 73636 91520 73642
rect 91468 73578 91520 73584
rect 91376 73568 91428 73574
rect 91376 73510 91428 73516
rect 91008 70440 91060 70446
rect 91572 70394 91600 77318
rect 91940 77042 91968 77590
rect 92020 77444 92072 77450
rect 92020 77386 92072 77392
rect 91928 77036 91980 77042
rect 91928 76978 91980 76984
rect 91836 74996 91888 75002
rect 91836 74938 91888 74944
rect 91848 74866 91876 74938
rect 91836 74860 91888 74866
rect 91836 74802 91888 74808
rect 91836 73568 91888 73574
rect 91836 73510 91888 73516
rect 91008 70382 91060 70388
rect 90640 70100 90692 70106
rect 90640 70042 90692 70048
rect 90364 70032 90416 70038
rect 90364 69974 90416 69980
rect 90376 69902 90404 69974
rect 90652 69970 90680 70042
rect 90640 69964 90692 69970
rect 90640 69906 90692 69912
rect 90364 69896 90416 69902
rect 90364 69838 90416 69844
rect 89720 69420 89772 69426
rect 89720 69362 89772 69368
rect 89076 69352 89128 69358
rect 89076 69294 89128 69300
rect 89088 67930 89116 69294
rect 89732 69018 89760 69362
rect 89720 69012 89772 69018
rect 89720 68954 89772 68960
rect 89260 68672 89312 68678
rect 89260 68614 89312 68620
rect 89076 67924 89128 67930
rect 89076 67866 89128 67872
rect 89272 67726 89300 68614
rect 91020 68406 91048 70382
rect 91480 70366 91600 70394
rect 91008 68400 91060 68406
rect 91008 68342 91060 68348
rect 89444 67924 89496 67930
rect 89444 67866 89496 67872
rect 90824 67924 90876 67930
rect 90824 67866 90876 67872
rect 89260 67720 89312 67726
rect 89260 67662 89312 67668
rect 89076 67584 89128 67590
rect 89076 67526 89128 67532
rect 88248 66496 88300 66502
rect 88248 66438 88300 66444
rect 88260 66162 88288 66438
rect 88616 66292 88668 66298
rect 88616 66234 88668 66240
rect 88248 66156 88300 66162
rect 88248 66098 88300 66104
rect 88628 66094 88656 66234
rect 89088 66230 89116 67526
rect 89272 66638 89300 67662
rect 89352 67584 89404 67590
rect 89352 67526 89404 67532
rect 89364 67386 89392 67526
rect 89352 67380 89404 67386
rect 89352 67322 89404 67328
rect 89352 67244 89404 67250
rect 89352 67186 89404 67192
rect 89364 66638 89392 67186
rect 89456 66842 89484 67866
rect 89720 67652 89772 67658
rect 89720 67594 89772 67600
rect 89996 67652 90048 67658
rect 89996 67594 90048 67600
rect 89444 66836 89496 66842
rect 89444 66778 89496 66784
rect 89260 66632 89312 66638
rect 89260 66574 89312 66580
rect 89352 66632 89404 66638
rect 89352 66574 89404 66580
rect 89076 66224 89128 66230
rect 89076 66166 89128 66172
rect 89272 66162 89300 66574
rect 89364 66298 89392 66574
rect 89352 66292 89404 66298
rect 89352 66234 89404 66240
rect 89732 66230 89760 67594
rect 89904 67312 89956 67318
rect 89904 67254 89956 67260
rect 89812 67040 89864 67046
rect 89812 66982 89864 66988
rect 89824 66842 89852 66982
rect 89812 66836 89864 66842
rect 89812 66778 89864 66784
rect 89916 66638 89944 67254
rect 89904 66632 89956 66638
rect 89904 66574 89956 66580
rect 90008 66570 90036 67594
rect 90180 67380 90232 67386
rect 90180 67322 90232 67328
rect 89996 66564 90048 66570
rect 89996 66506 90048 66512
rect 89904 66496 89956 66502
rect 89904 66438 89956 66444
rect 89916 66298 89944 66438
rect 89904 66292 89956 66298
rect 89904 66234 89956 66240
rect 89720 66224 89772 66230
rect 89720 66166 89772 66172
rect 90192 66162 90220 67322
rect 90640 66836 90692 66842
rect 90640 66778 90692 66784
rect 90652 66230 90680 66778
rect 90640 66224 90692 66230
rect 90640 66166 90692 66172
rect 89260 66156 89312 66162
rect 89260 66098 89312 66104
rect 90180 66156 90232 66162
rect 90180 66098 90232 66104
rect 90732 66156 90784 66162
rect 90732 66098 90784 66104
rect 88616 66088 88668 66094
rect 88168 66014 88288 66042
rect 88616 66030 88668 66036
rect 89272 66026 89300 66098
rect 88260 65958 88288 66014
rect 89260 66020 89312 66026
rect 89260 65962 89312 65968
rect 90744 65958 90772 66098
rect 90836 66094 90864 67866
rect 91020 67658 91048 68342
rect 91008 67652 91060 67658
rect 91008 67594 91060 67600
rect 91480 67318 91508 70366
rect 91560 69488 91612 69494
rect 91560 69430 91612 69436
rect 91572 68474 91600 69430
rect 91848 69426 91876 73510
rect 91836 69420 91888 69426
rect 91836 69362 91888 69368
rect 91744 69216 91796 69222
rect 91744 69158 91796 69164
rect 91756 68882 91784 69158
rect 91744 68876 91796 68882
rect 91744 68818 91796 68824
rect 91560 68468 91612 68474
rect 91560 68410 91612 68416
rect 91928 68400 91980 68406
rect 91928 68342 91980 68348
rect 91940 67930 91968 68342
rect 91928 67924 91980 67930
rect 91928 67866 91980 67872
rect 91468 67312 91520 67318
rect 91468 67254 91520 67260
rect 91192 67244 91244 67250
rect 91192 67186 91244 67192
rect 91204 66842 91232 67186
rect 91192 66836 91244 66842
rect 91192 66778 91244 66784
rect 91480 66706 91508 67254
rect 92032 66774 92060 77386
rect 92124 77042 92152 79426
rect 96804 79212 96856 79218
rect 96804 79154 96856 79160
rect 95884 78668 95936 78674
rect 95884 78610 95936 78616
rect 92388 78056 92440 78062
rect 92388 77998 92440 78004
rect 92202 77616 92258 77625
rect 92202 77551 92258 77560
rect 92216 77382 92244 77551
rect 92204 77376 92256 77382
rect 92204 77318 92256 77324
rect 92112 77036 92164 77042
rect 92112 76978 92164 76984
rect 92216 67114 92244 77318
rect 92400 75274 92428 77998
rect 94872 77716 94924 77722
rect 94872 77658 94924 77664
rect 94884 77518 94912 77658
rect 92480 77512 92532 77518
rect 92480 77454 92532 77460
rect 93952 77512 94004 77518
rect 93952 77454 94004 77460
rect 94872 77512 94924 77518
rect 94872 77454 94924 77460
rect 92492 76634 92520 77454
rect 93964 77382 93992 77454
rect 95240 77444 95292 77450
rect 95240 77386 95292 77392
rect 92572 77376 92624 77382
rect 92572 77318 92624 77324
rect 93952 77376 94004 77382
rect 93952 77318 94004 77324
rect 92584 76838 92612 77318
rect 93964 77042 93992 77318
rect 95252 77178 95280 77386
rect 95240 77172 95292 77178
rect 95240 77114 95292 77120
rect 93952 77036 94004 77042
rect 93952 76978 94004 76984
rect 92572 76832 92624 76838
rect 92572 76774 92624 76780
rect 92480 76628 92532 76634
rect 92480 76570 92532 76576
rect 92584 76294 92612 76774
rect 93492 76356 93544 76362
rect 93492 76298 93544 76304
rect 92572 76288 92624 76294
rect 92572 76230 92624 76236
rect 92584 75750 92612 76230
rect 93504 76090 93532 76298
rect 93492 76084 93544 76090
rect 93492 76026 93544 76032
rect 93400 76016 93452 76022
rect 93400 75958 93452 75964
rect 92572 75744 92624 75750
rect 92572 75686 92624 75692
rect 92388 75268 92440 75274
rect 92388 75210 92440 75216
rect 92400 74866 92428 75210
rect 92584 75206 92612 75686
rect 93412 75410 93440 75958
rect 93400 75404 93452 75410
rect 93400 75346 93452 75352
rect 93032 75268 93084 75274
rect 93032 75210 93084 75216
rect 92572 75200 92624 75206
rect 92572 75142 92624 75148
rect 92388 74860 92440 74866
rect 92388 74802 92440 74808
rect 92400 74610 92428 74802
rect 92400 74582 92520 74610
rect 92492 71738 92520 74582
rect 93044 74458 93072 75210
rect 93308 74996 93360 75002
rect 93308 74938 93360 74944
rect 93032 74452 93084 74458
rect 93032 74394 93084 74400
rect 93320 73914 93348 74938
rect 93964 74934 93992 76978
rect 94044 76832 94096 76838
rect 94044 76774 94096 76780
rect 94056 76022 94084 76774
rect 95424 76560 95476 76566
rect 95424 76502 95476 76508
rect 94044 76016 94096 76022
rect 94044 75958 94096 75964
rect 95436 75886 95464 76502
rect 95424 75880 95476 75886
rect 95424 75822 95476 75828
rect 93952 74928 94004 74934
rect 93952 74870 94004 74876
rect 94044 74860 94096 74866
rect 94044 74802 94096 74808
rect 93308 73908 93360 73914
rect 93308 73850 93360 73856
rect 93320 73778 93348 73850
rect 93308 73772 93360 73778
rect 93308 73714 93360 73720
rect 93860 73772 93912 73778
rect 93860 73714 93912 73720
rect 93320 73370 93348 73714
rect 93584 73568 93636 73574
rect 93584 73510 93636 73516
rect 93308 73364 93360 73370
rect 93308 73306 93360 73312
rect 92480 71732 92532 71738
rect 92480 71674 92532 71680
rect 92492 71126 92520 71674
rect 93320 71194 93348 73306
rect 93596 72078 93624 73510
rect 93872 73234 93900 73714
rect 93952 73568 94004 73574
rect 93952 73510 94004 73516
rect 93860 73228 93912 73234
rect 93860 73170 93912 73176
rect 93584 72072 93636 72078
rect 93584 72014 93636 72020
rect 93768 72004 93820 72010
rect 93768 71946 93820 71952
rect 93308 71188 93360 71194
rect 93308 71130 93360 71136
rect 92480 71120 92532 71126
rect 92480 71062 92532 71068
rect 93320 70990 93348 71130
rect 93308 70984 93360 70990
rect 93308 70926 93360 70932
rect 93400 70984 93452 70990
rect 93400 70926 93452 70932
rect 92940 70848 92992 70854
rect 92940 70790 92992 70796
rect 93032 70848 93084 70854
rect 93032 70790 93084 70796
rect 92480 69828 92532 69834
rect 92480 69770 92532 69776
rect 92296 69488 92348 69494
rect 92296 69430 92348 69436
rect 92308 68406 92336 69430
rect 92492 69426 92520 69770
rect 92952 69562 92980 70790
rect 92940 69556 92992 69562
rect 92940 69498 92992 69504
rect 93044 69426 93072 70790
rect 93216 70644 93268 70650
rect 93320 70632 93348 70926
rect 93268 70604 93348 70632
rect 93216 70586 93268 70592
rect 93412 70564 93440 70926
rect 93320 70536 93440 70564
rect 93320 70310 93348 70536
rect 93308 70304 93360 70310
rect 93308 70246 93360 70252
rect 92480 69420 92532 69426
rect 92480 69362 92532 69368
rect 93032 69420 93084 69426
rect 93032 69362 93084 69368
rect 92756 69216 92808 69222
rect 92756 69158 92808 69164
rect 92296 68400 92348 68406
rect 92296 68342 92348 68348
rect 92572 67312 92624 67318
rect 92572 67254 92624 67260
rect 92204 67108 92256 67114
rect 92204 67050 92256 67056
rect 92480 66836 92532 66842
rect 92400 66796 92480 66824
rect 92020 66768 92072 66774
rect 92020 66710 92072 66716
rect 91468 66700 91520 66706
rect 91468 66642 91520 66648
rect 92296 66564 92348 66570
rect 92296 66506 92348 66512
rect 92308 66298 92336 66506
rect 92296 66292 92348 66298
rect 92296 66234 92348 66240
rect 92400 66094 92428 66796
rect 92480 66778 92532 66784
rect 92584 66502 92612 67254
rect 92768 67250 92796 69158
rect 92940 68468 92992 68474
rect 92940 68410 92992 68416
rect 92952 67386 92980 68410
rect 92940 67380 92992 67386
rect 92940 67322 92992 67328
rect 93044 67318 93072 69362
rect 93320 69018 93348 70246
rect 93780 69834 93808 71946
rect 93872 71942 93900 73170
rect 93964 72214 93992 73510
rect 93952 72208 94004 72214
rect 93952 72150 94004 72156
rect 93860 71936 93912 71942
rect 93860 71878 93912 71884
rect 93860 71052 93912 71058
rect 93860 70994 93912 71000
rect 93872 70854 93900 70994
rect 94056 70922 94084 74802
rect 94412 74656 94464 74662
rect 94412 74598 94464 74604
rect 94424 73778 94452 74598
rect 94412 73772 94464 73778
rect 94412 73714 94464 73720
rect 94504 72752 94556 72758
rect 94504 72694 94556 72700
rect 94516 72282 94544 72694
rect 94504 72276 94556 72282
rect 94504 72218 94556 72224
rect 94320 72072 94372 72078
rect 94320 72014 94372 72020
rect 94332 71466 94360 72014
rect 95056 71936 95108 71942
rect 95056 71878 95108 71884
rect 94320 71460 94372 71466
rect 94320 71402 94372 71408
rect 94044 70916 94096 70922
rect 94044 70858 94096 70864
rect 93860 70848 93912 70854
rect 93860 70790 93912 70796
rect 94332 69902 94360 71402
rect 94872 71052 94924 71058
rect 94872 70994 94924 71000
rect 94884 69902 94912 70994
rect 94320 69896 94372 69902
rect 94320 69838 94372 69844
rect 94872 69896 94924 69902
rect 94872 69838 94924 69844
rect 93768 69828 93820 69834
rect 93768 69770 93820 69776
rect 94780 69760 94832 69766
rect 94780 69702 94832 69708
rect 93308 69012 93360 69018
rect 93308 68954 93360 68960
rect 94504 68672 94556 68678
rect 94504 68614 94556 68620
rect 93400 68128 93452 68134
rect 93400 68070 93452 68076
rect 93412 67386 93440 68070
rect 94412 67856 94464 67862
rect 94412 67798 94464 67804
rect 93400 67380 93452 67386
rect 93400 67322 93452 67328
rect 93032 67312 93084 67318
rect 93032 67254 93084 67260
rect 92756 67244 92808 67250
rect 92756 67186 92808 67192
rect 92768 66570 92796 67186
rect 92756 66564 92808 66570
rect 92756 66506 92808 66512
rect 92572 66496 92624 66502
rect 92572 66438 92624 66444
rect 92584 66162 92612 66438
rect 92572 66156 92624 66162
rect 92572 66098 92624 66104
rect 94136 66156 94188 66162
rect 94136 66098 94188 66104
rect 90824 66088 90876 66094
rect 90824 66030 90876 66036
rect 92388 66088 92440 66094
rect 92388 66030 92440 66036
rect 88248 65952 88300 65958
rect 88246 65920 88248 65929
rect 90732 65952 90784 65958
rect 88300 65920 88302 65929
rect 90732 65894 90784 65900
rect 88246 65855 88302 65864
rect 94148 65754 94176 66098
rect 94424 65958 94452 67798
rect 94516 67182 94544 68614
rect 94792 68406 94820 69702
rect 94780 68400 94832 68406
rect 94780 68342 94832 68348
rect 94504 67176 94556 67182
rect 94504 67118 94556 67124
rect 94780 67108 94832 67114
rect 94780 67050 94832 67056
rect 94792 66570 94820 67050
rect 94780 66564 94832 66570
rect 94780 66506 94832 66512
rect 94792 66162 94820 66506
rect 94780 66156 94832 66162
rect 94780 66098 94832 66104
rect 94412 65952 94464 65958
rect 94412 65894 94464 65900
rect 94136 65748 94188 65754
rect 94136 65690 94188 65696
rect 94884 65686 94912 69838
rect 94964 69352 95016 69358
rect 94964 69294 95016 69300
rect 94976 68814 95004 69294
rect 94964 68808 95016 68814
rect 94964 68750 95016 68756
rect 95068 68270 95096 71878
rect 95700 71392 95752 71398
rect 95700 71334 95752 71340
rect 95240 70032 95292 70038
rect 95240 69974 95292 69980
rect 95252 68882 95280 69974
rect 95712 69970 95740 71334
rect 95700 69964 95752 69970
rect 95700 69906 95752 69912
rect 95896 69358 95924 78610
rect 96374 77820 96682 77829
rect 96374 77818 96380 77820
rect 96436 77818 96460 77820
rect 96516 77818 96540 77820
rect 96596 77818 96620 77820
rect 96676 77818 96682 77820
rect 96436 77766 96438 77818
rect 96618 77766 96620 77818
rect 96374 77764 96380 77766
rect 96436 77764 96460 77766
rect 96516 77764 96540 77766
rect 96596 77764 96620 77766
rect 96676 77764 96682 77766
rect 96374 77755 96682 77764
rect 96528 77648 96580 77654
rect 96528 77590 96580 77596
rect 96540 77110 96568 77590
rect 96528 77104 96580 77110
rect 96528 77046 96580 77052
rect 96374 76732 96682 76741
rect 96374 76730 96380 76732
rect 96436 76730 96460 76732
rect 96516 76730 96540 76732
rect 96596 76730 96620 76732
rect 96676 76730 96682 76732
rect 96436 76678 96438 76730
rect 96618 76678 96620 76730
rect 96374 76676 96380 76678
rect 96436 76676 96460 76678
rect 96516 76676 96540 76678
rect 96596 76676 96620 76678
rect 96676 76676 96682 76678
rect 96374 76667 96682 76676
rect 96374 75644 96682 75653
rect 96374 75642 96380 75644
rect 96436 75642 96460 75644
rect 96516 75642 96540 75644
rect 96596 75642 96620 75644
rect 96676 75642 96682 75644
rect 96436 75590 96438 75642
rect 96618 75590 96620 75642
rect 96374 75588 96380 75590
rect 96436 75588 96460 75590
rect 96516 75588 96540 75590
rect 96596 75588 96620 75590
rect 96676 75588 96682 75590
rect 96374 75579 96682 75588
rect 96816 75546 96844 79154
rect 97908 77716 97960 77722
rect 97908 77658 97960 77664
rect 96896 77512 96948 77518
rect 96896 77454 96948 77460
rect 96908 77178 96936 77454
rect 97920 77450 97948 77658
rect 97908 77444 97960 77450
rect 97908 77386 97960 77392
rect 97632 77376 97684 77382
rect 97632 77318 97684 77324
rect 97034 77276 97342 77285
rect 97034 77274 97040 77276
rect 97096 77274 97120 77276
rect 97176 77274 97200 77276
rect 97256 77274 97280 77276
rect 97336 77274 97342 77276
rect 97096 77222 97098 77274
rect 97278 77222 97280 77274
rect 97034 77220 97040 77222
rect 97096 77220 97120 77222
rect 97176 77220 97200 77222
rect 97256 77220 97280 77222
rect 97336 77220 97342 77222
rect 97034 77211 97342 77220
rect 97644 77178 97672 77318
rect 96896 77172 96948 77178
rect 96896 77114 96948 77120
rect 97632 77172 97684 77178
rect 97632 77114 97684 77120
rect 98012 76634 98040 79630
rect 101968 77926 101996 80038
rect 102060 78674 102088 92195
rect 102048 78668 102100 78674
rect 102048 78610 102100 78616
rect 102152 77994 102180 136818
rect 105922 136572 106230 136581
rect 105922 136570 105928 136572
rect 105984 136570 106008 136572
rect 106064 136570 106088 136572
rect 106144 136570 106168 136572
rect 106224 136570 106230 136572
rect 105984 136518 105986 136570
rect 106166 136518 106168 136570
rect 105922 136516 105928 136518
rect 105984 136516 106008 136518
rect 106064 136516 106088 136518
rect 106144 136516 106168 136518
rect 106224 136516 106230 136518
rect 105922 136507 106230 136516
rect 104348 136128 104400 136134
rect 104348 136070 104400 136076
rect 103704 135924 103756 135930
rect 103704 135866 103756 135872
rect 102232 135856 102284 135862
rect 102232 135798 102284 135804
rect 102140 77988 102192 77994
rect 102140 77930 102192 77936
rect 101956 77920 102008 77926
rect 101956 77862 102008 77868
rect 99104 77716 99156 77722
rect 99104 77658 99156 77664
rect 99116 77382 99144 77658
rect 99104 77376 99156 77382
rect 99104 77318 99156 77324
rect 98736 77104 98788 77110
rect 98736 77046 98788 77052
rect 98460 76832 98512 76838
rect 98460 76774 98512 76780
rect 98000 76628 98052 76634
rect 98000 76570 98052 76576
rect 98276 76492 98328 76498
rect 98276 76434 98328 76440
rect 97724 76356 97776 76362
rect 97724 76298 97776 76304
rect 98184 76356 98236 76362
rect 98184 76298 98236 76304
rect 97034 76188 97342 76197
rect 97034 76186 97040 76188
rect 97096 76186 97120 76188
rect 97176 76186 97200 76188
rect 97256 76186 97280 76188
rect 97336 76186 97342 76188
rect 97096 76134 97098 76186
rect 97278 76134 97280 76186
rect 97034 76132 97040 76134
rect 97096 76132 97120 76134
rect 97176 76132 97200 76134
rect 97256 76132 97280 76134
rect 97336 76132 97342 76134
rect 97034 76123 97342 76132
rect 97736 75954 97764 76298
rect 96896 75948 96948 75954
rect 97724 75948 97776 75954
rect 96896 75890 96948 75896
rect 97644 75908 97724 75936
rect 96804 75540 96856 75546
rect 96804 75482 96856 75488
rect 96908 75410 96936 75890
rect 97540 75744 97592 75750
rect 97540 75686 97592 75692
rect 96896 75404 96948 75410
rect 96896 75346 96948 75352
rect 96804 75200 96856 75206
rect 96804 75142 96856 75148
rect 96712 74792 96764 74798
rect 96712 74734 96764 74740
rect 96374 74556 96682 74565
rect 96374 74554 96380 74556
rect 96436 74554 96460 74556
rect 96516 74554 96540 74556
rect 96596 74554 96620 74556
rect 96676 74554 96682 74556
rect 96436 74502 96438 74554
rect 96618 74502 96620 74554
rect 96374 74500 96380 74502
rect 96436 74500 96460 74502
rect 96516 74500 96540 74502
rect 96596 74500 96620 74502
rect 96676 74500 96682 74502
rect 96374 74491 96682 74500
rect 96724 74458 96752 74734
rect 96712 74452 96764 74458
rect 96712 74394 96764 74400
rect 96816 74322 96844 75142
rect 96908 75002 96936 75346
rect 97448 75200 97500 75206
rect 97448 75142 97500 75148
rect 97034 75100 97342 75109
rect 97034 75098 97040 75100
rect 97096 75098 97120 75100
rect 97176 75098 97200 75100
rect 97256 75098 97280 75100
rect 97336 75098 97342 75100
rect 97096 75046 97098 75098
rect 97278 75046 97280 75098
rect 97034 75044 97040 75046
rect 97096 75044 97120 75046
rect 97176 75044 97200 75046
rect 97256 75044 97280 75046
rect 97336 75044 97342 75046
rect 97034 75035 97342 75044
rect 97460 75002 97488 75142
rect 96896 74996 96948 75002
rect 96896 74938 96948 74944
rect 97448 74996 97500 75002
rect 97448 74938 97500 74944
rect 97552 74866 97580 75686
rect 97356 74860 97408 74866
rect 97356 74802 97408 74808
rect 97540 74860 97592 74866
rect 97540 74802 97592 74808
rect 97368 74662 97396 74802
rect 96896 74656 96948 74662
rect 96896 74598 96948 74604
rect 97356 74656 97408 74662
rect 97356 74598 97408 74604
rect 96804 74316 96856 74322
rect 96804 74258 96856 74264
rect 96374 73468 96682 73477
rect 96374 73466 96380 73468
rect 96436 73466 96460 73468
rect 96516 73466 96540 73468
rect 96596 73466 96620 73468
rect 96676 73466 96682 73468
rect 96436 73414 96438 73466
rect 96618 73414 96620 73466
rect 96374 73412 96380 73414
rect 96436 73412 96460 73414
rect 96516 73412 96540 73414
rect 96596 73412 96620 73414
rect 96676 73412 96682 73414
rect 96374 73403 96682 73412
rect 96908 73166 96936 74598
rect 97644 74338 97672 75908
rect 97724 75890 97776 75896
rect 98000 75880 98052 75886
rect 98000 75822 98052 75828
rect 98012 75546 98040 75822
rect 98196 75818 98224 76298
rect 98184 75812 98236 75818
rect 98184 75754 98236 75760
rect 98000 75540 98052 75546
rect 98000 75482 98052 75488
rect 97724 75472 97776 75478
rect 97724 75414 97776 75420
rect 97736 74866 97764 75414
rect 98288 75342 98316 76434
rect 98472 76430 98500 76774
rect 98460 76424 98512 76430
rect 98460 76366 98512 76372
rect 98644 76424 98696 76430
rect 98644 76366 98696 76372
rect 98472 76022 98500 76366
rect 98460 76016 98512 76022
rect 98460 75958 98512 75964
rect 98656 75954 98684 76366
rect 98748 75954 98776 77046
rect 99104 77036 99156 77042
rect 99104 76978 99156 76984
rect 99288 77036 99340 77042
rect 99288 76978 99340 76984
rect 100116 77036 100168 77042
rect 100116 76978 100168 76984
rect 100760 77036 100812 77042
rect 100760 76978 100812 76984
rect 99116 76634 99144 76978
rect 99196 76968 99248 76974
rect 99196 76910 99248 76916
rect 99104 76628 99156 76634
rect 99104 76570 99156 76576
rect 99012 76424 99064 76430
rect 99012 76366 99064 76372
rect 99024 75954 99052 76366
rect 99208 76362 99236 76910
rect 99300 76566 99328 76978
rect 99288 76560 99340 76566
rect 99288 76502 99340 76508
rect 99196 76356 99248 76362
rect 99196 76298 99248 76304
rect 98552 75948 98604 75954
rect 98552 75890 98604 75896
rect 98644 75948 98696 75954
rect 98644 75890 98696 75896
rect 98736 75948 98788 75954
rect 98736 75890 98788 75896
rect 99012 75948 99064 75954
rect 99012 75890 99064 75896
rect 98460 75880 98512 75886
rect 98460 75822 98512 75828
rect 98368 75744 98420 75750
rect 98368 75686 98420 75692
rect 98380 75342 98408 75686
rect 98276 75336 98328 75342
rect 98276 75278 98328 75284
rect 98368 75336 98420 75342
rect 98368 75278 98420 75284
rect 97908 75268 97960 75274
rect 97908 75210 97960 75216
rect 97920 75002 97948 75210
rect 98000 75200 98052 75206
rect 98000 75142 98052 75148
rect 98184 75200 98236 75206
rect 98184 75142 98236 75148
rect 97908 74996 97960 75002
rect 97908 74938 97960 74944
rect 97724 74860 97776 74866
rect 97724 74802 97776 74808
rect 97908 74792 97960 74798
rect 98012 74780 98040 75142
rect 97960 74752 98040 74780
rect 97908 74734 97960 74740
rect 97816 74656 97868 74662
rect 97816 74598 97868 74604
rect 97908 74656 97960 74662
rect 97908 74598 97960 74604
rect 97552 74310 97672 74338
rect 97448 74248 97500 74254
rect 97448 74190 97500 74196
rect 97034 74012 97342 74021
rect 97034 74010 97040 74012
rect 97096 74010 97120 74012
rect 97176 74010 97200 74012
rect 97256 74010 97280 74012
rect 97336 74010 97342 74012
rect 97096 73958 97098 74010
rect 97278 73958 97280 74010
rect 97034 73956 97040 73958
rect 97096 73956 97120 73958
rect 97176 73956 97200 73958
rect 97256 73956 97280 73958
rect 97336 73956 97342 73958
rect 97034 73947 97342 73956
rect 97460 73778 97488 74190
rect 97448 73772 97500 73778
rect 97448 73714 97500 73720
rect 97552 73166 97580 74310
rect 97724 74112 97776 74118
rect 97724 74054 97776 74060
rect 97736 73302 97764 74054
rect 97828 73846 97856 74598
rect 97920 74254 97948 74598
rect 98012 74322 98040 74752
rect 98000 74316 98052 74322
rect 98000 74258 98052 74264
rect 97908 74248 97960 74254
rect 97908 74190 97960 74196
rect 98196 73914 98224 75142
rect 98368 74860 98420 74866
rect 98368 74802 98420 74808
rect 98380 74458 98408 74802
rect 98472 74730 98500 75822
rect 98564 74934 98592 75890
rect 98656 75818 98684 75890
rect 98644 75812 98696 75818
rect 98644 75754 98696 75760
rect 98748 75806 99236 75834
rect 98656 75546 98684 75754
rect 98644 75540 98696 75546
rect 98644 75482 98696 75488
rect 98748 75426 98776 75806
rect 99208 75750 99236 75806
rect 99104 75744 99156 75750
rect 99104 75686 99156 75692
rect 99196 75744 99248 75750
rect 99196 75686 99248 75692
rect 98656 75398 98776 75426
rect 98552 74928 98604 74934
rect 98552 74870 98604 74876
rect 98460 74724 98512 74730
rect 98460 74666 98512 74672
rect 98368 74452 98420 74458
rect 98368 74394 98420 74400
rect 98656 74390 98684 75398
rect 98736 75268 98788 75274
rect 98736 75210 98788 75216
rect 98644 74384 98696 74390
rect 98644 74326 98696 74332
rect 98276 74248 98328 74254
rect 98276 74190 98328 74196
rect 98644 74248 98696 74254
rect 98644 74190 98696 74196
rect 98184 73908 98236 73914
rect 98184 73850 98236 73856
rect 98288 73846 98316 74190
rect 97816 73840 97868 73846
rect 97816 73782 97868 73788
rect 98276 73840 98328 73846
rect 98276 73782 98328 73788
rect 97724 73296 97776 73302
rect 97724 73238 97776 73244
rect 97736 73166 97764 73238
rect 96896 73160 96948 73166
rect 96896 73102 96948 73108
rect 97540 73160 97592 73166
rect 97540 73102 97592 73108
rect 97724 73160 97776 73166
rect 97724 73102 97776 73108
rect 97552 73030 97580 73102
rect 96160 73024 96212 73030
rect 96160 72966 96212 72972
rect 97448 73024 97500 73030
rect 97448 72966 97500 72972
rect 97540 73024 97592 73030
rect 97540 72966 97592 72972
rect 96068 72752 96120 72758
rect 96068 72694 96120 72700
rect 96080 69766 96108 72694
rect 96172 71670 96200 72966
rect 97034 72924 97342 72933
rect 97034 72922 97040 72924
rect 97096 72922 97120 72924
rect 97176 72922 97200 72924
rect 97256 72922 97280 72924
rect 97336 72922 97342 72924
rect 97096 72870 97098 72922
rect 97278 72870 97280 72922
rect 97034 72868 97040 72870
rect 97096 72868 97120 72870
rect 97176 72868 97200 72870
rect 97256 72868 97280 72870
rect 97336 72868 97342 72870
rect 97034 72859 97342 72868
rect 96374 72380 96682 72389
rect 96374 72378 96380 72380
rect 96436 72378 96460 72380
rect 96516 72378 96540 72380
rect 96596 72378 96620 72380
rect 96676 72378 96682 72380
rect 96436 72326 96438 72378
rect 96618 72326 96620 72378
rect 96374 72324 96380 72326
rect 96436 72324 96460 72326
rect 96516 72324 96540 72326
rect 96596 72324 96620 72326
rect 96676 72324 96682 72326
rect 96374 72315 96682 72324
rect 96804 72140 96856 72146
rect 96804 72082 96856 72088
rect 96712 72072 96764 72078
rect 96712 72014 96764 72020
rect 96160 71664 96212 71670
rect 96160 71606 96212 71612
rect 96172 69902 96200 71606
rect 96374 71292 96682 71301
rect 96374 71290 96380 71292
rect 96436 71290 96460 71292
rect 96516 71290 96540 71292
rect 96596 71290 96620 71292
rect 96676 71290 96682 71292
rect 96436 71238 96438 71290
rect 96618 71238 96620 71290
rect 96374 71236 96380 71238
rect 96436 71236 96460 71238
rect 96516 71236 96540 71238
rect 96596 71236 96620 71238
rect 96676 71236 96682 71238
rect 96374 71227 96682 71236
rect 96724 71194 96752 72014
rect 96816 71738 96844 72082
rect 97034 71836 97342 71845
rect 97034 71834 97040 71836
rect 97096 71834 97120 71836
rect 97176 71834 97200 71836
rect 97256 71834 97280 71836
rect 97336 71834 97342 71836
rect 97096 71782 97098 71834
rect 97278 71782 97280 71834
rect 97034 71780 97040 71782
rect 97096 71780 97120 71782
rect 97176 71780 97200 71782
rect 97256 71780 97280 71782
rect 97336 71780 97342 71782
rect 97034 71771 97342 71780
rect 96804 71732 96856 71738
rect 96804 71674 96856 71680
rect 97460 71466 97488 72966
rect 97632 72752 97684 72758
rect 97632 72694 97684 72700
rect 97644 72486 97672 72694
rect 97724 72684 97776 72690
rect 97828 72672 97856 73782
rect 98460 73772 98512 73778
rect 98460 73714 98512 73720
rect 98368 73704 98420 73710
rect 98368 73646 98420 73652
rect 98092 73160 98144 73166
rect 98092 73102 98144 73108
rect 98184 73160 98236 73166
rect 98184 73102 98236 73108
rect 97908 73092 97960 73098
rect 97908 73034 97960 73040
rect 97920 72826 97948 73034
rect 97908 72820 97960 72826
rect 97908 72762 97960 72768
rect 97776 72644 97856 72672
rect 97724 72626 97776 72632
rect 97632 72480 97684 72486
rect 97632 72422 97684 72428
rect 97632 72208 97684 72214
rect 97632 72150 97684 72156
rect 97540 71596 97592 71602
rect 97540 71538 97592 71544
rect 97448 71460 97500 71466
rect 97448 71402 97500 71408
rect 96712 71188 96764 71194
rect 96712 71130 96764 71136
rect 96804 70984 96856 70990
rect 96804 70926 96856 70932
rect 96816 70446 96844 70926
rect 97552 70854 97580 71538
rect 97644 71466 97672 72150
rect 97736 71584 97764 72626
rect 98104 72622 98132 73102
rect 98196 72826 98224 73102
rect 98276 73024 98328 73030
rect 98276 72966 98328 72972
rect 98184 72820 98236 72826
rect 98184 72762 98236 72768
rect 98092 72616 98144 72622
rect 98092 72558 98144 72564
rect 98288 72554 98316 72966
rect 98380 72690 98408 73646
rect 98472 73302 98500 73714
rect 98656 73642 98684 74190
rect 98748 73642 98776 75210
rect 99116 75002 99144 75686
rect 99196 75540 99248 75546
rect 99196 75482 99248 75488
rect 99104 74996 99156 75002
rect 99104 74938 99156 74944
rect 98826 74216 98882 74225
rect 98826 74151 98882 74160
rect 98840 73914 98868 74151
rect 98920 74112 98972 74118
rect 98920 74054 98972 74060
rect 98932 73914 98960 74054
rect 98828 73908 98880 73914
rect 98828 73850 98880 73856
rect 98920 73908 98972 73914
rect 98920 73850 98972 73856
rect 99012 73772 99064 73778
rect 99116 73760 99144 74938
rect 99208 74798 99236 75482
rect 99300 75478 99328 76502
rect 99564 76356 99616 76362
rect 99564 76298 99616 76304
rect 99576 75954 99604 76298
rect 100024 76288 100076 76294
rect 100024 76230 100076 76236
rect 100036 75954 100064 76230
rect 99564 75948 99616 75954
rect 99564 75890 99616 75896
rect 100024 75948 100076 75954
rect 100024 75890 100076 75896
rect 99288 75472 99340 75478
rect 99288 75414 99340 75420
rect 100036 75342 100064 75890
rect 99380 75336 99432 75342
rect 99380 75278 99432 75284
rect 100024 75336 100076 75342
rect 100024 75278 100076 75284
rect 99288 74860 99340 74866
rect 99288 74802 99340 74808
rect 99196 74792 99248 74798
rect 99196 74734 99248 74740
rect 99300 74458 99328 74802
rect 99288 74452 99340 74458
rect 99288 74394 99340 74400
rect 99196 74180 99248 74186
rect 99196 74122 99248 74128
rect 99064 73732 99144 73760
rect 99012 73714 99064 73720
rect 98644 73636 98696 73642
rect 98644 73578 98696 73584
rect 98736 73636 98788 73642
rect 98736 73578 98788 73584
rect 98550 73400 98606 73409
rect 98550 73335 98552 73344
rect 98604 73335 98606 73344
rect 98552 73306 98604 73312
rect 98460 73296 98512 73302
rect 98460 73238 98512 73244
rect 98748 72842 98776 73578
rect 99116 73273 99144 73732
rect 99102 73264 99158 73273
rect 99102 73199 99158 73208
rect 99208 73030 99236 74122
rect 99392 73778 99420 75278
rect 99472 75268 99524 75274
rect 99472 75210 99524 75216
rect 99932 75268 99984 75274
rect 99932 75210 99984 75216
rect 99484 74934 99512 75210
rect 99472 74928 99524 74934
rect 99524 74876 99604 74882
rect 99472 74870 99604 74876
rect 99484 74854 99604 74870
rect 99944 74866 99972 75210
rect 100036 74866 100064 75278
rect 100128 75002 100156 76978
rect 100576 76968 100628 76974
rect 100576 76910 100628 76916
rect 100392 76424 100444 76430
rect 100392 76366 100444 76372
rect 100404 75886 100432 76366
rect 100588 76090 100616 76910
rect 100772 76090 100800 76978
rect 101036 76832 101088 76838
rect 101036 76774 101088 76780
rect 101048 76498 101076 76774
rect 102244 76537 102272 135798
rect 103612 135720 103664 135726
rect 103612 135662 103664 135668
rect 103520 135652 103572 135658
rect 103520 135594 103572 135600
rect 102784 135516 102836 135522
rect 102784 135458 102836 135464
rect 102324 135448 102376 135454
rect 102324 135390 102376 135396
rect 102336 78198 102364 135390
rect 102796 96626 102824 135458
rect 102876 113280 102928 113286
rect 102876 113222 102928 113228
rect 102784 96620 102836 96626
rect 102784 96562 102836 96568
rect 102508 95192 102560 95198
rect 102508 95134 102560 95140
rect 102520 95097 102548 95134
rect 102506 95088 102562 95097
rect 102506 95023 102562 95032
rect 102416 93696 102468 93702
rect 102416 93638 102468 93644
rect 102428 93397 102456 93638
rect 102414 93388 102470 93397
rect 102414 93323 102470 93332
rect 102520 84194 102548 95023
rect 102784 91112 102836 91118
rect 102784 91054 102836 91060
rect 102428 84166 102548 84194
rect 102324 78192 102376 78198
rect 102324 78134 102376 78140
rect 102428 78062 102456 84166
rect 102796 79354 102824 91054
rect 102888 79490 102916 113222
rect 102968 96144 103020 96150
rect 102968 96086 103020 96092
rect 102876 79484 102928 79490
rect 102876 79426 102928 79432
rect 102980 79422 103008 96086
rect 102968 79416 103020 79422
rect 102968 79358 103020 79364
rect 102784 79348 102836 79354
rect 102784 79290 102836 79296
rect 102416 78056 102468 78062
rect 102416 77998 102468 78004
rect 102230 76528 102286 76537
rect 100944 76492 100996 76498
rect 100944 76434 100996 76440
rect 101036 76492 101088 76498
rect 102230 76463 102286 76472
rect 101036 76434 101088 76440
rect 100576 76084 100628 76090
rect 100576 76026 100628 76032
rect 100760 76084 100812 76090
rect 100760 76026 100812 76032
rect 100208 75880 100260 75886
rect 100208 75822 100260 75828
rect 100392 75880 100444 75886
rect 100392 75822 100444 75828
rect 100116 74996 100168 75002
rect 100116 74938 100168 74944
rect 99472 74792 99524 74798
rect 99472 74734 99524 74740
rect 99484 74497 99512 74734
rect 99470 74488 99526 74497
rect 99470 74423 99526 74432
rect 99288 73772 99340 73778
rect 99288 73714 99340 73720
rect 99380 73772 99432 73778
rect 99380 73714 99432 73720
rect 99300 73370 99328 73714
rect 99472 73636 99524 73642
rect 99472 73578 99524 73584
rect 99484 73409 99512 73578
rect 99470 73400 99526 73409
rect 99288 73364 99340 73370
rect 99576 73370 99604 74854
rect 99932 74860 99984 74866
rect 99932 74802 99984 74808
rect 100024 74860 100076 74866
rect 100024 74802 100076 74808
rect 99840 74792 99892 74798
rect 99840 74734 99892 74740
rect 99656 74656 99708 74662
rect 99656 74598 99708 74604
rect 99668 73710 99696 74598
rect 99748 74180 99800 74186
rect 99748 74122 99800 74128
rect 99760 73914 99788 74122
rect 99748 73908 99800 73914
rect 99748 73850 99800 73856
rect 99656 73704 99708 73710
rect 99656 73646 99708 73652
rect 99470 73335 99526 73344
rect 99564 73364 99616 73370
rect 99288 73306 99340 73312
rect 99564 73306 99616 73312
rect 99196 73024 99248 73030
rect 99196 72966 99248 72972
rect 98656 72814 98776 72842
rect 98460 72752 98512 72758
rect 98460 72694 98512 72700
rect 98368 72684 98420 72690
rect 98368 72626 98420 72632
rect 98276 72548 98328 72554
rect 98276 72490 98328 72496
rect 98000 72072 98052 72078
rect 98000 72014 98052 72020
rect 98092 72072 98144 72078
rect 98092 72014 98144 72020
rect 97908 71596 97960 71602
rect 97736 71556 97908 71584
rect 97908 71538 97960 71544
rect 97632 71460 97684 71466
rect 97632 71402 97684 71408
rect 96896 70848 96948 70854
rect 96896 70790 96948 70796
rect 97540 70848 97592 70854
rect 97540 70790 97592 70796
rect 96908 70632 96936 70790
rect 97034 70748 97342 70757
rect 97034 70746 97040 70748
rect 97096 70746 97120 70748
rect 97176 70746 97200 70748
rect 97256 70746 97280 70748
rect 97336 70746 97342 70748
rect 97096 70694 97098 70746
rect 97278 70694 97280 70746
rect 97034 70692 97040 70694
rect 97096 70692 97120 70694
rect 97176 70692 97200 70694
rect 97256 70692 97280 70694
rect 97336 70692 97342 70694
rect 97034 70683 97342 70692
rect 97080 70644 97132 70650
rect 96908 70604 97080 70632
rect 97080 70586 97132 70592
rect 97092 70514 97120 70586
rect 97080 70508 97132 70514
rect 97080 70450 97132 70456
rect 97264 70508 97316 70514
rect 97264 70450 97316 70456
rect 96804 70440 96856 70446
rect 96804 70382 96856 70388
rect 96374 70204 96682 70213
rect 96374 70202 96380 70204
rect 96436 70202 96460 70204
rect 96516 70202 96540 70204
rect 96596 70202 96620 70204
rect 96676 70202 96682 70204
rect 96436 70150 96438 70202
rect 96618 70150 96620 70202
rect 96374 70148 96380 70150
rect 96436 70148 96460 70150
rect 96516 70148 96540 70150
rect 96596 70148 96620 70150
rect 96676 70148 96682 70150
rect 96374 70139 96682 70148
rect 97276 70038 97304 70450
rect 97448 70440 97500 70446
rect 97448 70382 97500 70388
rect 97264 70032 97316 70038
rect 97264 69974 97316 69980
rect 96160 69896 96212 69902
rect 96160 69838 96212 69844
rect 96068 69760 96120 69766
rect 96068 69702 96120 69708
rect 95884 69352 95936 69358
rect 95884 69294 95936 69300
rect 95976 69012 96028 69018
rect 95976 68954 96028 68960
rect 95240 68876 95292 68882
rect 95240 68818 95292 68824
rect 95516 68876 95568 68882
rect 95516 68818 95568 68824
rect 95148 68672 95200 68678
rect 95148 68614 95200 68620
rect 95056 68264 95108 68270
rect 95056 68206 95108 68212
rect 95160 68134 95188 68614
rect 95240 68332 95292 68338
rect 95240 68274 95292 68280
rect 95148 68128 95200 68134
rect 95148 68070 95200 68076
rect 94964 67788 95016 67794
rect 94964 67730 95016 67736
rect 94976 65958 95004 67730
rect 95252 67386 95280 68274
rect 95332 68128 95384 68134
rect 95332 68070 95384 68076
rect 95344 67726 95372 68070
rect 95332 67720 95384 67726
rect 95332 67662 95384 67668
rect 95332 67584 95384 67590
rect 95332 67526 95384 67532
rect 95240 67380 95292 67386
rect 95240 67322 95292 67328
rect 95240 66700 95292 66706
rect 95240 66642 95292 66648
rect 95252 66230 95280 66642
rect 95240 66224 95292 66230
rect 95240 66166 95292 66172
rect 95344 66162 95372 67526
rect 95528 67182 95556 68818
rect 95792 68196 95844 68202
rect 95792 68138 95844 68144
rect 95700 67788 95752 67794
rect 95700 67730 95752 67736
rect 95516 67176 95568 67182
rect 95516 67118 95568 67124
rect 95712 66842 95740 67730
rect 95700 66836 95752 66842
rect 95700 66778 95752 66784
rect 95608 66632 95660 66638
rect 95608 66574 95660 66580
rect 95424 66496 95476 66502
rect 95424 66438 95476 66444
rect 95436 66298 95464 66438
rect 95620 66298 95648 66574
rect 95804 66298 95832 68138
rect 95884 68128 95936 68134
rect 95884 68070 95936 68076
rect 95896 67794 95924 68070
rect 95884 67788 95936 67794
rect 95884 67730 95936 67736
rect 95988 67250 96016 68954
rect 96080 68814 96108 69702
rect 96172 68882 96200 69838
rect 97460 69834 97488 70382
rect 97552 70106 97580 70790
rect 97644 70446 97672 71402
rect 97908 71392 97960 71398
rect 97908 71334 97960 71340
rect 97724 71120 97776 71126
rect 97722 71088 97724 71097
rect 97776 71088 97778 71097
rect 97722 71023 97778 71032
rect 97724 70984 97776 70990
rect 97776 70944 97856 70972
rect 97724 70926 97776 70932
rect 97828 70514 97856 70944
rect 97920 70938 97948 71334
rect 98012 71058 98040 72014
rect 98104 71738 98132 72014
rect 98092 71732 98144 71738
rect 98092 71674 98144 71680
rect 98288 71618 98316 72490
rect 98380 72010 98408 72626
rect 98472 72214 98500 72694
rect 98552 72616 98604 72622
rect 98552 72558 98604 72564
rect 98460 72208 98512 72214
rect 98460 72150 98512 72156
rect 98564 72078 98592 72558
rect 98552 72072 98604 72078
rect 98552 72014 98604 72020
rect 98368 72004 98420 72010
rect 98368 71946 98420 71952
rect 98656 71942 98684 72814
rect 98736 72684 98788 72690
rect 98736 72626 98788 72632
rect 98748 72146 98776 72626
rect 99576 72622 99604 73306
rect 99654 73264 99710 73273
rect 99654 73199 99710 73208
rect 99668 73166 99696 73199
rect 99656 73160 99708 73166
rect 99852 73114 99880 74734
rect 99944 74322 99972 74802
rect 99932 74316 99984 74322
rect 99932 74258 99984 74264
rect 99944 74118 99972 74258
rect 99932 74112 99984 74118
rect 99932 74054 99984 74060
rect 99932 73908 99984 73914
rect 99932 73850 99984 73856
rect 99944 73234 99972 73850
rect 99932 73228 99984 73234
rect 99932 73170 99984 73176
rect 99656 73102 99708 73108
rect 99760 73086 99880 73114
rect 99564 72616 99616 72622
rect 99564 72558 99616 72564
rect 99104 72276 99156 72282
rect 99104 72218 99156 72224
rect 98736 72140 98788 72146
rect 98736 72082 98788 72088
rect 98644 71936 98696 71942
rect 98644 71878 98696 71884
rect 99012 71936 99064 71942
rect 99012 71878 99064 71884
rect 98920 71732 98972 71738
rect 98920 71674 98972 71680
rect 98104 71590 98316 71618
rect 98552 71664 98604 71670
rect 98552 71606 98604 71612
rect 98368 71596 98420 71602
rect 98104 71534 98132 71590
rect 98368 71538 98420 71544
rect 98092 71528 98144 71534
rect 98092 71470 98144 71476
rect 98000 71052 98052 71058
rect 98000 70994 98052 71000
rect 97920 70910 98040 70938
rect 98012 70854 98040 70910
rect 97908 70848 97960 70854
rect 97908 70790 97960 70796
rect 98000 70848 98052 70854
rect 98000 70790 98052 70796
rect 97920 70582 97948 70790
rect 97908 70576 97960 70582
rect 97908 70518 97960 70524
rect 97816 70508 97868 70514
rect 97816 70450 97868 70456
rect 97632 70440 97684 70446
rect 97632 70382 97684 70388
rect 97540 70100 97592 70106
rect 97540 70042 97592 70048
rect 97538 70000 97594 70009
rect 97828 69970 97856 70450
rect 97908 70440 97960 70446
rect 97908 70382 97960 70388
rect 97920 70038 97948 70382
rect 98104 70378 98132 71470
rect 98182 71088 98238 71097
rect 98182 71023 98238 71032
rect 98276 71052 98328 71058
rect 98196 70514 98224 71023
rect 98276 70994 98328 71000
rect 98184 70508 98236 70514
rect 98184 70450 98236 70456
rect 98288 70394 98316 70994
rect 98380 70582 98408 71538
rect 98564 71466 98592 71606
rect 98552 71460 98604 71466
rect 98552 71402 98604 71408
rect 98564 71126 98592 71402
rect 98932 71398 98960 71674
rect 99024 71534 99052 71878
rect 99012 71528 99064 71534
rect 99012 71470 99064 71476
rect 99116 71466 99144 72218
rect 99576 72010 99604 72558
rect 99196 72004 99248 72010
rect 99196 71946 99248 71952
rect 99564 72004 99616 72010
rect 99564 71946 99616 71952
rect 99208 71670 99236 71946
rect 99196 71664 99248 71670
rect 99196 71606 99248 71612
rect 99760 71602 99788 73086
rect 100036 72826 100064 74802
rect 100128 73574 100156 74938
rect 100220 74866 100248 75822
rect 100300 75812 100352 75818
rect 100300 75754 100352 75760
rect 100312 75206 100340 75754
rect 100404 75274 100432 75822
rect 100956 75410 100984 76434
rect 101128 76424 101180 76430
rect 101128 76366 101180 76372
rect 100944 75404 100996 75410
rect 100944 75346 100996 75352
rect 100392 75268 100444 75274
rect 100392 75210 100444 75216
rect 100300 75200 100352 75206
rect 100300 75142 100352 75148
rect 100484 75200 100536 75206
rect 100484 75142 100536 75148
rect 100496 74866 100524 75142
rect 100956 75002 100984 75346
rect 100944 74996 100996 75002
rect 100944 74938 100996 74944
rect 101140 74866 101168 76366
rect 103532 75993 103560 135594
rect 103624 77081 103652 135662
rect 103610 77072 103666 77081
rect 103610 77007 103666 77016
rect 103716 76401 103744 135866
rect 103796 135788 103848 135794
rect 103796 135730 103848 135736
rect 103808 76945 103836 135730
rect 104072 133952 104124 133958
rect 104072 133894 104124 133900
rect 103886 129840 103942 129849
rect 103886 129775 103888 129784
rect 103940 129775 103942 129784
rect 103888 129746 103940 129752
rect 103888 92608 103940 92614
rect 103888 92550 103940 92556
rect 103900 92313 103928 92550
rect 103886 92304 103942 92313
rect 103886 92239 103942 92248
rect 103794 76936 103850 76945
rect 103794 76871 103850 76880
rect 103702 76392 103758 76401
rect 103702 76327 103758 76336
rect 103518 75984 103574 75993
rect 103518 75919 103574 75928
rect 104084 75886 104112 133894
rect 104360 113626 104388 136070
rect 106658 136028 106966 136037
rect 106658 136026 106664 136028
rect 106720 136026 106744 136028
rect 106800 136026 106824 136028
rect 106880 136026 106904 136028
rect 106960 136026 106966 136028
rect 106720 135974 106722 136026
rect 106902 135974 106904 136026
rect 106658 135972 106664 135974
rect 106720 135972 106744 135974
rect 106800 135972 106824 135974
rect 106880 135972 106904 135974
rect 106960 135972 106966 135974
rect 106658 135963 106966 135972
rect 104624 135584 104676 135590
rect 104624 135526 104676 135532
rect 104532 133748 104584 133754
rect 104532 133690 104584 133696
rect 104348 113620 104400 113626
rect 104348 113562 104400 113568
rect 104360 113490 104388 113562
rect 104348 113484 104400 113490
rect 104348 113426 104400 113432
rect 104544 113354 104572 133690
rect 104532 113348 104584 113354
rect 104532 113290 104584 113296
rect 104544 113082 104572 113290
rect 104532 113076 104584 113082
rect 104532 113018 104584 113024
rect 104636 101046 104664 135526
rect 105922 135484 106230 135493
rect 105922 135482 105928 135484
rect 105984 135482 106008 135484
rect 106064 135482 106088 135484
rect 106144 135482 106168 135484
rect 106224 135482 106230 135484
rect 105984 135430 105986 135482
rect 106166 135430 106168 135482
rect 105922 135428 105928 135430
rect 105984 135428 106008 135430
rect 106064 135428 106088 135430
rect 106144 135428 106168 135430
rect 106224 135428 106230 135430
rect 105922 135419 106230 135428
rect 106658 134940 106966 134949
rect 106658 134938 106664 134940
rect 106720 134938 106744 134940
rect 106800 134938 106824 134940
rect 106880 134938 106904 134940
rect 106960 134938 106966 134940
rect 106720 134886 106722 134938
rect 106902 134886 106904 134938
rect 106658 134884 106664 134886
rect 106720 134884 106744 134886
rect 106800 134884 106824 134886
rect 106880 134884 106904 134886
rect 106960 134884 106966 134886
rect 106658 134875 106966 134884
rect 105922 134396 106230 134405
rect 105922 134394 105928 134396
rect 105984 134394 106008 134396
rect 106064 134394 106088 134396
rect 106144 134394 106168 134396
rect 106224 134394 106230 134396
rect 105984 134342 105986 134394
rect 106166 134342 106168 134394
rect 105922 134340 105928 134342
rect 105984 134340 106008 134342
rect 106064 134340 106088 134342
rect 106144 134340 106168 134342
rect 106224 134340 106230 134342
rect 105922 134331 106230 134340
rect 106658 133852 106966 133861
rect 106658 133850 106664 133852
rect 106720 133850 106744 133852
rect 106800 133850 106824 133852
rect 106880 133850 106904 133852
rect 106960 133850 106966 133852
rect 106720 133798 106722 133850
rect 106902 133798 106904 133850
rect 106658 133796 106664 133798
rect 106720 133796 106744 133798
rect 106800 133796 106824 133798
rect 106880 133796 106904 133798
rect 106960 133796 106966 133798
rect 106658 133787 106966 133796
rect 105922 133308 106230 133317
rect 105922 133306 105928 133308
rect 105984 133306 106008 133308
rect 106064 133306 106088 133308
rect 106144 133306 106168 133308
rect 106224 133306 106230 133308
rect 105984 133254 105986 133306
rect 106166 133254 106168 133306
rect 105922 133252 105928 133254
rect 105984 133252 106008 133254
rect 106064 133252 106088 133254
rect 106144 133252 106168 133254
rect 106224 133252 106230 133254
rect 105922 133243 106230 133252
rect 106658 132764 106966 132773
rect 106658 132762 106664 132764
rect 106720 132762 106744 132764
rect 106800 132762 106824 132764
rect 106880 132762 106904 132764
rect 106960 132762 106966 132764
rect 106720 132710 106722 132762
rect 106902 132710 106904 132762
rect 106658 132708 106664 132710
rect 106720 132708 106744 132710
rect 106800 132708 106824 132710
rect 106880 132708 106904 132710
rect 106960 132708 106966 132710
rect 106658 132699 106966 132708
rect 105922 132220 106230 132229
rect 105922 132218 105928 132220
rect 105984 132218 106008 132220
rect 106064 132218 106088 132220
rect 106144 132218 106168 132220
rect 106224 132218 106230 132220
rect 105984 132166 105986 132218
rect 106166 132166 106168 132218
rect 105922 132164 105928 132166
rect 105984 132164 106008 132166
rect 106064 132164 106088 132166
rect 106144 132164 106168 132166
rect 106224 132164 106230 132166
rect 105922 132155 106230 132164
rect 106658 131676 106966 131685
rect 106658 131674 106664 131676
rect 106720 131674 106744 131676
rect 106800 131674 106824 131676
rect 106880 131674 106904 131676
rect 106960 131674 106966 131676
rect 106720 131622 106722 131674
rect 106902 131622 106904 131674
rect 106658 131620 106664 131622
rect 106720 131620 106744 131622
rect 106800 131620 106824 131622
rect 106880 131620 106904 131622
rect 106960 131620 106966 131622
rect 106658 131611 106966 131620
rect 105922 131132 106230 131141
rect 105922 131130 105928 131132
rect 105984 131130 106008 131132
rect 106064 131130 106088 131132
rect 106144 131130 106168 131132
rect 106224 131130 106230 131132
rect 105984 131078 105986 131130
rect 106166 131078 106168 131130
rect 105922 131076 105928 131078
rect 105984 131076 106008 131078
rect 106064 131076 106088 131078
rect 106144 131076 106168 131078
rect 106224 131076 106230 131078
rect 105922 131067 106230 131076
rect 106658 130588 106966 130597
rect 106658 130586 106664 130588
rect 106720 130586 106744 130588
rect 106800 130586 106824 130588
rect 106880 130586 106904 130588
rect 106960 130586 106966 130588
rect 106720 130534 106722 130586
rect 106902 130534 106904 130586
rect 106658 130532 106664 130534
rect 106720 130532 106744 130534
rect 106800 130532 106824 130534
rect 106880 130532 106904 130534
rect 106960 130532 106966 130534
rect 106658 130523 106966 130532
rect 105922 130044 106230 130053
rect 105922 130042 105928 130044
rect 105984 130042 106008 130044
rect 106064 130042 106088 130044
rect 106144 130042 106168 130044
rect 106224 130042 106230 130044
rect 105984 129990 105986 130042
rect 106166 129990 106168 130042
rect 105922 129988 105928 129990
rect 105984 129988 106008 129990
rect 106064 129988 106088 129990
rect 106144 129988 106168 129990
rect 106224 129988 106230 129990
rect 105922 129979 106230 129988
rect 106658 129500 106966 129509
rect 106658 129498 106664 129500
rect 106720 129498 106744 129500
rect 106800 129498 106824 129500
rect 106880 129498 106904 129500
rect 106960 129498 106966 129500
rect 106720 129446 106722 129498
rect 106902 129446 106904 129498
rect 106658 129444 106664 129446
rect 106720 129444 106744 129446
rect 106800 129444 106824 129446
rect 106880 129444 106904 129446
rect 106960 129444 106966 129446
rect 106658 129435 106966 129444
rect 105922 128956 106230 128965
rect 105922 128954 105928 128956
rect 105984 128954 106008 128956
rect 106064 128954 106088 128956
rect 106144 128954 106168 128956
rect 106224 128954 106230 128956
rect 105984 128902 105986 128954
rect 106166 128902 106168 128954
rect 105922 128900 105928 128902
rect 105984 128900 106008 128902
rect 106064 128900 106088 128902
rect 106144 128900 106168 128902
rect 106224 128900 106230 128902
rect 105922 128891 106230 128900
rect 106658 128412 106966 128421
rect 106658 128410 106664 128412
rect 106720 128410 106744 128412
rect 106800 128410 106824 128412
rect 106880 128410 106904 128412
rect 106960 128410 106966 128412
rect 106720 128358 106722 128410
rect 106902 128358 106904 128410
rect 106658 128356 106664 128358
rect 106720 128356 106744 128358
rect 106800 128356 106824 128358
rect 106880 128356 106904 128358
rect 106960 128356 106966 128358
rect 106658 128347 106966 128356
rect 105922 127868 106230 127877
rect 105922 127866 105928 127868
rect 105984 127866 106008 127868
rect 106064 127866 106088 127868
rect 106144 127866 106168 127868
rect 106224 127866 106230 127868
rect 105984 127814 105986 127866
rect 106166 127814 106168 127866
rect 105922 127812 105928 127814
rect 105984 127812 106008 127814
rect 106064 127812 106088 127814
rect 106144 127812 106168 127814
rect 106224 127812 106230 127814
rect 105922 127803 106230 127812
rect 106658 127324 106966 127333
rect 106658 127322 106664 127324
rect 106720 127322 106744 127324
rect 106800 127322 106824 127324
rect 106880 127322 106904 127324
rect 106960 127322 106966 127324
rect 106720 127270 106722 127322
rect 106902 127270 106904 127322
rect 106658 127268 106664 127270
rect 106720 127268 106744 127270
rect 106800 127268 106824 127270
rect 106880 127268 106904 127270
rect 106960 127268 106966 127270
rect 106658 127259 106966 127268
rect 105922 126780 106230 126789
rect 105922 126778 105928 126780
rect 105984 126778 106008 126780
rect 106064 126778 106088 126780
rect 106144 126778 106168 126780
rect 106224 126778 106230 126780
rect 105984 126726 105986 126778
rect 106166 126726 106168 126778
rect 105922 126724 105928 126726
rect 105984 126724 106008 126726
rect 106064 126724 106088 126726
rect 106144 126724 106168 126726
rect 106224 126724 106230 126726
rect 105922 126715 106230 126724
rect 106658 126236 106966 126245
rect 106658 126234 106664 126236
rect 106720 126234 106744 126236
rect 106800 126234 106824 126236
rect 106880 126234 106904 126236
rect 106960 126234 106966 126236
rect 106720 126182 106722 126234
rect 106902 126182 106904 126234
rect 106658 126180 106664 126182
rect 106720 126180 106744 126182
rect 106800 126180 106824 126182
rect 106880 126180 106904 126182
rect 106960 126180 106966 126182
rect 106658 126171 106966 126180
rect 105922 125692 106230 125701
rect 105922 125690 105928 125692
rect 105984 125690 106008 125692
rect 106064 125690 106088 125692
rect 106144 125690 106168 125692
rect 106224 125690 106230 125692
rect 105984 125638 105986 125690
rect 106166 125638 106168 125690
rect 105922 125636 105928 125638
rect 105984 125636 106008 125638
rect 106064 125636 106088 125638
rect 106144 125636 106168 125638
rect 106224 125636 106230 125638
rect 105922 125627 106230 125636
rect 106658 125148 106966 125157
rect 106658 125146 106664 125148
rect 106720 125146 106744 125148
rect 106800 125146 106824 125148
rect 106880 125146 106904 125148
rect 106960 125146 106966 125148
rect 106720 125094 106722 125146
rect 106902 125094 106904 125146
rect 106658 125092 106664 125094
rect 106720 125092 106744 125094
rect 106800 125092 106824 125094
rect 106880 125092 106904 125094
rect 106960 125092 106966 125094
rect 106658 125083 106966 125092
rect 105922 124604 106230 124613
rect 105922 124602 105928 124604
rect 105984 124602 106008 124604
rect 106064 124602 106088 124604
rect 106144 124602 106168 124604
rect 106224 124602 106230 124604
rect 105984 124550 105986 124602
rect 106166 124550 106168 124602
rect 105922 124548 105928 124550
rect 105984 124548 106008 124550
rect 106064 124548 106088 124550
rect 106144 124548 106168 124550
rect 106224 124548 106230 124550
rect 105922 124539 106230 124548
rect 106658 124060 106966 124069
rect 106658 124058 106664 124060
rect 106720 124058 106744 124060
rect 106800 124058 106824 124060
rect 106880 124058 106904 124060
rect 106960 124058 106966 124060
rect 106720 124006 106722 124058
rect 106902 124006 106904 124058
rect 106658 124004 106664 124006
rect 106720 124004 106744 124006
rect 106800 124004 106824 124006
rect 106880 124004 106904 124006
rect 106960 124004 106966 124006
rect 106658 123995 106966 124004
rect 105922 123516 106230 123525
rect 105922 123514 105928 123516
rect 105984 123514 106008 123516
rect 106064 123514 106088 123516
rect 106144 123514 106168 123516
rect 106224 123514 106230 123516
rect 105984 123462 105986 123514
rect 106166 123462 106168 123514
rect 105922 123460 105928 123462
rect 105984 123460 106008 123462
rect 106064 123460 106088 123462
rect 106144 123460 106168 123462
rect 106224 123460 106230 123462
rect 105922 123451 106230 123460
rect 106658 122972 106966 122981
rect 106658 122970 106664 122972
rect 106720 122970 106744 122972
rect 106800 122970 106824 122972
rect 106880 122970 106904 122972
rect 106960 122970 106966 122972
rect 106720 122918 106722 122970
rect 106902 122918 106904 122970
rect 106658 122916 106664 122918
rect 106720 122916 106744 122918
rect 106800 122916 106824 122918
rect 106880 122916 106904 122918
rect 106960 122916 106966 122918
rect 106658 122907 106966 122916
rect 105922 122428 106230 122437
rect 105922 122426 105928 122428
rect 105984 122426 106008 122428
rect 106064 122426 106088 122428
rect 106144 122426 106168 122428
rect 106224 122426 106230 122428
rect 105984 122374 105986 122426
rect 106166 122374 106168 122426
rect 105922 122372 105928 122374
rect 105984 122372 106008 122374
rect 106064 122372 106088 122374
rect 106144 122372 106168 122374
rect 106224 122372 106230 122374
rect 105922 122363 106230 122372
rect 106658 121884 106966 121893
rect 106658 121882 106664 121884
rect 106720 121882 106744 121884
rect 106800 121882 106824 121884
rect 106880 121882 106904 121884
rect 106960 121882 106966 121884
rect 106720 121830 106722 121882
rect 106902 121830 106904 121882
rect 106658 121828 106664 121830
rect 106720 121828 106744 121830
rect 106800 121828 106824 121830
rect 106880 121828 106904 121830
rect 106960 121828 106966 121830
rect 106658 121819 106966 121828
rect 105922 121340 106230 121349
rect 105922 121338 105928 121340
rect 105984 121338 106008 121340
rect 106064 121338 106088 121340
rect 106144 121338 106168 121340
rect 106224 121338 106230 121340
rect 105984 121286 105986 121338
rect 106166 121286 106168 121338
rect 105922 121284 105928 121286
rect 105984 121284 106008 121286
rect 106064 121284 106088 121286
rect 106144 121284 106168 121286
rect 106224 121284 106230 121286
rect 105922 121275 106230 121284
rect 106658 120796 106966 120805
rect 106658 120794 106664 120796
rect 106720 120794 106744 120796
rect 106800 120794 106824 120796
rect 106880 120794 106904 120796
rect 106960 120794 106966 120796
rect 106720 120742 106722 120794
rect 106902 120742 106904 120794
rect 106658 120740 106664 120742
rect 106720 120740 106744 120742
rect 106800 120740 106824 120742
rect 106880 120740 106904 120742
rect 106960 120740 106966 120742
rect 106658 120731 106966 120740
rect 105922 120252 106230 120261
rect 105922 120250 105928 120252
rect 105984 120250 106008 120252
rect 106064 120250 106088 120252
rect 106144 120250 106168 120252
rect 106224 120250 106230 120252
rect 105984 120198 105986 120250
rect 106166 120198 106168 120250
rect 105922 120196 105928 120198
rect 105984 120196 106008 120198
rect 106064 120196 106088 120198
rect 106144 120196 106168 120198
rect 106224 120196 106230 120198
rect 105922 120187 106230 120196
rect 106658 119708 106966 119717
rect 106658 119706 106664 119708
rect 106720 119706 106744 119708
rect 106800 119706 106824 119708
rect 106880 119706 106904 119708
rect 106960 119706 106966 119708
rect 106720 119654 106722 119706
rect 106902 119654 106904 119706
rect 106658 119652 106664 119654
rect 106720 119652 106744 119654
rect 106800 119652 106824 119654
rect 106880 119652 106904 119654
rect 106960 119652 106966 119654
rect 106658 119643 106966 119652
rect 105922 119164 106230 119173
rect 105922 119162 105928 119164
rect 105984 119162 106008 119164
rect 106064 119162 106088 119164
rect 106144 119162 106168 119164
rect 106224 119162 106230 119164
rect 105984 119110 105986 119162
rect 106166 119110 106168 119162
rect 105922 119108 105928 119110
rect 105984 119108 106008 119110
rect 106064 119108 106088 119110
rect 106144 119108 106168 119110
rect 106224 119108 106230 119110
rect 105922 119099 106230 119108
rect 106658 118620 106966 118629
rect 106658 118618 106664 118620
rect 106720 118618 106744 118620
rect 106800 118618 106824 118620
rect 106880 118618 106904 118620
rect 106960 118618 106966 118620
rect 106720 118566 106722 118618
rect 106902 118566 106904 118618
rect 106658 118564 106664 118566
rect 106720 118564 106744 118566
rect 106800 118564 106824 118566
rect 106880 118564 106904 118566
rect 106960 118564 106966 118566
rect 106658 118555 106966 118564
rect 105922 118076 106230 118085
rect 105922 118074 105928 118076
rect 105984 118074 106008 118076
rect 106064 118074 106088 118076
rect 106144 118074 106168 118076
rect 106224 118074 106230 118076
rect 105984 118022 105986 118074
rect 106166 118022 106168 118074
rect 105922 118020 105928 118022
rect 105984 118020 106008 118022
rect 106064 118020 106088 118022
rect 106144 118020 106168 118022
rect 106224 118020 106230 118022
rect 105922 118011 106230 118020
rect 106658 117532 106966 117541
rect 106658 117530 106664 117532
rect 106720 117530 106744 117532
rect 106800 117530 106824 117532
rect 106880 117530 106904 117532
rect 106960 117530 106966 117532
rect 106720 117478 106722 117530
rect 106902 117478 106904 117530
rect 106658 117476 106664 117478
rect 106720 117476 106744 117478
rect 106800 117476 106824 117478
rect 106880 117476 106904 117478
rect 106960 117476 106966 117478
rect 106658 117467 106966 117476
rect 105922 116988 106230 116997
rect 105922 116986 105928 116988
rect 105984 116986 106008 116988
rect 106064 116986 106088 116988
rect 106144 116986 106168 116988
rect 106224 116986 106230 116988
rect 105984 116934 105986 116986
rect 106166 116934 106168 116986
rect 105922 116932 105928 116934
rect 105984 116932 106008 116934
rect 106064 116932 106088 116934
rect 106144 116932 106168 116934
rect 106224 116932 106230 116934
rect 105922 116923 106230 116932
rect 106658 116444 106966 116453
rect 106658 116442 106664 116444
rect 106720 116442 106744 116444
rect 106800 116442 106824 116444
rect 106880 116442 106904 116444
rect 106960 116442 106966 116444
rect 106720 116390 106722 116442
rect 106902 116390 106904 116442
rect 106658 116388 106664 116390
rect 106720 116388 106744 116390
rect 106800 116388 106824 116390
rect 106880 116388 106904 116390
rect 106960 116388 106966 116390
rect 106658 116379 106966 116388
rect 105922 115900 106230 115909
rect 105922 115898 105928 115900
rect 105984 115898 106008 115900
rect 106064 115898 106088 115900
rect 106144 115898 106168 115900
rect 106224 115898 106230 115900
rect 105984 115846 105986 115898
rect 106166 115846 106168 115898
rect 105922 115844 105928 115846
rect 105984 115844 106008 115846
rect 106064 115844 106088 115846
rect 106144 115844 106168 115846
rect 106224 115844 106230 115846
rect 105922 115835 106230 115844
rect 106658 115356 106966 115365
rect 106658 115354 106664 115356
rect 106720 115354 106744 115356
rect 106800 115354 106824 115356
rect 106880 115354 106904 115356
rect 106960 115354 106966 115356
rect 106720 115302 106722 115354
rect 106902 115302 106904 115354
rect 106658 115300 106664 115302
rect 106720 115300 106744 115302
rect 106800 115300 106824 115302
rect 106880 115300 106904 115302
rect 106960 115300 106966 115302
rect 106658 115291 106966 115300
rect 105922 114812 106230 114821
rect 105922 114810 105928 114812
rect 105984 114810 106008 114812
rect 106064 114810 106088 114812
rect 106144 114810 106168 114812
rect 106224 114810 106230 114812
rect 105984 114758 105986 114810
rect 106166 114758 106168 114810
rect 105922 114756 105928 114758
rect 105984 114756 106008 114758
rect 106064 114756 106088 114758
rect 106144 114756 106168 114758
rect 106224 114756 106230 114758
rect 105922 114747 106230 114756
rect 106658 114268 106966 114277
rect 106658 114266 106664 114268
rect 106720 114266 106744 114268
rect 106800 114266 106824 114268
rect 106880 114266 106904 114268
rect 106960 114266 106966 114268
rect 106720 114214 106722 114266
rect 106902 114214 106904 114266
rect 106658 114212 106664 114214
rect 106720 114212 106744 114214
rect 106800 114212 106824 114214
rect 106880 114212 106904 114214
rect 106960 114212 106966 114214
rect 106658 114203 106966 114212
rect 105922 113724 106230 113733
rect 105922 113722 105928 113724
rect 105984 113722 106008 113724
rect 106064 113722 106088 113724
rect 106144 113722 106168 113724
rect 106224 113722 106230 113724
rect 105984 113670 105986 113722
rect 106166 113670 106168 113722
rect 105922 113668 105928 113670
rect 105984 113668 106008 113670
rect 106064 113668 106088 113670
rect 106144 113668 106168 113670
rect 106224 113668 106230 113670
rect 105922 113659 106230 113668
rect 105636 113620 105688 113626
rect 105636 113562 105688 113568
rect 105648 107098 105676 113562
rect 106658 113180 106966 113189
rect 106658 113178 106664 113180
rect 106720 113178 106744 113180
rect 106800 113178 106824 113180
rect 106880 113178 106904 113180
rect 106960 113178 106966 113180
rect 106720 113126 106722 113178
rect 106902 113126 106904 113178
rect 106658 113124 106664 113126
rect 106720 113124 106744 113126
rect 106800 113124 106824 113126
rect 106880 113124 106904 113126
rect 106960 113124 106966 113126
rect 106658 113115 106966 113124
rect 105922 112636 106230 112645
rect 105922 112634 105928 112636
rect 105984 112634 106008 112636
rect 106064 112634 106088 112636
rect 106144 112634 106168 112636
rect 106224 112634 106230 112636
rect 105984 112582 105986 112634
rect 106166 112582 106168 112634
rect 105922 112580 105928 112582
rect 105984 112580 106008 112582
rect 106064 112580 106088 112582
rect 106144 112580 106168 112582
rect 106224 112580 106230 112582
rect 105922 112571 106230 112580
rect 106658 112092 106966 112101
rect 106658 112090 106664 112092
rect 106720 112090 106744 112092
rect 106800 112090 106824 112092
rect 106880 112090 106904 112092
rect 106960 112090 106966 112092
rect 106720 112038 106722 112090
rect 106902 112038 106904 112090
rect 106658 112036 106664 112038
rect 106720 112036 106744 112038
rect 106800 112036 106824 112038
rect 106880 112036 106904 112038
rect 106960 112036 106966 112038
rect 106658 112027 106966 112036
rect 105922 111548 106230 111557
rect 105922 111546 105928 111548
rect 105984 111546 106008 111548
rect 106064 111546 106088 111548
rect 106144 111546 106168 111548
rect 106224 111546 106230 111548
rect 105984 111494 105986 111546
rect 106166 111494 106168 111546
rect 105922 111492 105928 111494
rect 105984 111492 106008 111494
rect 106064 111492 106088 111494
rect 106144 111492 106168 111494
rect 106224 111492 106230 111494
rect 105922 111483 106230 111492
rect 106658 111004 106966 111013
rect 106658 111002 106664 111004
rect 106720 111002 106744 111004
rect 106800 111002 106824 111004
rect 106880 111002 106904 111004
rect 106960 111002 106966 111004
rect 106720 110950 106722 111002
rect 106902 110950 106904 111002
rect 106658 110948 106664 110950
rect 106720 110948 106744 110950
rect 106800 110948 106824 110950
rect 106880 110948 106904 110950
rect 106960 110948 106966 110950
rect 106658 110939 106966 110948
rect 105922 110460 106230 110469
rect 105922 110458 105928 110460
rect 105984 110458 106008 110460
rect 106064 110458 106088 110460
rect 106144 110458 106168 110460
rect 106224 110458 106230 110460
rect 105984 110406 105986 110458
rect 106166 110406 106168 110458
rect 105922 110404 105928 110406
rect 105984 110404 106008 110406
rect 106064 110404 106088 110406
rect 106144 110404 106168 110406
rect 106224 110404 106230 110406
rect 105922 110395 106230 110404
rect 106658 109916 106966 109925
rect 106658 109914 106664 109916
rect 106720 109914 106744 109916
rect 106800 109914 106824 109916
rect 106880 109914 106904 109916
rect 106960 109914 106966 109916
rect 106720 109862 106722 109914
rect 106902 109862 106904 109914
rect 106658 109860 106664 109862
rect 106720 109860 106744 109862
rect 106800 109860 106824 109862
rect 106880 109860 106904 109862
rect 106960 109860 106966 109862
rect 106658 109851 106966 109860
rect 105922 109372 106230 109381
rect 105922 109370 105928 109372
rect 105984 109370 106008 109372
rect 106064 109370 106088 109372
rect 106144 109370 106168 109372
rect 106224 109370 106230 109372
rect 105984 109318 105986 109370
rect 106166 109318 106168 109370
rect 105922 109316 105928 109318
rect 105984 109316 106008 109318
rect 106064 109316 106088 109318
rect 106144 109316 106168 109318
rect 106224 109316 106230 109318
rect 105922 109307 106230 109316
rect 106658 108828 106966 108837
rect 106658 108826 106664 108828
rect 106720 108826 106744 108828
rect 106800 108826 106824 108828
rect 106880 108826 106904 108828
rect 106960 108826 106966 108828
rect 106720 108774 106722 108826
rect 106902 108774 106904 108826
rect 106658 108772 106664 108774
rect 106720 108772 106744 108774
rect 106800 108772 106824 108774
rect 106880 108772 106904 108774
rect 106960 108772 106966 108774
rect 106658 108763 106966 108772
rect 105922 108284 106230 108293
rect 105922 108282 105928 108284
rect 105984 108282 106008 108284
rect 106064 108282 106088 108284
rect 106144 108282 106168 108284
rect 106224 108282 106230 108284
rect 105984 108230 105986 108282
rect 106166 108230 106168 108282
rect 105922 108228 105928 108230
rect 105984 108228 106008 108230
rect 106064 108228 106088 108230
rect 106144 108228 106168 108230
rect 106224 108228 106230 108230
rect 105922 108219 106230 108228
rect 106658 107740 106966 107749
rect 106658 107738 106664 107740
rect 106720 107738 106744 107740
rect 106800 107738 106824 107740
rect 106880 107738 106904 107740
rect 106960 107738 106966 107740
rect 106720 107686 106722 107738
rect 106902 107686 106904 107738
rect 106658 107684 106664 107686
rect 106720 107684 106744 107686
rect 106800 107684 106824 107686
rect 106880 107684 106904 107686
rect 106960 107684 106966 107686
rect 106658 107675 106966 107684
rect 105922 107196 106230 107205
rect 105922 107194 105928 107196
rect 105984 107194 106008 107196
rect 106064 107194 106088 107196
rect 106144 107194 106168 107196
rect 106224 107194 106230 107196
rect 105984 107142 105986 107194
rect 106166 107142 106168 107194
rect 105922 107140 105928 107142
rect 105984 107140 106008 107142
rect 106064 107140 106088 107142
rect 106144 107140 106168 107142
rect 106224 107140 106230 107142
rect 105922 107131 106230 107140
rect 105636 107092 105688 107098
rect 105636 107034 105688 107040
rect 105820 107092 105872 107098
rect 105820 107034 105872 107040
rect 105084 106820 105136 106826
rect 105084 106762 105136 106768
rect 104624 101040 104676 101046
rect 104624 100982 104676 100988
rect 104636 100570 104664 100982
rect 104624 100564 104676 100570
rect 104624 100506 104676 100512
rect 104348 96552 104400 96558
rect 104348 96494 104400 96500
rect 104360 96422 104388 96494
rect 104348 96416 104400 96422
rect 104348 96358 104400 96364
rect 104360 77722 104388 96358
rect 105096 91594 105124 106762
rect 105832 100910 105860 107034
rect 106658 106652 106966 106661
rect 106658 106650 106664 106652
rect 106720 106650 106744 106652
rect 106800 106650 106824 106652
rect 106880 106650 106904 106652
rect 106960 106650 106966 106652
rect 106720 106598 106722 106650
rect 106902 106598 106904 106650
rect 106658 106596 106664 106598
rect 106720 106596 106744 106598
rect 106800 106596 106824 106598
rect 106880 106596 106904 106598
rect 106960 106596 106966 106598
rect 106658 106587 106966 106596
rect 105922 106108 106230 106117
rect 105922 106106 105928 106108
rect 105984 106106 106008 106108
rect 106064 106106 106088 106108
rect 106144 106106 106168 106108
rect 106224 106106 106230 106108
rect 105984 106054 105986 106106
rect 106166 106054 106168 106106
rect 105922 106052 105928 106054
rect 105984 106052 106008 106054
rect 106064 106052 106088 106054
rect 106144 106052 106168 106054
rect 106224 106052 106230 106054
rect 105922 106043 106230 106052
rect 106658 105564 106966 105573
rect 106658 105562 106664 105564
rect 106720 105562 106744 105564
rect 106800 105562 106824 105564
rect 106880 105562 106904 105564
rect 106960 105562 106966 105564
rect 106720 105510 106722 105562
rect 106902 105510 106904 105562
rect 106658 105508 106664 105510
rect 106720 105508 106744 105510
rect 106800 105508 106824 105510
rect 106880 105508 106904 105510
rect 106960 105508 106966 105510
rect 106658 105499 106966 105508
rect 105922 105020 106230 105029
rect 105922 105018 105928 105020
rect 105984 105018 106008 105020
rect 106064 105018 106088 105020
rect 106144 105018 106168 105020
rect 106224 105018 106230 105020
rect 105984 104966 105986 105018
rect 106166 104966 106168 105018
rect 105922 104964 105928 104966
rect 105984 104964 106008 104966
rect 106064 104964 106088 104966
rect 106144 104964 106168 104966
rect 106224 104964 106230 104966
rect 105922 104955 106230 104964
rect 106658 104476 106966 104485
rect 106658 104474 106664 104476
rect 106720 104474 106744 104476
rect 106800 104474 106824 104476
rect 106880 104474 106904 104476
rect 106960 104474 106966 104476
rect 106720 104422 106722 104474
rect 106902 104422 106904 104474
rect 106658 104420 106664 104422
rect 106720 104420 106744 104422
rect 106800 104420 106824 104422
rect 106880 104420 106904 104422
rect 106960 104420 106966 104422
rect 106658 104411 106966 104420
rect 105922 103932 106230 103941
rect 105922 103930 105928 103932
rect 105984 103930 106008 103932
rect 106064 103930 106088 103932
rect 106144 103930 106168 103932
rect 106224 103930 106230 103932
rect 105984 103878 105986 103930
rect 106166 103878 106168 103930
rect 105922 103876 105928 103878
rect 105984 103876 106008 103878
rect 106064 103876 106088 103878
rect 106144 103876 106168 103878
rect 106224 103876 106230 103878
rect 105922 103867 106230 103876
rect 106658 103388 106966 103397
rect 106658 103386 106664 103388
rect 106720 103386 106744 103388
rect 106800 103386 106824 103388
rect 106880 103386 106904 103388
rect 106960 103386 106966 103388
rect 106720 103334 106722 103386
rect 106902 103334 106904 103386
rect 106658 103332 106664 103334
rect 106720 103332 106744 103334
rect 106800 103332 106824 103334
rect 106880 103332 106904 103334
rect 106960 103332 106966 103334
rect 106658 103323 106966 103332
rect 105922 102844 106230 102853
rect 105922 102842 105928 102844
rect 105984 102842 106008 102844
rect 106064 102842 106088 102844
rect 106144 102842 106168 102844
rect 106224 102842 106230 102844
rect 105984 102790 105986 102842
rect 106166 102790 106168 102842
rect 105922 102788 105928 102790
rect 105984 102788 106008 102790
rect 106064 102788 106088 102790
rect 106144 102788 106168 102790
rect 106224 102788 106230 102790
rect 105922 102779 106230 102788
rect 106658 102300 106966 102309
rect 106658 102298 106664 102300
rect 106720 102298 106744 102300
rect 106800 102298 106824 102300
rect 106880 102298 106904 102300
rect 106960 102298 106966 102300
rect 106720 102246 106722 102298
rect 106902 102246 106904 102298
rect 106658 102244 106664 102246
rect 106720 102244 106744 102246
rect 106800 102244 106824 102246
rect 106880 102244 106904 102246
rect 106960 102244 106966 102246
rect 106658 102235 106966 102244
rect 105922 101756 106230 101765
rect 105922 101754 105928 101756
rect 105984 101754 106008 101756
rect 106064 101754 106088 101756
rect 106144 101754 106168 101756
rect 106224 101754 106230 101756
rect 105984 101702 105986 101754
rect 106166 101702 106168 101754
rect 105922 101700 105928 101702
rect 105984 101700 106008 101702
rect 106064 101700 106088 101702
rect 106144 101700 106168 101702
rect 106224 101700 106230 101702
rect 105922 101691 106230 101700
rect 106658 101212 106966 101221
rect 106658 101210 106664 101212
rect 106720 101210 106744 101212
rect 106800 101210 106824 101212
rect 106880 101210 106904 101212
rect 106960 101210 106966 101212
rect 106720 101158 106722 101210
rect 106902 101158 106904 101210
rect 106658 101156 106664 101158
rect 106720 101156 106744 101158
rect 106800 101156 106824 101158
rect 106880 101156 106904 101158
rect 106960 101156 106966 101158
rect 106658 101147 106966 101156
rect 105820 100904 105872 100910
rect 105820 100846 105872 100852
rect 105636 100836 105688 100842
rect 105636 100778 105688 100784
rect 105648 96490 105676 100778
rect 105820 100768 105872 100774
rect 105820 100710 105872 100716
rect 105636 96484 105688 96490
rect 105636 96426 105688 96432
rect 105728 96416 105780 96422
rect 105728 96358 105780 96364
rect 105740 96150 105768 96358
rect 105728 96144 105780 96150
rect 105728 96086 105780 96092
rect 105084 91588 105136 91594
rect 105084 91530 105136 91536
rect 104348 77716 104400 77722
rect 104348 77658 104400 77664
rect 105096 77586 105124 91530
rect 105832 80102 105860 100710
rect 105922 100668 106230 100677
rect 105922 100666 105928 100668
rect 105984 100666 106008 100668
rect 106064 100666 106088 100668
rect 106144 100666 106168 100668
rect 106224 100666 106230 100668
rect 105984 100614 105986 100666
rect 106166 100614 106168 100666
rect 105922 100612 105928 100614
rect 105984 100612 106008 100614
rect 106064 100612 106088 100614
rect 106144 100612 106168 100614
rect 106224 100612 106230 100614
rect 105922 100603 106230 100612
rect 106658 100124 106966 100133
rect 106658 100122 106664 100124
rect 106720 100122 106744 100124
rect 106800 100122 106824 100124
rect 106880 100122 106904 100124
rect 106960 100122 106966 100124
rect 106720 100070 106722 100122
rect 106902 100070 106904 100122
rect 106658 100068 106664 100070
rect 106720 100068 106744 100070
rect 106800 100068 106824 100070
rect 106880 100068 106904 100070
rect 106960 100068 106966 100070
rect 106658 100059 106966 100068
rect 105922 99580 106230 99589
rect 105922 99578 105928 99580
rect 105984 99578 106008 99580
rect 106064 99578 106088 99580
rect 106144 99578 106168 99580
rect 106224 99578 106230 99580
rect 105984 99526 105986 99578
rect 106166 99526 106168 99578
rect 105922 99524 105928 99526
rect 105984 99524 106008 99526
rect 106064 99524 106088 99526
rect 106144 99524 106168 99526
rect 106224 99524 106230 99526
rect 105922 99515 106230 99524
rect 106658 99036 106966 99045
rect 106658 99034 106664 99036
rect 106720 99034 106744 99036
rect 106800 99034 106824 99036
rect 106880 99034 106904 99036
rect 106960 99034 106966 99036
rect 106720 98982 106722 99034
rect 106902 98982 106904 99034
rect 106658 98980 106664 98982
rect 106720 98980 106744 98982
rect 106800 98980 106824 98982
rect 106880 98980 106904 98982
rect 106960 98980 106966 98982
rect 106658 98971 106966 98980
rect 105922 98492 106230 98501
rect 105922 98490 105928 98492
rect 105984 98490 106008 98492
rect 106064 98490 106088 98492
rect 106144 98490 106168 98492
rect 106224 98490 106230 98492
rect 105984 98438 105986 98490
rect 106166 98438 106168 98490
rect 105922 98436 105928 98438
rect 105984 98436 106008 98438
rect 106064 98436 106088 98438
rect 106144 98436 106168 98438
rect 106224 98436 106230 98438
rect 105922 98427 106230 98436
rect 106658 97948 106966 97957
rect 106658 97946 106664 97948
rect 106720 97946 106744 97948
rect 106800 97946 106824 97948
rect 106880 97946 106904 97948
rect 106960 97946 106966 97948
rect 106720 97894 106722 97946
rect 106902 97894 106904 97946
rect 106658 97892 106664 97894
rect 106720 97892 106744 97894
rect 106800 97892 106824 97894
rect 106880 97892 106904 97894
rect 106960 97892 106966 97894
rect 106658 97883 106966 97892
rect 105922 97404 106230 97413
rect 105922 97402 105928 97404
rect 105984 97402 106008 97404
rect 106064 97402 106088 97404
rect 106144 97402 106168 97404
rect 106224 97402 106230 97404
rect 105984 97350 105986 97402
rect 106166 97350 106168 97402
rect 105922 97348 105928 97350
rect 105984 97348 106008 97350
rect 106064 97348 106088 97350
rect 106144 97348 106168 97350
rect 106224 97348 106230 97350
rect 105922 97339 106230 97348
rect 106658 96860 106966 96869
rect 106658 96858 106664 96860
rect 106720 96858 106744 96860
rect 106800 96858 106824 96860
rect 106880 96858 106904 96860
rect 106960 96858 106966 96860
rect 106720 96806 106722 96858
rect 106902 96806 106904 96858
rect 106658 96804 106664 96806
rect 106720 96804 106744 96806
rect 106800 96804 106824 96806
rect 106880 96804 106904 96806
rect 106960 96804 106966 96806
rect 106658 96795 106966 96804
rect 105922 96316 106230 96325
rect 105922 96314 105928 96316
rect 105984 96314 106008 96316
rect 106064 96314 106088 96316
rect 106144 96314 106168 96316
rect 106224 96314 106230 96316
rect 105984 96262 105986 96314
rect 106166 96262 106168 96314
rect 105922 96260 105928 96262
rect 105984 96260 106008 96262
rect 106064 96260 106088 96262
rect 106144 96260 106168 96262
rect 106224 96260 106230 96262
rect 105922 96251 106230 96260
rect 106658 95772 106966 95781
rect 106658 95770 106664 95772
rect 106720 95770 106744 95772
rect 106800 95770 106824 95772
rect 106880 95770 106904 95772
rect 106960 95770 106966 95772
rect 106720 95718 106722 95770
rect 106902 95718 106904 95770
rect 106658 95716 106664 95718
rect 106720 95716 106744 95718
rect 106800 95716 106824 95718
rect 106880 95716 106904 95718
rect 106960 95716 106966 95718
rect 106658 95707 106966 95716
rect 105922 95228 106230 95237
rect 105922 95226 105928 95228
rect 105984 95226 106008 95228
rect 106064 95226 106088 95228
rect 106144 95226 106168 95228
rect 106224 95226 106230 95228
rect 105984 95174 105986 95226
rect 106166 95174 106168 95226
rect 105922 95172 105928 95174
rect 105984 95172 106008 95174
rect 106064 95172 106088 95174
rect 106144 95172 106168 95174
rect 106224 95172 106230 95174
rect 105922 95163 106230 95172
rect 106658 94684 106966 94693
rect 106658 94682 106664 94684
rect 106720 94682 106744 94684
rect 106800 94682 106824 94684
rect 106880 94682 106904 94684
rect 106960 94682 106966 94684
rect 106720 94630 106722 94682
rect 106902 94630 106904 94682
rect 106658 94628 106664 94630
rect 106720 94628 106744 94630
rect 106800 94628 106824 94630
rect 106880 94628 106904 94630
rect 106960 94628 106966 94630
rect 106658 94619 106966 94628
rect 105922 94140 106230 94149
rect 105922 94138 105928 94140
rect 105984 94138 106008 94140
rect 106064 94138 106088 94140
rect 106144 94138 106168 94140
rect 106224 94138 106230 94140
rect 105984 94086 105986 94138
rect 106166 94086 106168 94138
rect 105922 94084 105928 94086
rect 105984 94084 106008 94086
rect 106064 94084 106088 94086
rect 106144 94084 106168 94086
rect 106224 94084 106230 94086
rect 105922 94075 106230 94084
rect 106658 93596 106966 93605
rect 106658 93594 106664 93596
rect 106720 93594 106744 93596
rect 106800 93594 106824 93596
rect 106880 93594 106904 93596
rect 106960 93594 106966 93596
rect 106720 93542 106722 93594
rect 106902 93542 106904 93594
rect 106658 93540 106664 93542
rect 106720 93540 106744 93542
rect 106800 93540 106824 93542
rect 106880 93540 106904 93542
rect 106960 93540 106966 93542
rect 106658 93531 106966 93540
rect 105922 93052 106230 93061
rect 105922 93050 105928 93052
rect 105984 93050 106008 93052
rect 106064 93050 106088 93052
rect 106144 93050 106168 93052
rect 106224 93050 106230 93052
rect 105984 92998 105986 93050
rect 106166 92998 106168 93050
rect 105922 92996 105928 92998
rect 105984 92996 106008 92998
rect 106064 92996 106088 92998
rect 106144 92996 106168 92998
rect 106224 92996 106230 92998
rect 105922 92987 106230 92996
rect 106658 92508 106966 92517
rect 106658 92506 106664 92508
rect 106720 92506 106744 92508
rect 106800 92506 106824 92508
rect 106880 92506 106904 92508
rect 106960 92506 106966 92508
rect 106720 92454 106722 92506
rect 106902 92454 106904 92506
rect 106658 92452 106664 92454
rect 106720 92452 106744 92454
rect 106800 92452 106824 92454
rect 106880 92452 106904 92454
rect 106960 92452 106966 92454
rect 106658 92443 106966 92452
rect 105922 91964 106230 91973
rect 105922 91962 105928 91964
rect 105984 91962 106008 91964
rect 106064 91962 106088 91964
rect 106144 91962 106168 91964
rect 106224 91962 106230 91964
rect 105984 91910 105986 91962
rect 106166 91910 106168 91962
rect 105922 91908 105928 91910
rect 105984 91908 106008 91910
rect 106064 91908 106088 91910
rect 106144 91908 106168 91910
rect 106224 91908 106230 91910
rect 105922 91899 106230 91908
rect 106658 91420 106966 91429
rect 106658 91418 106664 91420
rect 106720 91418 106744 91420
rect 106800 91418 106824 91420
rect 106880 91418 106904 91420
rect 106960 91418 106966 91420
rect 106720 91366 106722 91418
rect 106902 91366 106904 91418
rect 106658 91364 106664 91366
rect 106720 91364 106744 91366
rect 106800 91364 106824 91366
rect 106880 91364 106904 91366
rect 106960 91364 106966 91366
rect 106658 91355 106966 91364
rect 105922 90876 106230 90885
rect 105922 90874 105928 90876
rect 105984 90874 106008 90876
rect 106064 90874 106088 90876
rect 106144 90874 106168 90876
rect 106224 90874 106230 90876
rect 105984 90822 105986 90874
rect 106166 90822 106168 90874
rect 105922 90820 105928 90822
rect 105984 90820 106008 90822
rect 106064 90820 106088 90822
rect 106144 90820 106168 90822
rect 106224 90820 106230 90822
rect 105922 90811 106230 90820
rect 106658 90332 106966 90341
rect 106658 90330 106664 90332
rect 106720 90330 106744 90332
rect 106800 90330 106824 90332
rect 106880 90330 106904 90332
rect 106960 90330 106966 90332
rect 106720 90278 106722 90330
rect 106902 90278 106904 90330
rect 106658 90276 106664 90278
rect 106720 90276 106744 90278
rect 106800 90276 106824 90278
rect 106880 90276 106904 90278
rect 106960 90276 106966 90278
rect 106658 90267 106966 90276
rect 105922 89788 106230 89797
rect 105922 89786 105928 89788
rect 105984 89786 106008 89788
rect 106064 89786 106088 89788
rect 106144 89786 106168 89788
rect 106224 89786 106230 89788
rect 105984 89734 105986 89786
rect 106166 89734 106168 89786
rect 105922 89732 105928 89734
rect 105984 89732 106008 89734
rect 106064 89732 106088 89734
rect 106144 89732 106168 89734
rect 106224 89732 106230 89734
rect 105922 89723 106230 89732
rect 106658 89244 106966 89253
rect 106658 89242 106664 89244
rect 106720 89242 106744 89244
rect 106800 89242 106824 89244
rect 106880 89242 106904 89244
rect 106960 89242 106966 89244
rect 106720 89190 106722 89242
rect 106902 89190 106904 89242
rect 106658 89188 106664 89190
rect 106720 89188 106744 89190
rect 106800 89188 106824 89190
rect 106880 89188 106904 89190
rect 106960 89188 106966 89190
rect 106658 89179 106966 89188
rect 105922 88700 106230 88709
rect 105922 88698 105928 88700
rect 105984 88698 106008 88700
rect 106064 88698 106088 88700
rect 106144 88698 106168 88700
rect 106224 88698 106230 88700
rect 105984 88646 105986 88698
rect 106166 88646 106168 88698
rect 105922 88644 105928 88646
rect 105984 88644 106008 88646
rect 106064 88644 106088 88646
rect 106144 88644 106168 88646
rect 106224 88644 106230 88646
rect 105922 88635 106230 88644
rect 106658 88156 106966 88165
rect 106658 88154 106664 88156
rect 106720 88154 106744 88156
rect 106800 88154 106824 88156
rect 106880 88154 106904 88156
rect 106960 88154 106966 88156
rect 106720 88102 106722 88154
rect 106902 88102 106904 88154
rect 106658 88100 106664 88102
rect 106720 88100 106744 88102
rect 106800 88100 106824 88102
rect 106880 88100 106904 88102
rect 106960 88100 106966 88102
rect 106658 88091 106966 88100
rect 105922 87612 106230 87621
rect 105922 87610 105928 87612
rect 105984 87610 106008 87612
rect 106064 87610 106088 87612
rect 106144 87610 106168 87612
rect 106224 87610 106230 87612
rect 105984 87558 105986 87610
rect 106166 87558 106168 87610
rect 105922 87556 105928 87558
rect 105984 87556 106008 87558
rect 106064 87556 106088 87558
rect 106144 87556 106168 87558
rect 106224 87556 106230 87558
rect 105922 87547 106230 87556
rect 106658 87068 106966 87077
rect 106658 87066 106664 87068
rect 106720 87066 106744 87068
rect 106800 87066 106824 87068
rect 106880 87066 106904 87068
rect 106960 87066 106966 87068
rect 106720 87014 106722 87066
rect 106902 87014 106904 87066
rect 106658 87012 106664 87014
rect 106720 87012 106744 87014
rect 106800 87012 106824 87014
rect 106880 87012 106904 87014
rect 106960 87012 106966 87014
rect 106658 87003 106966 87012
rect 105922 86524 106230 86533
rect 105922 86522 105928 86524
rect 105984 86522 106008 86524
rect 106064 86522 106088 86524
rect 106144 86522 106168 86524
rect 106224 86522 106230 86524
rect 105984 86470 105986 86522
rect 106166 86470 106168 86522
rect 105922 86468 105928 86470
rect 105984 86468 106008 86470
rect 106064 86468 106088 86470
rect 106144 86468 106168 86470
rect 106224 86468 106230 86470
rect 105922 86459 106230 86468
rect 106658 85980 106966 85989
rect 106658 85978 106664 85980
rect 106720 85978 106744 85980
rect 106800 85978 106824 85980
rect 106880 85978 106904 85980
rect 106960 85978 106966 85980
rect 106720 85926 106722 85978
rect 106902 85926 106904 85978
rect 106658 85924 106664 85926
rect 106720 85924 106744 85926
rect 106800 85924 106824 85926
rect 106880 85924 106904 85926
rect 106960 85924 106966 85926
rect 106658 85915 106966 85924
rect 105922 85436 106230 85445
rect 105922 85434 105928 85436
rect 105984 85434 106008 85436
rect 106064 85434 106088 85436
rect 106144 85434 106168 85436
rect 106224 85434 106230 85436
rect 105984 85382 105986 85434
rect 106166 85382 106168 85434
rect 105922 85380 105928 85382
rect 105984 85380 106008 85382
rect 106064 85380 106088 85382
rect 106144 85380 106168 85382
rect 106224 85380 106230 85382
rect 105922 85371 106230 85380
rect 106658 84892 106966 84901
rect 106658 84890 106664 84892
rect 106720 84890 106744 84892
rect 106800 84890 106824 84892
rect 106880 84890 106904 84892
rect 106960 84890 106966 84892
rect 106720 84838 106722 84890
rect 106902 84838 106904 84890
rect 106658 84836 106664 84838
rect 106720 84836 106744 84838
rect 106800 84836 106824 84838
rect 106880 84836 106904 84838
rect 106960 84836 106966 84838
rect 106658 84827 106966 84836
rect 105922 84348 106230 84357
rect 105922 84346 105928 84348
rect 105984 84346 106008 84348
rect 106064 84346 106088 84348
rect 106144 84346 106168 84348
rect 106224 84346 106230 84348
rect 105984 84294 105986 84346
rect 106166 84294 106168 84346
rect 105922 84292 105928 84294
rect 105984 84292 106008 84294
rect 106064 84292 106088 84294
rect 106144 84292 106168 84294
rect 106224 84292 106230 84294
rect 105922 84283 106230 84292
rect 106658 83804 106966 83813
rect 106658 83802 106664 83804
rect 106720 83802 106744 83804
rect 106800 83802 106824 83804
rect 106880 83802 106904 83804
rect 106960 83802 106966 83804
rect 106720 83750 106722 83802
rect 106902 83750 106904 83802
rect 106658 83748 106664 83750
rect 106720 83748 106744 83750
rect 106800 83748 106824 83750
rect 106880 83748 106904 83750
rect 106960 83748 106966 83750
rect 106658 83739 106966 83748
rect 105922 83260 106230 83269
rect 105922 83258 105928 83260
rect 105984 83258 106008 83260
rect 106064 83258 106088 83260
rect 106144 83258 106168 83260
rect 106224 83258 106230 83260
rect 105984 83206 105986 83258
rect 106166 83206 106168 83258
rect 105922 83204 105928 83206
rect 105984 83204 106008 83206
rect 106064 83204 106088 83206
rect 106144 83204 106168 83206
rect 106224 83204 106230 83206
rect 105922 83195 106230 83204
rect 106658 82716 106966 82725
rect 106658 82714 106664 82716
rect 106720 82714 106744 82716
rect 106800 82714 106824 82716
rect 106880 82714 106904 82716
rect 106960 82714 106966 82716
rect 106720 82662 106722 82714
rect 106902 82662 106904 82714
rect 106658 82660 106664 82662
rect 106720 82660 106744 82662
rect 106800 82660 106824 82662
rect 106880 82660 106904 82662
rect 106960 82660 106966 82662
rect 106658 82651 106966 82660
rect 105922 82172 106230 82181
rect 105922 82170 105928 82172
rect 105984 82170 106008 82172
rect 106064 82170 106088 82172
rect 106144 82170 106168 82172
rect 106224 82170 106230 82172
rect 105984 82118 105986 82170
rect 106166 82118 106168 82170
rect 105922 82116 105928 82118
rect 105984 82116 106008 82118
rect 106064 82116 106088 82118
rect 106144 82116 106168 82118
rect 106224 82116 106230 82118
rect 105922 82107 106230 82116
rect 106658 81628 106966 81637
rect 106658 81626 106664 81628
rect 106720 81626 106744 81628
rect 106800 81626 106824 81628
rect 106880 81626 106904 81628
rect 106960 81626 106966 81628
rect 106720 81574 106722 81626
rect 106902 81574 106904 81626
rect 106658 81572 106664 81574
rect 106720 81572 106744 81574
rect 106800 81572 106824 81574
rect 106880 81572 106904 81574
rect 106960 81572 106966 81574
rect 106658 81563 106966 81572
rect 105922 81084 106230 81093
rect 105922 81082 105928 81084
rect 105984 81082 106008 81084
rect 106064 81082 106088 81084
rect 106144 81082 106168 81084
rect 106224 81082 106230 81084
rect 105984 81030 105986 81082
rect 106166 81030 106168 81082
rect 105922 81028 105928 81030
rect 105984 81028 106008 81030
rect 106064 81028 106088 81030
rect 106144 81028 106168 81030
rect 106224 81028 106230 81030
rect 105922 81019 106230 81028
rect 107752 80776 107804 80782
rect 107752 80718 107804 80724
rect 108488 80776 108540 80782
rect 108488 80718 108540 80724
rect 106658 80540 106966 80549
rect 106658 80538 106664 80540
rect 106720 80538 106744 80540
rect 106800 80538 106824 80540
rect 106880 80538 106904 80540
rect 106960 80538 106966 80540
rect 106720 80486 106722 80538
rect 106902 80486 106904 80538
rect 106658 80484 106664 80486
rect 106720 80484 106744 80486
rect 106800 80484 106824 80486
rect 106880 80484 106904 80486
rect 106960 80484 106966 80486
rect 106658 80475 106966 80484
rect 105820 80096 105872 80102
rect 105820 80038 105872 80044
rect 105922 79996 106230 80005
rect 105922 79994 105928 79996
rect 105984 79994 106008 79996
rect 106064 79994 106088 79996
rect 106144 79994 106168 79996
rect 106224 79994 106230 79996
rect 105984 79942 105986 79994
rect 106166 79942 106168 79994
rect 105922 79940 105928 79942
rect 105984 79940 106008 79942
rect 106064 79940 106088 79942
rect 106144 79940 106168 79942
rect 106224 79940 106230 79942
rect 105922 79931 106230 79940
rect 106658 79452 106966 79461
rect 106658 79450 106664 79452
rect 106720 79450 106744 79452
rect 106800 79450 106824 79452
rect 106880 79450 106904 79452
rect 106960 79450 106966 79452
rect 106720 79398 106722 79450
rect 106902 79398 106904 79450
rect 106658 79396 106664 79398
rect 106720 79396 106744 79398
rect 106800 79396 106824 79398
rect 106880 79396 106904 79398
rect 106960 79396 106966 79398
rect 106658 79387 106966 79396
rect 105922 78908 106230 78917
rect 105922 78906 105928 78908
rect 105984 78906 106008 78908
rect 106064 78906 106088 78908
rect 106144 78906 106168 78908
rect 106224 78906 106230 78908
rect 105984 78854 105986 78906
rect 106166 78854 106168 78906
rect 105922 78852 105928 78854
rect 105984 78852 106008 78854
rect 106064 78852 106088 78854
rect 106144 78852 106168 78854
rect 106224 78852 106230 78854
rect 105922 78843 106230 78852
rect 107660 78600 107712 78606
rect 107660 78542 107712 78548
rect 106658 78364 106966 78373
rect 106658 78362 106664 78364
rect 106720 78362 106744 78364
rect 106800 78362 106824 78364
rect 106880 78362 106904 78364
rect 106960 78362 106966 78364
rect 106720 78310 106722 78362
rect 106902 78310 106904 78362
rect 106658 78308 106664 78310
rect 106720 78308 106744 78310
rect 106800 78308 106824 78310
rect 106880 78308 106904 78310
rect 106960 78308 106966 78310
rect 106658 78299 106966 78308
rect 105922 77820 106230 77829
rect 105922 77818 105928 77820
rect 105984 77818 106008 77820
rect 106064 77818 106088 77820
rect 106144 77818 106168 77820
rect 106224 77818 106230 77820
rect 105984 77766 105986 77818
rect 106166 77766 106168 77818
rect 105922 77764 105928 77766
rect 105984 77764 106008 77766
rect 106064 77764 106088 77766
rect 106144 77764 106168 77766
rect 106224 77764 106230 77766
rect 105922 77755 106230 77764
rect 105084 77580 105136 77586
rect 105084 77522 105136 77528
rect 106658 77276 106966 77285
rect 106658 77274 106664 77276
rect 106720 77274 106744 77276
rect 106800 77274 106824 77276
rect 106880 77274 106904 77276
rect 106960 77274 106966 77276
rect 106720 77222 106722 77274
rect 106902 77222 106904 77274
rect 106658 77220 106664 77222
rect 106720 77220 106744 77222
rect 106800 77220 106824 77222
rect 106880 77220 106904 77222
rect 106960 77220 106966 77222
rect 106658 77211 106966 77220
rect 107672 76906 107700 78542
rect 107660 76900 107712 76906
rect 107660 76842 107712 76848
rect 101680 75880 101732 75886
rect 101680 75822 101732 75828
rect 104072 75880 104124 75886
rect 104072 75822 104124 75828
rect 101692 75546 101720 75822
rect 101680 75540 101732 75546
rect 101680 75482 101732 75488
rect 104164 75540 104216 75546
rect 104164 75482 104216 75488
rect 104808 75540 104860 75546
rect 104808 75482 104860 75488
rect 103520 75472 103572 75478
rect 101968 75410 102088 75426
rect 103520 75414 103572 75420
rect 103980 75472 104032 75478
rect 103980 75414 104032 75420
rect 101404 75404 101456 75410
rect 101404 75346 101456 75352
rect 101956 75404 102088 75410
rect 102008 75398 102088 75404
rect 101956 75346 102008 75352
rect 101220 75200 101272 75206
rect 101220 75142 101272 75148
rect 101232 75002 101260 75142
rect 101220 74996 101272 75002
rect 101220 74938 101272 74944
rect 101416 74866 101444 75346
rect 101956 75268 102008 75274
rect 101956 75210 102008 75216
rect 101864 74996 101916 75002
rect 101864 74938 101916 74944
rect 100208 74860 100260 74866
rect 100208 74802 100260 74808
rect 100300 74860 100352 74866
rect 100300 74802 100352 74808
rect 100484 74860 100536 74866
rect 100484 74802 100536 74808
rect 100668 74860 100720 74866
rect 100668 74802 100720 74808
rect 101128 74860 101180 74866
rect 101128 74802 101180 74808
rect 101404 74860 101456 74866
rect 101404 74802 101456 74808
rect 100312 74746 100340 74802
rect 100680 74746 100708 74802
rect 100208 74724 100260 74730
rect 100208 74666 100260 74672
rect 100312 74718 100708 74746
rect 100220 74338 100248 74666
rect 100312 74662 100340 74718
rect 100300 74656 100352 74662
rect 100300 74598 100352 74604
rect 100760 74656 100812 74662
rect 100760 74598 100812 74604
rect 100390 74488 100446 74497
rect 100390 74423 100446 74432
rect 100404 74390 100432 74423
rect 100392 74384 100444 74390
rect 100220 74310 100340 74338
rect 100392 74326 100444 74332
rect 100772 74322 100800 74598
rect 101876 74322 101904 74938
rect 101968 74866 101996 75210
rect 102060 74866 102088 75398
rect 103152 75404 103204 75410
rect 103152 75346 103204 75352
rect 103336 75404 103388 75410
rect 103336 75346 103388 75352
rect 102968 75336 103020 75342
rect 102968 75278 103020 75284
rect 102876 75268 102928 75274
rect 102876 75210 102928 75216
rect 101956 74860 102008 74866
rect 101956 74802 102008 74808
rect 102048 74860 102100 74866
rect 102048 74802 102100 74808
rect 102508 74860 102560 74866
rect 102508 74802 102560 74808
rect 101968 74458 101996 74802
rect 101956 74452 102008 74458
rect 101956 74394 102008 74400
rect 102060 74390 102088 74802
rect 102048 74384 102100 74390
rect 102048 74326 102100 74332
rect 102140 74384 102192 74390
rect 102140 74326 102192 74332
rect 100208 74248 100260 74254
rect 100206 74216 100208 74225
rect 100260 74216 100262 74225
rect 100206 74151 100262 74160
rect 100116 73568 100168 73574
rect 100116 73510 100168 73516
rect 100116 73296 100168 73302
rect 100116 73238 100168 73244
rect 100024 72820 100076 72826
rect 100024 72762 100076 72768
rect 100024 72616 100076 72622
rect 100024 72558 100076 72564
rect 100036 72078 100064 72558
rect 100024 72072 100076 72078
rect 100024 72014 100076 72020
rect 99748 71596 99800 71602
rect 99748 71538 99800 71544
rect 99840 71596 99892 71602
rect 99840 71538 99892 71544
rect 99104 71460 99156 71466
rect 99104 71402 99156 71408
rect 98920 71392 98972 71398
rect 98920 71334 98972 71340
rect 99380 71392 99432 71398
rect 99380 71334 99432 71340
rect 98828 71188 98880 71194
rect 98828 71130 98880 71136
rect 98552 71120 98604 71126
rect 98552 71062 98604 71068
rect 98644 70984 98696 70990
rect 98644 70926 98696 70932
rect 98736 70984 98788 70990
rect 98840 70961 98868 71130
rect 98736 70926 98788 70932
rect 98826 70952 98882 70961
rect 98460 70848 98512 70854
rect 98460 70790 98512 70796
rect 98368 70576 98420 70582
rect 98368 70518 98420 70524
rect 98472 70496 98500 70790
rect 98552 70508 98604 70514
rect 98472 70468 98552 70496
rect 98552 70450 98604 70456
rect 98092 70372 98144 70378
rect 98092 70314 98144 70320
rect 98196 70366 98316 70394
rect 97908 70032 97960 70038
rect 97908 69974 97960 69980
rect 97538 69935 97594 69944
rect 97816 69964 97868 69970
rect 97552 69902 97580 69935
rect 97816 69906 97868 69912
rect 97540 69896 97592 69902
rect 97540 69838 97592 69844
rect 97448 69828 97500 69834
rect 97448 69770 97500 69776
rect 96804 69760 96856 69766
rect 96804 69702 96856 69708
rect 96374 69116 96682 69125
rect 96374 69114 96380 69116
rect 96436 69114 96460 69116
rect 96516 69114 96540 69116
rect 96596 69114 96620 69116
rect 96676 69114 96682 69116
rect 96436 69062 96438 69114
rect 96618 69062 96620 69114
rect 96374 69060 96380 69062
rect 96436 69060 96460 69062
rect 96516 69060 96540 69062
rect 96596 69060 96620 69062
rect 96676 69060 96682 69062
rect 96374 69051 96682 69060
rect 96160 68876 96212 68882
rect 96160 68818 96212 68824
rect 96068 68808 96120 68814
rect 96068 68750 96120 68756
rect 96080 68474 96108 68750
rect 96068 68468 96120 68474
rect 96068 68410 96120 68416
rect 96080 68134 96108 68410
rect 96172 68338 96200 68818
rect 96160 68332 96212 68338
rect 96160 68274 96212 68280
rect 96252 68332 96304 68338
rect 96252 68274 96304 68280
rect 96068 68128 96120 68134
rect 96068 68070 96120 68076
rect 96264 67726 96292 68274
rect 96712 68128 96764 68134
rect 96712 68070 96764 68076
rect 96374 68028 96682 68037
rect 96374 68026 96380 68028
rect 96436 68026 96460 68028
rect 96516 68026 96540 68028
rect 96596 68026 96620 68028
rect 96676 68026 96682 68028
rect 96436 67974 96438 68026
rect 96618 67974 96620 68026
rect 96374 67972 96380 67974
rect 96436 67972 96460 67974
rect 96516 67972 96540 67974
rect 96596 67972 96620 67974
rect 96676 67972 96682 67974
rect 96374 67963 96682 67972
rect 96252 67720 96304 67726
rect 96252 67662 96304 67668
rect 95976 67244 96028 67250
rect 95976 67186 96028 67192
rect 96160 67040 96212 67046
rect 96160 66982 96212 66988
rect 95976 66836 96028 66842
rect 95976 66778 96028 66784
rect 95884 66496 95936 66502
rect 95884 66438 95936 66444
rect 95424 66292 95476 66298
rect 95424 66234 95476 66240
rect 95608 66292 95660 66298
rect 95608 66234 95660 66240
rect 95792 66292 95844 66298
rect 95792 66234 95844 66240
rect 95332 66156 95384 66162
rect 95332 66098 95384 66104
rect 95804 65958 95832 66234
rect 95896 66230 95924 66438
rect 95884 66224 95936 66230
rect 95884 66166 95936 66172
rect 95884 66020 95936 66026
rect 95884 65962 95936 65968
rect 94964 65952 95016 65958
rect 94964 65894 95016 65900
rect 95792 65952 95844 65958
rect 95792 65894 95844 65900
rect 94872 65680 94924 65686
rect 94872 65622 94924 65628
rect 95896 64161 95924 65962
rect 95988 65958 96016 66778
rect 96172 66706 96200 66982
rect 96374 66940 96682 66949
rect 96374 66938 96380 66940
rect 96436 66938 96460 66940
rect 96516 66938 96540 66940
rect 96596 66938 96620 66940
rect 96676 66938 96682 66940
rect 96436 66886 96438 66938
rect 96618 66886 96620 66938
rect 96374 66884 96380 66886
rect 96436 66884 96460 66886
rect 96516 66884 96540 66886
rect 96596 66884 96620 66886
rect 96676 66884 96682 66886
rect 96374 66875 96682 66884
rect 96068 66700 96120 66706
rect 96068 66642 96120 66648
rect 96160 66700 96212 66706
rect 96160 66642 96212 66648
rect 96080 66162 96108 66642
rect 96724 66230 96752 68070
rect 96816 67386 96844 69702
rect 97034 69660 97342 69669
rect 97034 69658 97040 69660
rect 97096 69658 97120 69660
rect 97176 69658 97200 69660
rect 97256 69658 97280 69660
rect 97336 69658 97342 69660
rect 97096 69606 97098 69658
rect 97278 69606 97280 69658
rect 97034 69604 97040 69606
rect 97096 69604 97120 69606
rect 97176 69604 97200 69606
rect 97256 69604 97280 69606
rect 97336 69604 97342 69606
rect 97034 69595 97342 69604
rect 97448 68808 97500 68814
rect 97448 68750 97500 68756
rect 96896 68672 96948 68678
rect 96896 68614 96948 68620
rect 96804 67380 96856 67386
rect 96804 67322 96856 67328
rect 96908 67182 96936 68614
rect 97034 68572 97342 68581
rect 97034 68570 97040 68572
rect 97096 68570 97120 68572
rect 97176 68570 97200 68572
rect 97256 68570 97280 68572
rect 97336 68570 97342 68572
rect 97096 68518 97098 68570
rect 97278 68518 97280 68570
rect 97034 68516 97040 68518
rect 97096 68516 97120 68518
rect 97176 68516 97200 68518
rect 97256 68516 97280 68518
rect 97336 68516 97342 68518
rect 97034 68507 97342 68516
rect 97460 68338 97488 68750
rect 97448 68332 97500 68338
rect 97448 68274 97500 68280
rect 97552 67697 97580 69838
rect 97828 69562 97856 69906
rect 98196 69834 98224 70366
rect 98656 70038 98684 70926
rect 98644 70032 98696 70038
rect 98644 69974 98696 69980
rect 98184 69828 98236 69834
rect 98184 69770 98236 69776
rect 97816 69556 97868 69562
rect 97816 69498 97868 69504
rect 98000 68740 98052 68746
rect 98000 68682 98052 68688
rect 97908 68672 97960 68678
rect 97908 68614 97960 68620
rect 97632 68332 97684 68338
rect 97632 68274 97684 68280
rect 97538 67688 97594 67697
rect 97538 67623 97594 67632
rect 97034 67484 97342 67493
rect 97034 67482 97040 67484
rect 97096 67482 97120 67484
rect 97176 67482 97200 67484
rect 97256 67482 97280 67484
rect 97336 67482 97342 67484
rect 97096 67430 97098 67482
rect 97278 67430 97280 67482
rect 97034 67428 97040 67430
rect 97096 67428 97120 67430
rect 97176 67428 97200 67430
rect 97256 67428 97280 67430
rect 97336 67428 97342 67430
rect 97034 67419 97342 67428
rect 96896 67176 96948 67182
rect 96896 67118 96948 67124
rect 96908 67046 96936 67118
rect 96896 67040 96948 67046
rect 96896 66982 96948 66988
rect 97080 67040 97132 67046
rect 97080 66982 97132 66988
rect 96712 66224 96764 66230
rect 96712 66166 96764 66172
rect 96068 66156 96120 66162
rect 96068 66098 96120 66104
rect 96908 66026 96936 66982
rect 97092 66638 97120 66982
rect 97448 66700 97500 66706
rect 97448 66642 97500 66648
rect 97080 66632 97132 66638
rect 97080 66574 97132 66580
rect 97034 66396 97342 66405
rect 97034 66394 97040 66396
rect 97096 66394 97120 66396
rect 97176 66394 97200 66396
rect 97256 66394 97280 66396
rect 97336 66394 97342 66396
rect 97096 66342 97098 66394
rect 97278 66342 97280 66394
rect 97034 66340 97040 66342
rect 97096 66340 97120 66342
rect 97176 66340 97200 66342
rect 97256 66340 97280 66342
rect 97336 66340 97342 66342
rect 97034 66331 97342 66340
rect 97460 66298 97488 66642
rect 97448 66292 97500 66298
rect 97448 66234 97500 66240
rect 97552 66162 97580 67623
rect 97644 66774 97672 68274
rect 97920 68270 97948 68614
rect 98012 68406 98040 68682
rect 98196 68474 98224 69770
rect 98748 69426 98776 70926
rect 98826 70887 98882 70896
rect 98276 69420 98328 69426
rect 98276 69362 98328 69368
rect 98736 69420 98788 69426
rect 98736 69362 98788 69368
rect 98288 69018 98316 69362
rect 98276 69012 98328 69018
rect 98276 68954 98328 68960
rect 98748 68746 98776 69362
rect 98736 68740 98788 68746
rect 98736 68682 98788 68688
rect 98184 68468 98236 68474
rect 98184 68410 98236 68416
rect 98000 68400 98052 68406
rect 98000 68342 98052 68348
rect 98552 68332 98604 68338
rect 98552 68274 98604 68280
rect 97908 68264 97960 68270
rect 97908 68206 97960 68212
rect 97920 67794 97948 68206
rect 98564 67794 98592 68274
rect 98736 67924 98788 67930
rect 98736 67866 98788 67872
rect 97908 67788 97960 67794
rect 97908 67730 97960 67736
rect 98552 67788 98604 67794
rect 98552 67730 98604 67736
rect 97632 66768 97684 66774
rect 97632 66710 97684 66716
rect 97632 66564 97684 66570
rect 97632 66506 97684 66512
rect 97644 66298 97672 66506
rect 97632 66292 97684 66298
rect 97632 66234 97684 66240
rect 97540 66156 97592 66162
rect 97540 66098 97592 66104
rect 97920 66094 97948 67730
rect 98276 67652 98328 67658
rect 98276 67594 98328 67600
rect 98288 66638 98316 67594
rect 98564 66706 98592 67730
rect 98552 66700 98604 66706
rect 98552 66642 98604 66648
rect 98276 66632 98328 66638
rect 98276 66574 98328 66580
rect 98564 66162 98592 66642
rect 98748 66638 98776 67866
rect 98840 67862 98868 70887
rect 98932 70854 98960 71334
rect 99392 71194 99420 71334
rect 99380 71188 99432 71194
rect 99380 71130 99432 71136
rect 99656 71052 99708 71058
rect 99656 70994 99708 71000
rect 99472 70984 99524 70990
rect 99472 70926 99524 70932
rect 98920 70848 98972 70854
rect 98920 70790 98972 70796
rect 99484 70650 99512 70926
rect 99472 70644 99524 70650
rect 99472 70586 99524 70592
rect 99668 70582 99696 70994
rect 99656 70576 99708 70582
rect 99656 70518 99708 70524
rect 99380 70508 99432 70514
rect 99380 70450 99432 70456
rect 99196 70440 99248 70446
rect 99196 70382 99248 70388
rect 99208 70106 99236 70382
rect 99392 70106 99420 70450
rect 99748 70304 99800 70310
rect 99748 70246 99800 70252
rect 99196 70100 99248 70106
rect 99196 70042 99248 70048
rect 99380 70100 99432 70106
rect 99380 70042 99432 70048
rect 99760 69902 99788 70246
rect 99852 70106 99880 71538
rect 100036 71194 100064 72014
rect 100024 71188 100076 71194
rect 100024 71130 100076 71136
rect 100024 70984 100076 70990
rect 100128 70972 100156 73238
rect 100220 73166 100248 74151
rect 100312 73914 100340 74310
rect 100760 74316 100812 74322
rect 100760 74258 100812 74264
rect 101864 74316 101916 74322
rect 101864 74258 101916 74264
rect 100576 74248 100628 74254
rect 100574 74216 100576 74225
rect 100628 74216 100630 74225
rect 100574 74151 100630 74160
rect 100300 73908 100352 73914
rect 100300 73850 100352 73856
rect 100312 73710 100340 73850
rect 100588 73846 100616 74151
rect 100576 73840 100628 73846
rect 100576 73782 100628 73788
rect 100772 73778 100800 74258
rect 101312 74248 101364 74254
rect 101312 74190 101364 74196
rect 101680 74248 101732 74254
rect 101680 74190 101732 74196
rect 101128 73840 101180 73846
rect 101128 73782 101180 73788
rect 100484 73772 100536 73778
rect 100484 73714 100536 73720
rect 100760 73772 100812 73778
rect 100760 73714 100812 73720
rect 100300 73704 100352 73710
rect 100300 73646 100352 73652
rect 100392 73704 100444 73710
rect 100392 73646 100444 73652
rect 100300 73568 100352 73574
rect 100300 73510 100352 73516
rect 100312 73370 100340 73510
rect 100404 73370 100432 73646
rect 100300 73364 100352 73370
rect 100300 73306 100352 73312
rect 100392 73364 100444 73370
rect 100392 73306 100444 73312
rect 100208 73160 100260 73166
rect 100208 73102 100260 73108
rect 100496 73030 100524 73714
rect 100668 73160 100720 73166
rect 100668 73102 100720 73108
rect 100484 73024 100536 73030
rect 100484 72966 100536 72972
rect 100680 72690 100708 73102
rect 100852 72820 100904 72826
rect 100852 72762 100904 72768
rect 100392 72684 100444 72690
rect 100392 72626 100444 72632
rect 100668 72684 100720 72690
rect 100668 72626 100720 72632
rect 100300 72072 100352 72078
rect 100300 72014 100352 72020
rect 100312 71738 100340 72014
rect 100404 71738 100432 72626
rect 100576 71936 100628 71942
rect 100576 71878 100628 71884
rect 100300 71732 100352 71738
rect 100300 71674 100352 71680
rect 100392 71732 100444 71738
rect 100392 71674 100444 71680
rect 100300 71528 100352 71534
rect 100300 71470 100352 71476
rect 100312 71194 100340 71470
rect 100588 71466 100616 71878
rect 100576 71460 100628 71466
rect 100576 71402 100628 71408
rect 100300 71188 100352 71194
rect 100300 71130 100352 71136
rect 100076 70944 100156 70972
rect 100024 70926 100076 70932
rect 100036 70854 100064 70926
rect 100024 70848 100076 70854
rect 100024 70790 100076 70796
rect 99840 70100 99892 70106
rect 99840 70042 99892 70048
rect 100036 70009 100064 70790
rect 100208 70508 100260 70514
rect 100208 70450 100260 70456
rect 100220 70106 100248 70450
rect 100208 70100 100260 70106
rect 100208 70042 100260 70048
rect 100022 70000 100078 70009
rect 100022 69935 100078 69944
rect 99012 69896 99064 69902
rect 99472 69896 99524 69902
rect 99064 69856 99144 69884
rect 99012 69838 99064 69844
rect 99116 69426 99144 69856
rect 99472 69838 99524 69844
rect 99748 69896 99800 69902
rect 99748 69838 99800 69844
rect 100484 69896 100536 69902
rect 100588 69884 100616 71402
rect 100680 71398 100708 72626
rect 100864 72146 100892 72762
rect 101140 72690 101168 73782
rect 101324 73642 101352 74190
rect 101588 74112 101640 74118
rect 101588 74054 101640 74060
rect 101600 73846 101628 74054
rect 101588 73840 101640 73846
rect 101588 73782 101640 73788
rect 101312 73636 101364 73642
rect 101312 73578 101364 73584
rect 101220 73092 101272 73098
rect 101220 73034 101272 73040
rect 101232 72826 101260 73034
rect 101220 72820 101272 72826
rect 101220 72762 101272 72768
rect 101128 72684 101180 72690
rect 101128 72626 101180 72632
rect 101324 72554 101352 73578
rect 101588 73296 101640 73302
rect 101588 73238 101640 73244
rect 101496 73024 101548 73030
rect 101496 72966 101548 72972
rect 101508 72622 101536 72966
rect 101600 72690 101628 73238
rect 101588 72684 101640 72690
rect 101588 72626 101640 72632
rect 101496 72616 101548 72622
rect 101496 72558 101548 72564
rect 101312 72548 101364 72554
rect 101312 72490 101364 72496
rect 100852 72140 100904 72146
rect 100852 72082 100904 72088
rect 100864 71602 100892 72082
rect 101220 72072 101272 72078
rect 101220 72014 101272 72020
rect 100852 71596 100904 71602
rect 100852 71538 100904 71544
rect 100668 71392 100720 71398
rect 100668 71334 100720 71340
rect 101036 70984 101088 70990
rect 101034 70952 101036 70961
rect 101088 70952 101090 70961
rect 101034 70887 101090 70896
rect 100536 69856 100616 69884
rect 100484 69838 100536 69844
rect 99484 69562 99512 69838
rect 99656 69760 99708 69766
rect 99656 69702 99708 69708
rect 99472 69556 99524 69562
rect 99472 69498 99524 69504
rect 98920 69420 98972 69426
rect 98920 69362 98972 69368
rect 99104 69420 99156 69426
rect 99380 69420 99432 69426
rect 99156 69380 99380 69408
rect 99104 69362 99156 69368
rect 99380 69362 99432 69368
rect 98932 69222 98960 69362
rect 98920 69216 98972 69222
rect 98920 69158 98972 69164
rect 98828 67856 98880 67862
rect 98828 67798 98880 67804
rect 98932 67658 98960 69158
rect 99196 68740 99248 68746
rect 99196 68682 99248 68688
rect 99208 67862 99236 68682
rect 99288 68332 99340 68338
rect 99288 68274 99340 68280
rect 99300 67930 99328 68274
rect 99484 68270 99512 69498
rect 99564 69488 99616 69494
rect 99564 69430 99616 69436
rect 99576 69204 99604 69430
rect 99668 69426 99696 69702
rect 99760 69426 99788 69838
rect 100024 69760 100076 69766
rect 100024 69702 100076 69708
rect 100116 69760 100168 69766
rect 100116 69702 100168 69708
rect 99656 69420 99708 69426
rect 99656 69362 99708 69368
rect 99748 69420 99800 69426
rect 99748 69362 99800 69368
rect 99656 69216 99708 69222
rect 99576 69176 99656 69204
rect 99656 69158 99708 69164
rect 99668 68678 99696 69158
rect 99748 68808 99800 68814
rect 99748 68750 99800 68756
rect 99656 68672 99708 68678
rect 99656 68614 99708 68620
rect 99564 68332 99616 68338
rect 99564 68274 99616 68280
rect 99472 68264 99524 68270
rect 99472 68206 99524 68212
rect 99288 67924 99340 67930
rect 99288 67866 99340 67872
rect 99196 67856 99248 67862
rect 99196 67798 99248 67804
rect 99472 67788 99524 67794
rect 99472 67730 99524 67736
rect 99104 67720 99156 67726
rect 99104 67662 99156 67668
rect 98920 67652 98972 67658
rect 98920 67594 98972 67600
rect 99116 67386 99144 67662
rect 99104 67380 99156 67386
rect 99104 67322 99156 67328
rect 99484 66706 99512 67730
rect 99576 67386 99604 68274
rect 99760 67862 99788 68750
rect 99932 68400 99984 68406
rect 99932 68342 99984 68348
rect 99840 68332 99892 68338
rect 99840 68274 99892 68280
rect 99748 67856 99800 67862
rect 99748 67798 99800 67804
rect 99748 67652 99800 67658
rect 99748 67594 99800 67600
rect 99656 67584 99708 67590
rect 99656 67526 99708 67532
rect 99564 67380 99616 67386
rect 99564 67322 99616 67328
rect 99576 66706 99604 67322
rect 99668 67250 99696 67526
rect 99656 67244 99708 67250
rect 99656 67186 99708 67192
rect 99472 66700 99524 66706
rect 99472 66642 99524 66648
rect 99564 66700 99616 66706
rect 99564 66642 99616 66648
rect 98736 66632 98788 66638
rect 98736 66574 98788 66580
rect 99656 66632 99708 66638
rect 99656 66574 99708 66580
rect 98748 66162 98776 66574
rect 99668 66162 99696 66574
rect 98552 66156 98604 66162
rect 98552 66098 98604 66104
rect 98736 66156 98788 66162
rect 98736 66098 98788 66104
rect 99380 66156 99432 66162
rect 99380 66098 99432 66104
rect 99656 66156 99708 66162
rect 99656 66098 99708 66104
rect 97908 66088 97960 66094
rect 97908 66030 97960 66036
rect 99392 66026 99420 66098
rect 99760 66026 99788 67594
rect 99852 67318 99880 68274
rect 99840 67312 99892 67318
rect 99840 67254 99892 67260
rect 99852 66774 99880 67254
rect 99944 66842 99972 68342
rect 100036 67930 100064 69702
rect 100128 68474 100156 69702
rect 100484 69216 100536 69222
rect 100484 69158 100536 69164
rect 100300 68944 100352 68950
rect 100298 68912 100300 68921
rect 100352 68912 100354 68921
rect 100298 68847 100354 68856
rect 100300 68808 100352 68814
rect 100300 68750 100352 68756
rect 100312 68474 100340 68750
rect 100116 68468 100168 68474
rect 100116 68410 100168 68416
rect 100300 68468 100352 68474
rect 100300 68410 100352 68416
rect 100208 68332 100260 68338
rect 100128 68292 100208 68320
rect 100024 67924 100076 67930
rect 100024 67866 100076 67872
rect 100128 67810 100156 68292
rect 100208 68274 100260 68280
rect 100300 68196 100352 68202
rect 100300 68138 100352 68144
rect 100036 67782 100156 67810
rect 100036 67318 100064 67782
rect 100312 67658 100340 68138
rect 100300 67652 100352 67658
rect 100300 67594 100352 67600
rect 100024 67312 100076 67318
rect 100024 67254 100076 67260
rect 100116 67176 100168 67182
rect 100116 67118 100168 67124
rect 100128 66842 100156 67118
rect 99932 66836 99984 66842
rect 99932 66778 99984 66784
rect 100116 66836 100168 66842
rect 100116 66778 100168 66784
rect 99840 66768 99892 66774
rect 99840 66710 99892 66716
rect 99932 66496 99984 66502
rect 99932 66438 99984 66444
rect 99944 66094 99972 66438
rect 100312 66094 100340 67594
rect 100496 66706 100524 69158
rect 100588 68134 100616 69856
rect 100852 69896 100904 69902
rect 100852 69838 100904 69844
rect 100944 69896 100996 69902
rect 100944 69838 100996 69844
rect 100760 69828 100812 69834
rect 100760 69770 100812 69776
rect 100772 69426 100800 69770
rect 100864 69494 100892 69838
rect 100956 69766 100984 69838
rect 100944 69760 100996 69766
rect 100944 69702 100996 69708
rect 100956 69562 100984 69702
rect 100944 69556 100996 69562
rect 100944 69498 100996 69504
rect 100852 69488 100904 69494
rect 100852 69430 100904 69436
rect 100760 69420 100812 69426
rect 100760 69362 100812 69368
rect 100852 69352 100904 69358
rect 100852 69294 100904 69300
rect 100864 69018 100892 69294
rect 101128 69216 101180 69222
rect 101128 69158 101180 69164
rect 100852 69012 100904 69018
rect 100852 68954 100904 68960
rect 100864 68377 100892 68954
rect 101140 68814 101168 69158
rect 101232 68814 101260 72014
rect 101404 72004 101456 72010
rect 101404 71946 101456 71952
rect 101416 71738 101444 71946
rect 101404 71732 101456 71738
rect 101404 71674 101456 71680
rect 101312 70508 101364 70514
rect 101312 70450 101364 70456
rect 101324 69902 101352 70450
rect 101416 69970 101444 71674
rect 101692 71584 101720 74190
rect 101772 73772 101824 73778
rect 101772 73714 101824 73720
rect 101784 73302 101812 73714
rect 101876 73370 101904 74258
rect 101956 74112 102008 74118
rect 101956 74054 102008 74060
rect 101864 73364 101916 73370
rect 101864 73306 101916 73312
rect 101772 73296 101824 73302
rect 101772 73238 101824 73244
rect 101864 73228 101916 73234
rect 101864 73170 101916 73176
rect 101772 73024 101824 73030
rect 101772 72966 101824 72972
rect 101784 72282 101812 72966
rect 101876 72690 101904 73170
rect 101864 72684 101916 72690
rect 101864 72626 101916 72632
rect 101772 72276 101824 72282
rect 101772 72218 101824 72224
rect 101772 71596 101824 71602
rect 101692 71556 101772 71584
rect 101772 71538 101824 71544
rect 101784 70854 101812 71538
rect 101864 71120 101916 71126
rect 101864 71062 101916 71068
rect 101772 70848 101824 70854
rect 101772 70790 101824 70796
rect 101876 70446 101904 71062
rect 101968 70990 101996 74054
rect 102152 73914 102180 74326
rect 102140 73908 102192 73914
rect 102140 73850 102192 73856
rect 102520 73817 102548 74802
rect 102888 74798 102916 75210
rect 102980 74934 103008 75278
rect 103060 75200 103112 75206
rect 103060 75142 103112 75148
rect 102968 74928 103020 74934
rect 102968 74870 103020 74876
rect 102876 74792 102928 74798
rect 102876 74734 102928 74740
rect 103072 74322 103100 75142
rect 103164 74662 103192 75346
rect 103348 75274 103376 75346
rect 103336 75268 103388 75274
rect 103336 75210 103388 75216
rect 103152 74656 103204 74662
rect 103152 74598 103204 74604
rect 103060 74316 103112 74322
rect 103060 74258 103112 74264
rect 102876 74112 102928 74118
rect 102876 74054 102928 74060
rect 102888 73846 102916 74054
rect 102876 73840 102928 73846
rect 102506 73808 102562 73817
rect 102876 73782 102928 73788
rect 103072 73778 103100 74258
rect 102506 73743 102562 73752
rect 102784 73772 102836 73778
rect 102520 73098 102548 73743
rect 102784 73714 102836 73720
rect 103060 73772 103112 73778
rect 103060 73714 103112 73720
rect 102796 73234 102824 73714
rect 103164 73302 103192 74598
rect 103244 74248 103296 74254
rect 103244 74190 103296 74196
rect 103152 73296 103204 73302
rect 103152 73238 103204 73244
rect 102784 73228 102836 73234
rect 102784 73170 102836 73176
rect 102508 73092 102560 73098
rect 102508 73034 102560 73040
rect 102324 72140 102376 72146
rect 102324 72082 102376 72088
rect 102336 71942 102364 72082
rect 102520 72078 102548 73034
rect 102796 72758 102824 73170
rect 103256 73166 103284 74190
rect 103348 73370 103376 75210
rect 103428 74860 103480 74866
rect 103428 74802 103480 74808
rect 103440 74662 103468 74802
rect 103428 74656 103480 74662
rect 103428 74598 103480 74604
rect 103428 74452 103480 74458
rect 103428 74394 103480 74400
rect 103440 73914 103468 74394
rect 103532 74322 103560 75414
rect 103796 74928 103848 74934
rect 103796 74870 103848 74876
rect 103704 74724 103756 74730
rect 103704 74666 103756 74672
rect 103612 74656 103664 74662
rect 103612 74598 103664 74604
rect 103520 74316 103572 74322
rect 103520 74258 103572 74264
rect 103428 73908 103480 73914
rect 103428 73850 103480 73856
rect 103440 73778 103468 73850
rect 103532 73846 103560 74258
rect 103520 73840 103572 73846
rect 103520 73782 103572 73788
rect 103428 73772 103480 73778
rect 103428 73714 103480 73720
rect 103624 73710 103652 74598
rect 103612 73704 103664 73710
rect 103612 73646 103664 73652
rect 103520 73568 103572 73574
rect 103520 73510 103572 73516
rect 103336 73364 103388 73370
rect 103336 73306 103388 73312
rect 103244 73160 103296 73166
rect 103244 73102 103296 73108
rect 102784 72752 102836 72758
rect 102784 72694 102836 72700
rect 103060 72480 103112 72486
rect 103060 72422 103112 72428
rect 103152 72480 103204 72486
rect 103152 72422 103204 72428
rect 103072 72078 103100 72422
rect 103164 72078 103192 72422
rect 103256 72282 103284 73102
rect 103336 72616 103388 72622
rect 103336 72558 103388 72564
rect 103428 72616 103480 72622
rect 103428 72558 103480 72564
rect 103244 72276 103296 72282
rect 103244 72218 103296 72224
rect 102508 72072 102560 72078
rect 102508 72014 102560 72020
rect 103060 72072 103112 72078
rect 103060 72014 103112 72020
rect 103152 72072 103204 72078
rect 103152 72014 103204 72020
rect 102324 71936 102376 71942
rect 102324 71878 102376 71884
rect 102784 71936 102836 71942
rect 102784 71878 102836 71884
rect 102796 71602 102824 71878
rect 103256 71602 103284 72218
rect 103348 72010 103376 72558
rect 103440 72078 103468 72558
rect 103532 72554 103560 73510
rect 103612 72684 103664 72690
rect 103716 72672 103744 74666
rect 103808 73642 103836 74870
rect 103992 74866 104020 75414
rect 104176 75342 104204 75482
rect 104164 75336 104216 75342
rect 104164 75278 104216 75284
rect 104072 75268 104124 75274
rect 104072 75210 104124 75216
rect 104084 75002 104112 75210
rect 104072 74996 104124 75002
rect 104072 74938 104124 74944
rect 103980 74860 104032 74866
rect 103980 74802 104032 74808
rect 104072 74860 104124 74866
rect 104072 74802 104124 74808
rect 103980 74656 104032 74662
rect 103980 74598 104032 74604
rect 103796 73636 103848 73642
rect 103796 73578 103848 73584
rect 103808 73234 103836 73578
rect 103992 73302 104020 74598
rect 103980 73296 104032 73302
rect 103980 73238 104032 73244
rect 103796 73228 103848 73234
rect 103796 73170 103848 73176
rect 103808 72826 103836 73170
rect 103796 72820 103848 72826
rect 103796 72762 103848 72768
rect 103796 72684 103848 72690
rect 103716 72644 103796 72672
rect 103612 72626 103664 72632
rect 103796 72626 103848 72632
rect 103624 72570 103652 72626
rect 103520 72548 103572 72554
rect 103624 72542 103744 72570
rect 103520 72490 103572 72496
rect 103532 72078 103560 72490
rect 103716 72486 103744 72542
rect 103704 72480 103756 72486
rect 103704 72422 103756 72428
rect 103428 72072 103480 72078
rect 103428 72014 103480 72020
rect 103520 72072 103572 72078
rect 103520 72014 103572 72020
rect 103336 72004 103388 72010
rect 103336 71946 103388 71952
rect 103808 71942 103836 72626
rect 103992 72146 104020 73238
rect 104084 72214 104112 74802
rect 104176 74390 104204 75278
rect 104348 75200 104400 75206
rect 104348 75142 104400 75148
rect 104440 75200 104492 75206
rect 104440 75142 104492 75148
rect 104360 74730 104388 75142
rect 104452 74934 104480 75142
rect 104440 74928 104492 74934
rect 104440 74870 104492 74876
rect 104348 74724 104400 74730
rect 104348 74666 104400 74672
rect 104164 74384 104216 74390
rect 104164 74326 104216 74332
rect 104360 74186 104388 74666
rect 104452 74254 104480 74870
rect 104820 74866 104848 75482
rect 107764 75342 107792 80718
rect 108500 80374 108528 80718
rect 108488 80368 108540 80374
rect 108486 80336 108488 80345
rect 108540 80336 108542 80345
rect 108486 80271 108542 80280
rect 108394 79656 108450 79665
rect 108394 79591 108450 79600
rect 108408 79558 108436 79591
rect 108396 79552 108448 79558
rect 108396 79494 108448 79500
rect 108396 79008 108448 79014
rect 108394 78976 108396 78985
rect 108448 78976 108450 78985
rect 108394 78911 108450 78920
rect 108396 78464 108448 78470
rect 108396 78406 108448 78412
rect 108408 78305 108436 78406
rect 108394 78296 108450 78305
rect 108394 78231 108450 78240
rect 108212 78124 108264 78130
rect 108212 78066 108264 78072
rect 108224 77654 108252 78066
rect 108396 77920 108448 77926
rect 108396 77862 108448 77868
rect 108212 77648 108264 77654
rect 108408 77625 108436 77862
rect 108212 77590 108264 77596
rect 108394 77616 108450 77625
rect 108394 77551 108450 77560
rect 108394 76936 108450 76945
rect 108394 76871 108396 76880
rect 108448 76871 108450 76880
rect 108396 76842 108448 76848
rect 107936 76288 107988 76294
rect 108396 76288 108448 76294
rect 107936 76230 107988 76236
rect 108394 76256 108396 76265
rect 108448 76256 108450 76265
rect 107948 75750 107976 76230
rect 108394 76191 108450 76200
rect 108396 76084 108448 76090
rect 108396 76026 108448 76032
rect 107936 75744 107988 75750
rect 107936 75686 107988 75692
rect 108408 75585 108436 76026
rect 108394 75576 108450 75585
rect 108394 75511 108450 75520
rect 107752 75336 107804 75342
rect 107752 75278 107804 75284
rect 105268 75200 105320 75206
rect 105268 75142 105320 75148
rect 108396 75200 108448 75206
rect 108396 75142 108448 75148
rect 104808 74860 104860 74866
rect 104808 74802 104860 74808
rect 104624 74792 104676 74798
rect 104992 74792 105044 74798
rect 104624 74734 104676 74740
rect 104912 74752 104992 74780
rect 104532 74384 104584 74390
rect 104532 74326 104584 74332
rect 104440 74248 104492 74254
rect 104440 74190 104492 74196
rect 104348 74180 104400 74186
rect 104348 74122 104400 74128
rect 104440 73908 104492 73914
rect 104440 73850 104492 73856
rect 104452 73234 104480 73850
rect 104440 73228 104492 73234
rect 104440 73170 104492 73176
rect 104256 73024 104308 73030
rect 104256 72966 104308 72972
rect 104268 72622 104296 72966
rect 104544 72758 104572 74326
rect 104636 73846 104664 74734
rect 104912 74254 104940 74752
rect 104992 74734 105044 74740
rect 105280 74254 105308 75142
rect 108408 74905 108436 75142
rect 108394 74896 108450 74905
rect 108394 74831 108450 74840
rect 105360 74656 105412 74662
rect 105360 74598 105412 74604
rect 105372 74322 105400 74598
rect 105360 74316 105412 74322
rect 105360 74258 105412 74264
rect 105452 74316 105504 74322
rect 105452 74258 105504 74264
rect 104900 74248 104952 74254
rect 104900 74190 104952 74196
rect 105268 74248 105320 74254
rect 105268 74190 105320 74196
rect 104624 73840 104676 73846
rect 104624 73782 104676 73788
rect 104714 73808 104770 73817
rect 104714 73743 104716 73752
rect 104768 73743 104770 73752
rect 104716 73714 104768 73720
rect 104912 73710 104940 74190
rect 104992 74112 105044 74118
rect 104992 74054 105044 74060
rect 104900 73704 104952 73710
rect 104900 73646 104952 73652
rect 104624 73636 104676 73642
rect 104624 73578 104676 73584
rect 104636 73370 104664 73578
rect 104624 73364 104676 73370
rect 104624 73306 104676 73312
rect 104624 73160 104676 73166
rect 104624 73102 104676 73108
rect 104636 72826 104664 73102
rect 104624 72820 104676 72826
rect 104624 72762 104676 72768
rect 104532 72752 104584 72758
rect 104532 72694 104584 72700
rect 104256 72616 104308 72622
rect 104256 72558 104308 72564
rect 104072 72208 104124 72214
rect 104072 72150 104124 72156
rect 103980 72140 104032 72146
rect 103980 72082 104032 72088
rect 104532 72072 104584 72078
rect 104532 72014 104584 72020
rect 103520 71936 103572 71942
rect 103520 71878 103572 71884
rect 103796 71936 103848 71942
rect 103796 71878 103848 71884
rect 104440 71936 104492 71942
rect 104440 71878 104492 71884
rect 102140 71596 102192 71602
rect 102140 71538 102192 71544
rect 102784 71596 102836 71602
rect 102784 71538 102836 71544
rect 103244 71596 103296 71602
rect 103244 71538 103296 71544
rect 102152 70990 102180 71538
rect 102796 70990 102824 71538
rect 103428 71460 103480 71466
rect 103428 71402 103480 71408
rect 103440 70990 103468 71402
rect 101956 70984 102008 70990
rect 101956 70926 102008 70932
rect 102140 70984 102192 70990
rect 102140 70926 102192 70932
rect 102784 70984 102836 70990
rect 102784 70926 102836 70932
rect 103428 70984 103480 70990
rect 103532 70961 103560 71878
rect 104452 71602 104480 71878
rect 104544 71738 104572 72014
rect 104532 71732 104584 71738
rect 104532 71674 104584 71680
rect 104636 71602 104664 72762
rect 104808 72684 104860 72690
rect 104808 72626 104860 72632
rect 104716 72616 104768 72622
rect 104716 72558 104768 72564
rect 104728 72282 104756 72558
rect 104716 72276 104768 72282
rect 104716 72218 104768 72224
rect 104728 71602 104756 72218
rect 104820 71942 104848 72626
rect 104900 72004 104952 72010
rect 104900 71946 104952 71952
rect 104808 71936 104860 71942
rect 104808 71878 104860 71884
rect 104912 71670 104940 71946
rect 104900 71664 104952 71670
rect 104900 71606 104952 71612
rect 105004 71618 105032 74054
rect 105464 73914 105492 74258
rect 108394 74216 108450 74225
rect 108394 74151 108450 74160
rect 108408 74118 108436 74151
rect 108396 74112 108448 74118
rect 108396 74054 108448 74060
rect 105452 73908 105504 73914
rect 105452 73850 105504 73856
rect 105912 73908 105964 73914
rect 105912 73850 105964 73856
rect 105176 73772 105228 73778
rect 105176 73714 105228 73720
rect 105360 73772 105412 73778
rect 105544 73772 105596 73778
rect 105360 73714 105412 73720
rect 105464 73732 105544 73760
rect 105188 72826 105216 73714
rect 105268 73636 105320 73642
rect 105268 73578 105320 73584
rect 105280 73030 105308 73578
rect 105268 73024 105320 73030
rect 105268 72966 105320 72972
rect 105176 72820 105228 72826
rect 105176 72762 105228 72768
rect 105188 72554 105216 72762
rect 105176 72548 105228 72554
rect 105176 72490 105228 72496
rect 105280 72078 105308 72966
rect 105372 72826 105400 73714
rect 105464 73302 105492 73732
rect 105544 73714 105596 73720
rect 105452 73296 105504 73302
rect 105452 73238 105504 73244
rect 105464 72826 105492 73238
rect 105636 73160 105688 73166
rect 105636 73102 105688 73108
rect 105648 73030 105676 73102
rect 105636 73024 105688 73030
rect 105636 72966 105688 72972
rect 105360 72820 105412 72826
rect 105360 72762 105412 72768
rect 105452 72820 105504 72826
rect 105452 72762 105504 72768
rect 105464 72690 105492 72762
rect 105452 72684 105504 72690
rect 105452 72626 105504 72632
rect 105648 72078 105676 72966
rect 105924 72690 105952 73850
rect 108488 73772 108540 73778
rect 108488 73714 108540 73720
rect 108500 73545 108528 73714
rect 108486 73536 108542 73545
rect 108486 73471 108542 73480
rect 108120 73160 108172 73166
rect 108120 73102 108172 73108
rect 108488 73160 108540 73166
rect 108488 73102 108540 73108
rect 106004 72820 106056 72826
rect 106004 72762 106056 72768
rect 105912 72684 105964 72690
rect 105912 72626 105964 72632
rect 106016 72486 106044 72762
rect 105820 72480 105872 72486
rect 105820 72422 105872 72428
rect 106004 72480 106056 72486
rect 106004 72422 106056 72428
rect 106096 72480 106148 72486
rect 106096 72422 106148 72428
rect 105832 72078 105860 72422
rect 106004 72140 106056 72146
rect 106004 72082 106056 72088
rect 105268 72072 105320 72078
rect 105268 72014 105320 72020
rect 105360 72072 105412 72078
rect 105636 72072 105688 72078
rect 105360 72014 105412 72020
rect 105464 72032 105636 72060
rect 105004 71602 105124 71618
rect 105372 71602 105400 72014
rect 103796 71596 103848 71602
rect 103796 71538 103848 71544
rect 104440 71596 104492 71602
rect 104440 71538 104492 71544
rect 104624 71596 104676 71602
rect 104624 71538 104676 71544
rect 104716 71596 104768 71602
rect 104716 71538 104768 71544
rect 104992 71596 105124 71602
rect 105044 71590 105124 71596
rect 104992 71538 105044 71544
rect 103808 71058 103836 71538
rect 104992 71460 105044 71466
rect 104992 71402 105044 71408
rect 103888 71392 103940 71398
rect 103888 71334 103940 71340
rect 104900 71392 104952 71398
rect 104900 71334 104952 71340
rect 103612 71052 103664 71058
rect 103612 70994 103664 71000
rect 103796 71052 103848 71058
rect 103796 70994 103848 71000
rect 103428 70926 103480 70932
rect 103518 70952 103574 70961
rect 101864 70440 101916 70446
rect 101864 70382 101916 70388
rect 101968 70106 101996 70926
rect 102152 70514 102180 70926
rect 103060 70916 103112 70922
rect 103518 70887 103574 70896
rect 103060 70858 103112 70864
rect 102140 70508 102192 70514
rect 102140 70450 102192 70456
rect 102324 70372 102376 70378
rect 102324 70314 102376 70320
rect 101956 70100 102008 70106
rect 101956 70042 102008 70048
rect 101404 69964 101456 69970
rect 101404 69906 101456 69912
rect 101956 69964 102008 69970
rect 101956 69906 102008 69912
rect 101312 69896 101364 69902
rect 101312 69838 101364 69844
rect 101496 69896 101548 69902
rect 101496 69838 101548 69844
rect 101128 68808 101180 68814
rect 101128 68750 101180 68756
rect 101220 68808 101272 68814
rect 101220 68750 101272 68756
rect 100944 68740 100996 68746
rect 100996 68700 101076 68728
rect 100944 68682 100996 68688
rect 100850 68368 100906 68377
rect 100668 68332 100720 68338
rect 100850 68303 100852 68312
rect 100668 68274 100720 68280
rect 100904 68303 100906 68312
rect 100852 68274 100904 68280
rect 100576 68128 100628 68134
rect 100576 68070 100628 68076
rect 100576 67108 100628 67114
rect 100576 67050 100628 67056
rect 100588 66842 100616 67050
rect 100680 67046 100708 68274
rect 101048 68270 101076 68700
rect 101128 68672 101180 68678
rect 101128 68614 101180 68620
rect 101220 68672 101272 68678
rect 101220 68614 101272 68620
rect 101140 68338 101168 68614
rect 101232 68406 101260 68614
rect 101220 68400 101272 68406
rect 101220 68342 101272 68348
rect 101128 68332 101180 68338
rect 101128 68274 101180 68280
rect 101036 68264 101088 68270
rect 101036 68206 101088 68212
rect 100760 67856 100812 67862
rect 100760 67798 100812 67804
rect 100772 67130 100800 67798
rect 101048 67726 101076 68206
rect 101036 67720 101088 67726
rect 100850 67688 100906 67697
rect 101036 67662 101088 67668
rect 100850 67623 100906 67632
rect 100864 67590 100892 67623
rect 100852 67584 100904 67590
rect 100852 67526 100904 67532
rect 100864 67250 100892 67526
rect 101324 67318 101352 69838
rect 101508 69426 101536 69838
rect 101680 69828 101732 69834
rect 101680 69770 101732 69776
rect 101496 69420 101548 69426
rect 101496 69362 101548 69368
rect 101404 68876 101456 68882
rect 101404 68818 101456 68824
rect 101416 68406 101444 68818
rect 101404 68400 101456 68406
rect 101404 68342 101456 68348
rect 101692 67930 101720 69770
rect 101772 69216 101824 69222
rect 101772 69158 101824 69164
rect 101784 68882 101812 69158
rect 101772 68876 101824 68882
rect 101772 68818 101824 68824
rect 101864 68468 101916 68474
rect 101864 68410 101916 68416
rect 101680 67924 101732 67930
rect 101680 67866 101732 67872
rect 101772 67924 101824 67930
rect 101772 67866 101824 67872
rect 101680 67720 101732 67726
rect 101680 67662 101732 67668
rect 101312 67312 101364 67318
rect 101312 67254 101364 67260
rect 100852 67244 100904 67250
rect 100852 67186 100904 67192
rect 100944 67176 100996 67182
rect 100772 67124 100944 67130
rect 100772 67118 100996 67124
rect 100772 67102 100984 67118
rect 100668 67040 100720 67046
rect 100668 66982 100720 66988
rect 100576 66836 100628 66842
rect 100576 66778 100628 66784
rect 100484 66700 100536 66706
rect 100484 66642 100536 66648
rect 100680 66638 100708 66982
rect 100668 66632 100720 66638
rect 100668 66574 100720 66580
rect 100576 66496 100628 66502
rect 100576 66438 100628 66444
rect 99932 66088 99984 66094
rect 99932 66030 99984 66036
rect 100300 66088 100352 66094
rect 100300 66030 100352 66036
rect 96896 66020 96948 66026
rect 96896 65962 96948 65968
rect 99380 66020 99432 66026
rect 99380 65962 99432 65968
rect 99748 66020 99800 66026
rect 99748 65962 99800 65968
rect 100588 65958 100616 66438
rect 100772 66230 100800 67102
rect 100852 66700 100904 66706
rect 100852 66642 100904 66648
rect 100760 66224 100812 66230
rect 100760 66166 100812 66172
rect 100864 66162 100892 66642
rect 101692 66570 101720 67662
rect 101784 67250 101812 67866
rect 101876 67708 101904 68410
rect 101968 68202 101996 69906
rect 102232 69760 102284 69766
rect 102232 69702 102284 69708
rect 102048 69352 102100 69358
rect 102048 69294 102100 69300
rect 102060 68678 102088 69294
rect 102244 68882 102272 69702
rect 102336 69426 102364 70314
rect 102324 69420 102376 69426
rect 102324 69362 102376 69368
rect 102416 69352 102468 69358
rect 102416 69294 102468 69300
rect 102968 69352 103020 69358
rect 102968 69294 103020 69300
rect 102232 68876 102284 68882
rect 102232 68818 102284 68824
rect 102048 68672 102100 68678
rect 102048 68614 102100 68620
rect 101956 68196 102008 68202
rect 101956 68138 102008 68144
rect 101956 67720 102008 67726
rect 101876 67680 101956 67708
rect 101772 67244 101824 67250
rect 101772 67186 101824 67192
rect 101876 66774 101904 67680
rect 101956 67662 102008 67668
rect 101956 67312 102008 67318
rect 101956 67254 102008 67260
rect 101864 66768 101916 66774
rect 101864 66710 101916 66716
rect 101680 66564 101732 66570
rect 101680 66506 101732 66512
rect 101312 66496 101364 66502
rect 101312 66438 101364 66444
rect 101324 66230 101352 66438
rect 101312 66224 101364 66230
rect 101312 66166 101364 66172
rect 101968 66162 101996 67254
rect 102060 67046 102088 68614
rect 102428 68474 102456 69294
rect 102980 69018 103008 69294
rect 102968 69012 103020 69018
rect 102968 68954 103020 68960
rect 103072 68814 103100 70858
rect 103152 70848 103204 70854
rect 103152 70790 103204 70796
rect 103164 70446 103192 70790
rect 103152 70440 103204 70446
rect 103152 70382 103204 70388
rect 103164 68882 103192 70382
rect 103336 69760 103388 69766
rect 103336 69702 103388 69708
rect 103348 69426 103376 69702
rect 103532 69426 103560 70887
rect 103624 70650 103652 70994
rect 103612 70644 103664 70650
rect 103612 70586 103664 70592
rect 103624 69970 103652 70586
rect 103900 70514 103928 71334
rect 103888 70508 103940 70514
rect 103888 70450 103940 70456
rect 103612 69964 103664 69970
rect 103612 69906 103664 69912
rect 104912 69902 104940 71334
rect 105004 70446 105032 71402
rect 105096 70922 105124 71590
rect 105360 71596 105412 71602
rect 105360 71538 105412 71544
rect 105360 71392 105412 71398
rect 105360 71334 105412 71340
rect 105268 71052 105320 71058
rect 105268 70994 105320 71000
rect 105084 70916 105136 70922
rect 105084 70858 105136 70864
rect 105280 70650 105308 70994
rect 105268 70644 105320 70650
rect 105268 70586 105320 70592
rect 105084 70508 105136 70514
rect 105084 70450 105136 70456
rect 104992 70440 105044 70446
rect 104992 70382 105044 70388
rect 105004 69970 105032 70382
rect 104992 69964 105044 69970
rect 104992 69906 105044 69912
rect 105096 69902 105124 70450
rect 105176 70304 105228 70310
rect 105176 70246 105228 70252
rect 104900 69896 104952 69902
rect 104900 69838 104952 69844
rect 105084 69896 105136 69902
rect 105084 69838 105136 69844
rect 104900 69760 104952 69766
rect 104900 69702 104952 69708
rect 105188 69714 105216 70246
rect 105280 69902 105308 70586
rect 105372 70446 105400 71334
rect 105360 70440 105412 70446
rect 105360 70382 105412 70388
rect 105268 69896 105320 69902
rect 105268 69838 105320 69844
rect 103244 69420 103296 69426
rect 103244 69362 103296 69368
rect 103336 69420 103388 69426
rect 103336 69362 103388 69368
rect 103520 69420 103572 69426
rect 103520 69362 103572 69368
rect 104624 69420 104676 69426
rect 104624 69362 104676 69368
rect 103152 68876 103204 68882
rect 103152 68818 103204 68824
rect 103256 68814 103284 69362
rect 103060 68808 103112 68814
rect 103060 68750 103112 68756
rect 103244 68808 103296 68814
rect 103244 68750 103296 68756
rect 102876 68672 102928 68678
rect 102876 68614 102928 68620
rect 102324 68468 102376 68474
rect 102324 68410 102376 68416
rect 102416 68468 102468 68474
rect 102416 68410 102468 68416
rect 102232 68332 102284 68338
rect 102232 68274 102284 68280
rect 102138 67824 102194 67833
rect 102138 67759 102194 67768
rect 102152 67726 102180 67759
rect 102244 67726 102272 68274
rect 102336 67794 102364 68410
rect 102508 68196 102560 68202
rect 102508 68138 102560 68144
rect 102324 67788 102376 67794
rect 102324 67730 102376 67736
rect 102520 67726 102548 68138
rect 102692 67924 102744 67930
rect 102692 67866 102744 67872
rect 102704 67726 102732 67866
rect 102888 67862 102916 68614
rect 102876 67856 102928 67862
rect 102968 67856 103020 67862
rect 102876 67798 102928 67804
rect 102966 67824 102968 67833
rect 103020 67824 103022 67833
rect 102140 67720 102192 67726
rect 102140 67662 102192 67668
rect 102232 67720 102284 67726
rect 102232 67662 102284 67668
rect 102508 67720 102560 67726
rect 102692 67720 102744 67726
rect 102560 67680 102640 67708
rect 102508 67662 102560 67668
rect 102244 67250 102272 67662
rect 102416 67652 102468 67658
rect 102416 67594 102468 67600
rect 102428 67386 102456 67594
rect 102416 67380 102468 67386
rect 102416 67322 102468 67328
rect 102612 67250 102640 67680
rect 102692 67662 102744 67668
rect 102784 67720 102836 67726
rect 102784 67662 102836 67668
rect 102796 67386 102824 67662
rect 102784 67380 102836 67386
rect 102784 67322 102836 67328
rect 102888 67318 102916 67798
rect 102966 67759 103022 67768
rect 102876 67312 102928 67318
rect 103072 67266 103100 68750
rect 103348 68490 103376 69362
rect 103428 69216 103480 69222
rect 103428 69158 103480 69164
rect 103612 69216 103664 69222
rect 103612 69158 103664 69164
rect 104532 69216 104584 69222
rect 104532 69158 104584 69164
rect 103440 68814 103468 69158
rect 103624 68814 103652 69158
rect 103428 68808 103480 68814
rect 103428 68750 103480 68756
rect 103612 68808 103664 68814
rect 103612 68750 103664 68756
rect 103704 68808 103756 68814
rect 103704 68750 103756 68756
rect 103256 68462 103376 68490
rect 103152 67584 103204 67590
rect 103152 67526 103204 67532
rect 102876 67254 102928 67260
rect 102232 67244 102284 67250
rect 102232 67186 102284 67192
rect 102600 67244 102652 67250
rect 102600 67186 102652 67192
rect 102048 67040 102100 67046
rect 102048 66982 102100 66988
rect 102140 66836 102192 66842
rect 102140 66778 102192 66784
rect 100852 66156 100904 66162
rect 100852 66098 100904 66104
rect 101956 66156 102008 66162
rect 101956 66098 102008 66104
rect 95976 65952 96028 65958
rect 95976 65894 96028 65900
rect 100576 65952 100628 65958
rect 100576 65894 100628 65900
rect 96374 65852 96682 65861
rect 96374 65850 96380 65852
rect 96436 65850 96460 65852
rect 96516 65850 96540 65852
rect 96596 65850 96620 65852
rect 96676 65850 96682 65852
rect 96436 65798 96438 65850
rect 96618 65798 96620 65850
rect 96374 65796 96380 65798
rect 96436 65796 96460 65798
rect 96516 65796 96540 65798
rect 96596 65796 96620 65798
rect 96676 65796 96682 65798
rect 96374 65787 96682 65796
rect 95882 64152 95938 64161
rect 95882 64087 95938 64096
rect 77850 63880 77906 63889
rect 77850 63815 77906 63824
rect 102152 22778 102180 66778
rect 102244 66706 102272 67186
rect 102888 67046 102916 67254
rect 102980 67250 103100 67266
rect 102968 67244 103100 67250
rect 103020 67238 103100 67244
rect 102968 67186 103020 67192
rect 102876 67040 102928 67046
rect 102796 66988 102876 66994
rect 102796 66982 102928 66988
rect 102796 66966 102916 66982
rect 102796 66774 102824 66966
rect 102980 66858 103008 67186
rect 103164 67182 103192 67526
rect 103152 67176 103204 67182
rect 103152 67118 103204 67124
rect 102888 66830 103008 66858
rect 103164 66842 103192 67118
rect 103152 66836 103204 66842
rect 102784 66768 102836 66774
rect 102784 66710 102836 66716
rect 102232 66700 102284 66706
rect 102232 66642 102284 66648
rect 102796 66638 102824 66710
rect 102888 66638 102916 66830
rect 103152 66778 103204 66784
rect 103256 66706 103284 68462
rect 103336 68332 103388 68338
rect 103440 68320 103468 68750
rect 103624 68474 103652 68750
rect 103612 68468 103664 68474
rect 103612 68410 103664 68416
rect 103716 68338 103744 68750
rect 104440 68672 104492 68678
rect 104440 68614 104492 68620
rect 103388 68292 103468 68320
rect 103704 68332 103756 68338
rect 103336 68274 103388 68280
rect 103704 68274 103756 68280
rect 103980 68128 104032 68134
rect 103980 68070 104032 68076
rect 103704 67720 103756 67726
rect 103704 67662 103756 67668
rect 103336 67652 103388 67658
rect 103336 67594 103388 67600
rect 103244 66700 103296 66706
rect 103244 66642 103296 66648
rect 103348 66638 103376 67594
rect 103520 67312 103572 67318
rect 103520 67254 103572 67260
rect 102784 66632 102836 66638
rect 102784 66574 102836 66580
rect 102876 66632 102928 66638
rect 102876 66574 102928 66580
rect 103336 66632 103388 66638
rect 103336 66574 103388 66580
rect 102796 66230 102824 66574
rect 102784 66224 102836 66230
rect 102784 66166 102836 66172
rect 102888 66162 102916 66574
rect 102876 66156 102928 66162
rect 102876 66098 102928 66104
rect 103532 66094 103560 67254
rect 103716 67250 103744 67662
rect 103992 67318 104020 68070
rect 104452 67946 104480 68614
rect 104544 68270 104572 69158
rect 104636 68814 104664 69362
rect 104808 69012 104860 69018
rect 104808 68954 104860 68960
rect 104820 68814 104848 68954
rect 104624 68808 104676 68814
rect 104624 68750 104676 68756
rect 104808 68808 104860 68814
rect 104808 68750 104860 68756
rect 104532 68264 104584 68270
rect 104532 68206 104584 68212
rect 104636 68202 104664 68750
rect 104912 68746 104940 69702
rect 105188 69686 105308 69714
rect 104992 69420 105044 69426
rect 104992 69362 105044 69368
rect 105004 69018 105032 69362
rect 105280 69018 105308 69686
rect 104992 69012 105044 69018
rect 104992 68954 105044 68960
rect 105268 69012 105320 69018
rect 105268 68954 105320 68960
rect 104900 68740 104952 68746
rect 104900 68682 104952 68688
rect 105176 68740 105228 68746
rect 105176 68682 105228 68688
rect 104898 68368 104954 68377
rect 105188 68338 105216 68682
rect 105280 68474 105308 68954
rect 105372 68882 105400 70382
rect 105360 68876 105412 68882
rect 105360 68818 105412 68824
rect 105464 68746 105492 72032
rect 105636 72014 105688 72020
rect 105820 72072 105872 72078
rect 105820 72014 105872 72020
rect 106016 71942 106044 72082
rect 106108 72010 106136 72422
rect 107292 72208 107344 72214
rect 107292 72150 107344 72156
rect 106096 72004 106148 72010
rect 106096 71946 106148 71952
rect 105544 71936 105596 71942
rect 105544 71878 105596 71884
rect 105820 71936 105872 71942
rect 105820 71878 105872 71884
rect 106004 71936 106056 71942
rect 106004 71878 106056 71884
rect 105556 71058 105584 71878
rect 105728 71596 105780 71602
rect 105728 71538 105780 71544
rect 105544 71052 105596 71058
rect 105544 70994 105596 71000
rect 105556 70922 105584 70994
rect 105544 70916 105596 70922
rect 105544 70858 105596 70864
rect 105636 70848 105688 70854
rect 105636 70790 105688 70796
rect 105648 70582 105676 70790
rect 105544 70576 105596 70582
rect 105544 70518 105596 70524
rect 105636 70576 105688 70582
rect 105636 70518 105688 70524
rect 105556 70378 105584 70518
rect 105544 70372 105596 70378
rect 105544 70314 105596 70320
rect 105636 70304 105688 70310
rect 105636 70246 105688 70252
rect 105648 69834 105676 70246
rect 105740 70106 105768 71538
rect 105832 71194 105860 71878
rect 106016 71534 106044 71878
rect 106004 71528 106056 71534
rect 106004 71470 106056 71476
rect 106280 71392 106332 71398
rect 106280 71334 106332 71340
rect 105820 71188 105872 71194
rect 105820 71130 105872 71136
rect 105832 70990 105860 71130
rect 106004 71120 106056 71126
rect 106004 71062 106056 71068
rect 105820 70984 105872 70990
rect 105820 70926 105872 70932
rect 106016 70582 106044 71062
rect 106188 71052 106240 71058
rect 106188 70994 106240 71000
rect 106200 70650 106228 70994
rect 106188 70644 106240 70650
rect 106188 70586 106240 70592
rect 106004 70576 106056 70582
rect 106004 70518 106056 70524
rect 106292 70514 106320 71334
rect 107304 71194 107332 72150
rect 107292 71188 107344 71194
rect 107292 71130 107344 71136
rect 108132 70650 108160 73102
rect 108500 72865 108528 73102
rect 108486 72856 108542 72865
rect 108486 72791 108542 72800
rect 108488 72684 108540 72690
rect 108488 72626 108540 72632
rect 108304 72480 108356 72486
rect 108304 72422 108356 72428
rect 108316 71602 108344 72422
rect 108500 72185 108528 72626
rect 108486 72176 108542 72185
rect 108486 72111 108542 72120
rect 108304 71596 108356 71602
rect 108304 71538 108356 71544
rect 108488 71596 108540 71602
rect 108488 71538 108540 71544
rect 108500 71505 108528 71538
rect 108486 71496 108542 71505
rect 108486 71431 108542 71440
rect 108488 70984 108540 70990
rect 108488 70926 108540 70932
rect 108500 70825 108528 70926
rect 108486 70816 108542 70825
rect 108486 70751 108542 70760
rect 108120 70644 108172 70650
rect 108120 70586 108172 70592
rect 106280 70508 106332 70514
rect 106280 70450 106332 70456
rect 108488 70508 108540 70514
rect 108488 70450 108540 70456
rect 107936 70440 107988 70446
rect 107936 70382 107988 70388
rect 105728 70100 105780 70106
rect 105728 70042 105780 70048
rect 105636 69828 105688 69834
rect 105636 69770 105688 69776
rect 105452 68740 105504 68746
rect 105452 68682 105504 68688
rect 105268 68468 105320 68474
rect 105268 68410 105320 68416
rect 104898 68303 104900 68312
rect 104952 68303 104954 68312
rect 105176 68332 105228 68338
rect 104900 68274 104952 68280
rect 105176 68274 105228 68280
rect 105464 68270 105492 68682
rect 105452 68264 105504 68270
rect 105452 68206 105504 68212
rect 104624 68196 104676 68202
rect 104624 68138 104676 68144
rect 104452 67918 104664 67946
rect 107948 67930 107976 70382
rect 108500 70145 108528 70450
rect 108486 70136 108542 70145
rect 108486 70071 108542 70080
rect 108488 69896 108540 69902
rect 108488 69838 108540 69844
rect 108500 69465 108528 69838
rect 108486 69456 108542 69465
rect 108486 69391 108542 69400
rect 103980 67312 104032 67318
rect 103980 67254 104032 67260
rect 103704 67244 103756 67250
rect 103704 67186 103756 67192
rect 103716 66842 103744 67186
rect 103704 66836 103756 66842
rect 103704 66778 103756 66784
rect 104636 66570 104664 67918
rect 107936 67924 107988 67930
rect 107936 67866 107988 67872
rect 108488 67720 108540 67726
rect 108488 67662 108540 67668
rect 108500 67425 108528 67662
rect 108486 67416 108542 67425
rect 108486 67351 108542 67360
rect 104164 66564 104216 66570
rect 104164 66506 104216 66512
rect 104624 66564 104676 66570
rect 104624 66506 104676 66512
rect 103704 66496 103756 66502
rect 103704 66438 103756 66444
rect 103716 66162 103744 66438
rect 104176 66298 104204 66506
rect 103980 66292 104032 66298
rect 103980 66234 104032 66240
rect 104164 66292 104216 66298
rect 104164 66234 104216 66240
rect 103704 66156 103756 66162
rect 103704 66098 103756 66104
rect 103520 66088 103572 66094
rect 103520 66030 103572 66036
rect 103704 66020 103756 66026
rect 103704 65962 103756 65968
rect 103612 65748 103664 65754
rect 103612 65690 103664 65696
rect 102232 65680 102284 65686
rect 102232 65622 102284 65628
rect 102244 25097 102272 65622
rect 102600 25152 102652 25158
rect 102598 25120 102600 25129
rect 102652 25120 102654 25129
rect 102230 25088 102286 25097
rect 102598 25055 102654 25064
rect 102230 25023 102286 25032
rect 102784 23520 102836 23526
rect 102782 23488 102784 23497
rect 102836 23488 102838 23497
rect 102782 23423 102838 23432
rect 102140 22772 102192 22778
rect 102140 22714 102192 22720
rect 102152 22269 102180 22714
rect 102138 22260 102194 22269
rect 102138 22195 102194 22204
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29564 9761 29592 9862
rect 23478 9752 23534 9761
rect 23478 9687 23534 9696
rect 25778 9752 25834 9761
rect 25778 9687 25834 9696
rect 28170 9752 28226 9761
rect 28170 9687 28226 9696
rect 29550 9752 29606 9761
rect 29550 9687 29606 9696
rect 30470 9752 30526 9761
rect 30470 9687 30526 9696
rect 16028 9648 16080 9654
rect 16026 9616 16028 9625
rect 16080 9616 16082 9625
rect 9588 9580 9640 9586
rect 16026 9551 16082 9560
rect 16120 9580 16172 9586
rect 9588 9522 9640 9528
rect 16040 7546 16068 9551
rect 16120 9522 16172 9528
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1320 4865 1348 5170
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 1306 4856 1362 4865
rect 4214 4859 4522 4868
rect 1306 4791 1362 4800
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 16132 800 16160 9522
rect 23492 7546 23520 9687
rect 24674 9616 24730 9625
rect 24674 9551 24730 9560
rect 24688 8362 24716 9551
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24688 7546 24716 8298
rect 25792 7546 25820 9687
rect 26698 8936 26754 8945
rect 26698 8871 26754 8880
rect 26712 8838 26740 8871
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 26712 7546 26740 8774
rect 28184 7546 28212 9687
rect 29564 7546 29592 9687
rect 30484 7750 30512 9687
rect 90638 9616 90694 9625
rect 90638 9551 90694 9560
rect 90822 9616 90878 9625
rect 90822 9551 90878 9560
rect 90652 9042 90680 9551
rect 90836 9110 90864 9551
rect 90824 9104 90876 9110
rect 90824 9046 90876 9052
rect 90640 9036 90692 9042
rect 90640 8978 90692 8984
rect 90548 8968 90600 8974
rect 90548 8910 90600 8916
rect 90560 8401 90588 8910
rect 90546 8392 90602 8401
rect 90546 8327 90602 8336
rect 31666 8256 31722 8265
rect 31666 8191 31722 8200
rect 32954 8256 33010 8265
rect 32954 8191 33010 8200
rect 34242 8256 34298 8265
rect 34242 8191 34298 8200
rect 35438 8256 35494 8265
rect 35438 8191 35494 8200
rect 36358 8256 36414 8265
rect 36358 8191 36414 8200
rect 37462 8256 37518 8265
rect 37462 8191 37518 8200
rect 38750 8256 38806 8265
rect 38750 8191 38806 8200
rect 41326 8256 41382 8265
rect 41326 8191 41382 8200
rect 42154 8256 42210 8265
rect 42154 8191 42210 8200
rect 43442 8256 43498 8265
rect 43442 8191 43498 8200
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 30484 7546 30512 7686
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 23492 5030 23520 7482
rect 25792 6914 25820 7482
rect 28184 7274 28212 7482
rect 28172 7268 28224 7274
rect 28172 7210 28224 7216
rect 25792 6886 25912 6914
rect 25884 6118 25912 6886
rect 25872 6112 25924 6118
rect 25872 6054 25924 6060
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 31680 2650 31708 8191
rect 32968 2650 32996 8191
rect 34256 2650 34284 8191
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35452 2650 35480 8191
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 36372 2650 36400 8191
rect 37476 2650 37504 8191
rect 38764 2650 38792 8191
rect 39946 4584 40002 4593
rect 39946 4519 40002 4528
rect 39960 2650 39988 4519
rect 41340 2650 41368 8191
rect 42168 2650 42196 8191
rect 43456 2650 43484 8191
rect 66314 7644 66622 7653
rect 66314 7642 66320 7644
rect 66376 7642 66400 7644
rect 66456 7642 66480 7644
rect 66536 7642 66560 7644
rect 66616 7642 66622 7644
rect 66376 7590 66378 7642
rect 66558 7590 66560 7642
rect 66314 7588 66320 7590
rect 66376 7588 66400 7590
rect 66456 7588 66480 7590
rect 66536 7588 66560 7590
rect 66616 7588 66622 7590
rect 66314 7579 66622 7588
rect 90560 7546 90588 8327
rect 90652 7546 90680 8978
rect 90836 7546 90864 9046
rect 103624 8974 103652 65690
rect 103716 9042 103744 65962
rect 103992 9110 104020 66234
rect 104636 66162 104664 66506
rect 106658 66396 106966 66405
rect 106658 66394 106664 66396
rect 106720 66394 106744 66396
rect 106800 66394 106824 66396
rect 106880 66394 106904 66396
rect 106960 66394 106966 66396
rect 106720 66342 106722 66394
rect 106902 66342 106904 66394
rect 106658 66340 106664 66342
rect 106720 66340 106744 66342
rect 106800 66340 106824 66342
rect 106880 66340 106904 66342
rect 106960 66340 106966 66342
rect 106658 66331 106966 66340
rect 104624 66156 104676 66162
rect 104624 66098 104676 66104
rect 105922 65852 106230 65861
rect 105922 65850 105928 65852
rect 105984 65850 106008 65852
rect 106064 65850 106088 65852
rect 106144 65850 106168 65852
rect 106224 65850 106230 65852
rect 105984 65798 105986 65850
rect 106166 65798 106168 65850
rect 105922 65796 105928 65798
rect 105984 65796 106008 65798
rect 106064 65796 106088 65798
rect 106144 65796 106168 65798
rect 106224 65796 106230 65798
rect 105922 65787 106230 65796
rect 106658 65308 106966 65317
rect 106658 65306 106664 65308
rect 106720 65306 106744 65308
rect 106800 65306 106824 65308
rect 106880 65306 106904 65308
rect 106960 65306 106966 65308
rect 106720 65254 106722 65306
rect 106902 65254 106904 65306
rect 106658 65252 106664 65254
rect 106720 65252 106744 65254
rect 106800 65252 106824 65254
rect 106880 65252 106904 65254
rect 106960 65252 106966 65254
rect 106658 65243 106966 65252
rect 105922 64764 106230 64773
rect 105922 64762 105928 64764
rect 105984 64762 106008 64764
rect 106064 64762 106088 64764
rect 106144 64762 106168 64764
rect 106224 64762 106230 64764
rect 105984 64710 105986 64762
rect 106166 64710 106168 64762
rect 105922 64708 105928 64710
rect 105984 64708 106008 64710
rect 106064 64708 106088 64710
rect 106144 64708 106168 64710
rect 106224 64708 106230 64710
rect 105922 64699 106230 64708
rect 106658 64220 106966 64229
rect 106658 64218 106664 64220
rect 106720 64218 106744 64220
rect 106800 64218 106824 64220
rect 106880 64218 106904 64220
rect 106960 64218 106966 64220
rect 106720 64166 106722 64218
rect 106902 64166 106904 64218
rect 106658 64164 106664 64166
rect 106720 64164 106744 64166
rect 106800 64164 106824 64166
rect 106880 64164 106904 64166
rect 106960 64164 106966 64166
rect 106658 64155 106966 64164
rect 105922 63676 106230 63685
rect 105922 63674 105928 63676
rect 105984 63674 106008 63676
rect 106064 63674 106088 63676
rect 106144 63674 106168 63676
rect 106224 63674 106230 63676
rect 105984 63622 105986 63674
rect 106166 63622 106168 63674
rect 105922 63620 105928 63622
rect 105984 63620 106008 63622
rect 106064 63620 106088 63622
rect 106144 63620 106168 63622
rect 106224 63620 106230 63622
rect 105922 63611 106230 63620
rect 106658 63132 106966 63141
rect 106658 63130 106664 63132
rect 106720 63130 106744 63132
rect 106800 63130 106824 63132
rect 106880 63130 106904 63132
rect 106960 63130 106966 63132
rect 106720 63078 106722 63130
rect 106902 63078 106904 63130
rect 106658 63076 106664 63078
rect 106720 63076 106744 63078
rect 106800 63076 106824 63078
rect 106880 63076 106904 63078
rect 106960 63076 106966 63078
rect 106658 63067 106966 63076
rect 105922 62588 106230 62597
rect 105922 62586 105928 62588
rect 105984 62586 106008 62588
rect 106064 62586 106088 62588
rect 106144 62586 106168 62588
rect 106224 62586 106230 62588
rect 105984 62534 105986 62586
rect 106166 62534 106168 62586
rect 105922 62532 105928 62534
rect 105984 62532 106008 62534
rect 106064 62532 106088 62534
rect 106144 62532 106168 62534
rect 106224 62532 106230 62534
rect 105922 62523 106230 62532
rect 106658 62044 106966 62053
rect 106658 62042 106664 62044
rect 106720 62042 106744 62044
rect 106800 62042 106824 62044
rect 106880 62042 106904 62044
rect 106960 62042 106966 62044
rect 106720 61990 106722 62042
rect 106902 61990 106904 62042
rect 106658 61988 106664 61990
rect 106720 61988 106744 61990
rect 106800 61988 106824 61990
rect 106880 61988 106904 61990
rect 106960 61988 106966 61990
rect 106658 61979 106966 61988
rect 105922 61500 106230 61509
rect 105922 61498 105928 61500
rect 105984 61498 106008 61500
rect 106064 61498 106088 61500
rect 106144 61498 106168 61500
rect 106224 61498 106230 61500
rect 105984 61446 105986 61498
rect 106166 61446 106168 61498
rect 105922 61444 105928 61446
rect 105984 61444 106008 61446
rect 106064 61444 106088 61446
rect 106144 61444 106168 61446
rect 106224 61444 106230 61446
rect 105922 61435 106230 61444
rect 106658 60956 106966 60965
rect 106658 60954 106664 60956
rect 106720 60954 106744 60956
rect 106800 60954 106824 60956
rect 106880 60954 106904 60956
rect 106960 60954 106966 60956
rect 106720 60902 106722 60954
rect 106902 60902 106904 60954
rect 106658 60900 106664 60902
rect 106720 60900 106744 60902
rect 106800 60900 106824 60902
rect 106880 60900 106904 60902
rect 106960 60900 106966 60902
rect 106658 60891 106966 60900
rect 105922 60412 106230 60421
rect 105922 60410 105928 60412
rect 105984 60410 106008 60412
rect 106064 60410 106088 60412
rect 106144 60410 106168 60412
rect 106224 60410 106230 60412
rect 105984 60358 105986 60410
rect 106166 60358 106168 60410
rect 105922 60356 105928 60358
rect 105984 60356 106008 60358
rect 106064 60356 106088 60358
rect 106144 60356 106168 60358
rect 106224 60356 106230 60358
rect 105922 60347 106230 60356
rect 104348 60104 104400 60110
rect 104348 60046 104400 60052
rect 104360 59809 104388 60046
rect 106658 59868 106966 59877
rect 106658 59866 106664 59868
rect 106720 59866 106744 59868
rect 106800 59866 106824 59868
rect 106880 59866 106904 59868
rect 106960 59866 106966 59868
rect 106720 59814 106722 59866
rect 106902 59814 106904 59866
rect 106658 59812 106664 59814
rect 106720 59812 106744 59814
rect 106800 59812 106824 59814
rect 106880 59812 106904 59814
rect 106960 59812 106966 59814
rect 104346 59800 104402 59809
rect 106658 59803 106966 59812
rect 104346 59735 104402 59744
rect 105922 59324 106230 59333
rect 105922 59322 105928 59324
rect 105984 59322 106008 59324
rect 106064 59322 106088 59324
rect 106144 59322 106168 59324
rect 106224 59322 106230 59324
rect 105984 59270 105986 59322
rect 106166 59270 106168 59322
rect 105922 59268 105928 59270
rect 105984 59268 106008 59270
rect 106064 59268 106088 59270
rect 106144 59268 106168 59270
rect 106224 59268 106230 59270
rect 105922 59259 106230 59268
rect 106658 58780 106966 58789
rect 106658 58778 106664 58780
rect 106720 58778 106744 58780
rect 106800 58778 106824 58780
rect 106880 58778 106904 58780
rect 106960 58778 106966 58780
rect 106720 58726 106722 58778
rect 106902 58726 106904 58778
rect 106658 58724 106664 58726
rect 106720 58724 106744 58726
rect 106800 58724 106824 58726
rect 106880 58724 106904 58726
rect 106960 58724 106966 58726
rect 106658 58715 106966 58724
rect 105922 58236 106230 58245
rect 105922 58234 105928 58236
rect 105984 58234 106008 58236
rect 106064 58234 106088 58236
rect 106144 58234 106168 58236
rect 106224 58234 106230 58236
rect 105984 58182 105986 58234
rect 106166 58182 106168 58234
rect 105922 58180 105928 58182
rect 105984 58180 106008 58182
rect 106064 58180 106088 58182
rect 106144 58180 106168 58182
rect 106224 58180 106230 58182
rect 105922 58171 106230 58180
rect 106658 57692 106966 57701
rect 106658 57690 106664 57692
rect 106720 57690 106744 57692
rect 106800 57690 106824 57692
rect 106880 57690 106904 57692
rect 106960 57690 106966 57692
rect 106720 57638 106722 57690
rect 106902 57638 106904 57690
rect 106658 57636 106664 57638
rect 106720 57636 106744 57638
rect 106800 57636 106824 57638
rect 106880 57636 106904 57638
rect 106960 57636 106966 57638
rect 106658 57627 106966 57636
rect 105922 57148 106230 57157
rect 105922 57146 105928 57148
rect 105984 57146 106008 57148
rect 106064 57146 106088 57148
rect 106144 57146 106168 57148
rect 106224 57146 106230 57148
rect 105984 57094 105986 57146
rect 106166 57094 106168 57146
rect 105922 57092 105928 57094
rect 105984 57092 106008 57094
rect 106064 57092 106088 57094
rect 106144 57092 106168 57094
rect 106224 57092 106230 57094
rect 105922 57083 106230 57092
rect 106658 56604 106966 56613
rect 106658 56602 106664 56604
rect 106720 56602 106744 56604
rect 106800 56602 106824 56604
rect 106880 56602 106904 56604
rect 106960 56602 106966 56604
rect 106720 56550 106722 56602
rect 106902 56550 106904 56602
rect 106658 56548 106664 56550
rect 106720 56548 106744 56550
rect 106800 56548 106824 56550
rect 106880 56548 106904 56550
rect 106960 56548 106966 56550
rect 106658 56539 106966 56548
rect 105922 56060 106230 56069
rect 105922 56058 105928 56060
rect 105984 56058 106008 56060
rect 106064 56058 106088 56060
rect 106144 56058 106168 56060
rect 106224 56058 106230 56060
rect 105984 56006 105986 56058
rect 106166 56006 106168 56058
rect 105922 56004 105928 56006
rect 105984 56004 106008 56006
rect 106064 56004 106088 56006
rect 106144 56004 106168 56006
rect 106224 56004 106230 56006
rect 105922 55995 106230 56004
rect 106658 55516 106966 55525
rect 106658 55514 106664 55516
rect 106720 55514 106744 55516
rect 106800 55514 106824 55516
rect 106880 55514 106904 55516
rect 106960 55514 106966 55516
rect 106720 55462 106722 55514
rect 106902 55462 106904 55514
rect 106658 55460 106664 55462
rect 106720 55460 106744 55462
rect 106800 55460 106824 55462
rect 106880 55460 106904 55462
rect 106960 55460 106966 55462
rect 106658 55451 106966 55460
rect 105922 54972 106230 54981
rect 105922 54970 105928 54972
rect 105984 54970 106008 54972
rect 106064 54970 106088 54972
rect 106144 54970 106168 54972
rect 106224 54970 106230 54972
rect 105984 54918 105986 54970
rect 106166 54918 106168 54970
rect 105922 54916 105928 54918
rect 105984 54916 106008 54918
rect 106064 54916 106088 54918
rect 106144 54916 106168 54918
rect 106224 54916 106230 54918
rect 105922 54907 106230 54916
rect 106658 54428 106966 54437
rect 106658 54426 106664 54428
rect 106720 54426 106744 54428
rect 106800 54426 106824 54428
rect 106880 54426 106904 54428
rect 106960 54426 106966 54428
rect 106720 54374 106722 54426
rect 106902 54374 106904 54426
rect 106658 54372 106664 54374
rect 106720 54372 106744 54374
rect 106800 54372 106824 54374
rect 106880 54372 106904 54374
rect 106960 54372 106966 54374
rect 106658 54363 106966 54372
rect 105922 53884 106230 53893
rect 105922 53882 105928 53884
rect 105984 53882 106008 53884
rect 106064 53882 106088 53884
rect 106144 53882 106168 53884
rect 106224 53882 106230 53884
rect 105984 53830 105986 53882
rect 106166 53830 106168 53882
rect 105922 53828 105928 53830
rect 105984 53828 106008 53830
rect 106064 53828 106088 53830
rect 106144 53828 106168 53830
rect 106224 53828 106230 53830
rect 105922 53819 106230 53828
rect 106658 53340 106966 53349
rect 106658 53338 106664 53340
rect 106720 53338 106744 53340
rect 106800 53338 106824 53340
rect 106880 53338 106904 53340
rect 106960 53338 106966 53340
rect 106720 53286 106722 53338
rect 106902 53286 106904 53338
rect 106658 53284 106664 53286
rect 106720 53284 106744 53286
rect 106800 53284 106824 53286
rect 106880 53284 106904 53286
rect 106960 53284 106966 53286
rect 106658 53275 106966 53284
rect 105922 52796 106230 52805
rect 105922 52794 105928 52796
rect 105984 52794 106008 52796
rect 106064 52794 106088 52796
rect 106144 52794 106168 52796
rect 106224 52794 106230 52796
rect 105984 52742 105986 52794
rect 106166 52742 106168 52794
rect 105922 52740 105928 52742
rect 105984 52740 106008 52742
rect 106064 52740 106088 52742
rect 106144 52740 106168 52742
rect 106224 52740 106230 52742
rect 105922 52731 106230 52740
rect 106658 52252 106966 52261
rect 106658 52250 106664 52252
rect 106720 52250 106744 52252
rect 106800 52250 106824 52252
rect 106880 52250 106904 52252
rect 106960 52250 106966 52252
rect 106720 52198 106722 52250
rect 106902 52198 106904 52250
rect 106658 52196 106664 52198
rect 106720 52196 106744 52198
rect 106800 52196 106824 52198
rect 106880 52196 106904 52198
rect 106960 52196 106966 52198
rect 106658 52187 106966 52196
rect 105922 51708 106230 51717
rect 105922 51706 105928 51708
rect 105984 51706 106008 51708
rect 106064 51706 106088 51708
rect 106144 51706 106168 51708
rect 106224 51706 106230 51708
rect 105984 51654 105986 51706
rect 106166 51654 106168 51706
rect 105922 51652 105928 51654
rect 105984 51652 106008 51654
rect 106064 51652 106088 51654
rect 106144 51652 106168 51654
rect 106224 51652 106230 51654
rect 105922 51643 106230 51652
rect 106658 51164 106966 51173
rect 106658 51162 106664 51164
rect 106720 51162 106744 51164
rect 106800 51162 106824 51164
rect 106880 51162 106904 51164
rect 106960 51162 106966 51164
rect 106720 51110 106722 51162
rect 106902 51110 106904 51162
rect 106658 51108 106664 51110
rect 106720 51108 106744 51110
rect 106800 51108 106824 51110
rect 106880 51108 106904 51110
rect 106960 51108 106966 51110
rect 106658 51099 106966 51108
rect 105922 50620 106230 50629
rect 105922 50618 105928 50620
rect 105984 50618 106008 50620
rect 106064 50618 106088 50620
rect 106144 50618 106168 50620
rect 106224 50618 106230 50620
rect 105984 50566 105986 50618
rect 106166 50566 106168 50618
rect 105922 50564 105928 50566
rect 105984 50564 106008 50566
rect 106064 50564 106088 50566
rect 106144 50564 106168 50566
rect 106224 50564 106230 50566
rect 105922 50555 106230 50564
rect 106658 50076 106966 50085
rect 106658 50074 106664 50076
rect 106720 50074 106744 50076
rect 106800 50074 106824 50076
rect 106880 50074 106904 50076
rect 106960 50074 106966 50076
rect 106720 50022 106722 50074
rect 106902 50022 106904 50074
rect 106658 50020 106664 50022
rect 106720 50020 106744 50022
rect 106800 50020 106824 50022
rect 106880 50020 106904 50022
rect 106960 50020 106966 50022
rect 106658 50011 106966 50020
rect 105922 49532 106230 49541
rect 105922 49530 105928 49532
rect 105984 49530 106008 49532
rect 106064 49530 106088 49532
rect 106144 49530 106168 49532
rect 106224 49530 106230 49532
rect 105984 49478 105986 49530
rect 106166 49478 106168 49530
rect 105922 49476 105928 49478
rect 105984 49476 106008 49478
rect 106064 49476 106088 49478
rect 106144 49476 106168 49478
rect 106224 49476 106230 49478
rect 105922 49467 106230 49476
rect 106658 48988 106966 48997
rect 106658 48986 106664 48988
rect 106720 48986 106744 48988
rect 106800 48986 106824 48988
rect 106880 48986 106904 48988
rect 106960 48986 106966 48988
rect 106720 48934 106722 48986
rect 106902 48934 106904 48986
rect 106658 48932 106664 48934
rect 106720 48932 106744 48934
rect 106800 48932 106824 48934
rect 106880 48932 106904 48934
rect 106960 48932 106966 48934
rect 106658 48923 106966 48932
rect 105922 48444 106230 48453
rect 105922 48442 105928 48444
rect 105984 48442 106008 48444
rect 106064 48442 106088 48444
rect 106144 48442 106168 48444
rect 106224 48442 106230 48444
rect 105984 48390 105986 48442
rect 106166 48390 106168 48442
rect 105922 48388 105928 48390
rect 105984 48388 106008 48390
rect 106064 48388 106088 48390
rect 106144 48388 106168 48390
rect 106224 48388 106230 48390
rect 105922 48379 106230 48388
rect 106658 47900 106966 47909
rect 106658 47898 106664 47900
rect 106720 47898 106744 47900
rect 106800 47898 106824 47900
rect 106880 47898 106904 47900
rect 106960 47898 106966 47900
rect 106720 47846 106722 47898
rect 106902 47846 106904 47898
rect 106658 47844 106664 47846
rect 106720 47844 106744 47846
rect 106800 47844 106824 47846
rect 106880 47844 106904 47846
rect 106960 47844 106966 47846
rect 106658 47835 106966 47844
rect 105922 47356 106230 47365
rect 105922 47354 105928 47356
rect 105984 47354 106008 47356
rect 106064 47354 106088 47356
rect 106144 47354 106168 47356
rect 106224 47354 106230 47356
rect 105984 47302 105986 47354
rect 106166 47302 106168 47354
rect 105922 47300 105928 47302
rect 105984 47300 106008 47302
rect 106064 47300 106088 47302
rect 106144 47300 106168 47302
rect 106224 47300 106230 47302
rect 105922 47291 106230 47300
rect 106658 46812 106966 46821
rect 106658 46810 106664 46812
rect 106720 46810 106744 46812
rect 106800 46810 106824 46812
rect 106880 46810 106904 46812
rect 106960 46810 106966 46812
rect 106720 46758 106722 46810
rect 106902 46758 106904 46810
rect 106658 46756 106664 46758
rect 106720 46756 106744 46758
rect 106800 46756 106824 46758
rect 106880 46756 106904 46758
rect 106960 46756 106966 46758
rect 106658 46747 106966 46756
rect 105922 46268 106230 46277
rect 105922 46266 105928 46268
rect 105984 46266 106008 46268
rect 106064 46266 106088 46268
rect 106144 46266 106168 46268
rect 106224 46266 106230 46268
rect 105984 46214 105986 46266
rect 106166 46214 106168 46266
rect 105922 46212 105928 46214
rect 105984 46212 106008 46214
rect 106064 46212 106088 46214
rect 106144 46212 106168 46214
rect 106224 46212 106230 46214
rect 105922 46203 106230 46212
rect 106658 45724 106966 45733
rect 106658 45722 106664 45724
rect 106720 45722 106744 45724
rect 106800 45722 106824 45724
rect 106880 45722 106904 45724
rect 106960 45722 106966 45724
rect 106720 45670 106722 45722
rect 106902 45670 106904 45722
rect 106658 45668 106664 45670
rect 106720 45668 106744 45670
rect 106800 45668 106824 45670
rect 106880 45668 106904 45670
rect 106960 45668 106966 45670
rect 106658 45659 106966 45668
rect 105922 45180 106230 45189
rect 105922 45178 105928 45180
rect 105984 45178 106008 45180
rect 106064 45178 106088 45180
rect 106144 45178 106168 45180
rect 106224 45178 106230 45180
rect 105984 45126 105986 45178
rect 106166 45126 106168 45178
rect 105922 45124 105928 45126
rect 105984 45124 106008 45126
rect 106064 45124 106088 45126
rect 106144 45124 106168 45126
rect 106224 45124 106230 45126
rect 105922 45115 106230 45124
rect 106658 44636 106966 44645
rect 106658 44634 106664 44636
rect 106720 44634 106744 44636
rect 106800 44634 106824 44636
rect 106880 44634 106904 44636
rect 106960 44634 106966 44636
rect 106720 44582 106722 44634
rect 106902 44582 106904 44634
rect 106658 44580 106664 44582
rect 106720 44580 106744 44582
rect 106800 44580 106824 44582
rect 106880 44580 106904 44582
rect 106960 44580 106966 44582
rect 106658 44571 106966 44580
rect 105922 44092 106230 44101
rect 105922 44090 105928 44092
rect 105984 44090 106008 44092
rect 106064 44090 106088 44092
rect 106144 44090 106168 44092
rect 106224 44090 106230 44092
rect 105984 44038 105986 44090
rect 106166 44038 106168 44090
rect 105922 44036 105928 44038
rect 105984 44036 106008 44038
rect 106064 44036 106088 44038
rect 106144 44036 106168 44038
rect 106224 44036 106230 44038
rect 105922 44027 106230 44036
rect 106658 43548 106966 43557
rect 106658 43546 106664 43548
rect 106720 43546 106744 43548
rect 106800 43546 106824 43548
rect 106880 43546 106904 43548
rect 106960 43546 106966 43548
rect 106720 43494 106722 43546
rect 106902 43494 106904 43546
rect 106658 43492 106664 43494
rect 106720 43492 106744 43494
rect 106800 43492 106824 43494
rect 106880 43492 106904 43494
rect 106960 43492 106966 43494
rect 106658 43483 106966 43492
rect 105922 43004 106230 43013
rect 105922 43002 105928 43004
rect 105984 43002 106008 43004
rect 106064 43002 106088 43004
rect 106144 43002 106168 43004
rect 106224 43002 106230 43004
rect 105984 42950 105986 43002
rect 106166 42950 106168 43002
rect 105922 42948 105928 42950
rect 105984 42948 106008 42950
rect 106064 42948 106088 42950
rect 106144 42948 106168 42950
rect 106224 42948 106230 42950
rect 105922 42939 106230 42948
rect 106658 42460 106966 42469
rect 106658 42458 106664 42460
rect 106720 42458 106744 42460
rect 106800 42458 106824 42460
rect 106880 42458 106904 42460
rect 106960 42458 106966 42460
rect 106720 42406 106722 42458
rect 106902 42406 106904 42458
rect 106658 42404 106664 42406
rect 106720 42404 106744 42406
rect 106800 42404 106824 42406
rect 106880 42404 106904 42406
rect 106960 42404 106966 42406
rect 106658 42395 106966 42404
rect 105922 41916 106230 41925
rect 105922 41914 105928 41916
rect 105984 41914 106008 41916
rect 106064 41914 106088 41916
rect 106144 41914 106168 41916
rect 106224 41914 106230 41916
rect 105984 41862 105986 41914
rect 106166 41862 106168 41914
rect 105922 41860 105928 41862
rect 105984 41860 106008 41862
rect 106064 41860 106088 41862
rect 106144 41860 106168 41862
rect 106224 41860 106230 41862
rect 105922 41851 106230 41860
rect 106658 41372 106966 41381
rect 106658 41370 106664 41372
rect 106720 41370 106744 41372
rect 106800 41370 106824 41372
rect 106880 41370 106904 41372
rect 106960 41370 106966 41372
rect 106720 41318 106722 41370
rect 106902 41318 106904 41370
rect 106658 41316 106664 41318
rect 106720 41316 106744 41318
rect 106800 41316 106824 41318
rect 106880 41316 106904 41318
rect 106960 41316 106966 41318
rect 106658 41307 106966 41316
rect 105922 40828 106230 40837
rect 105922 40826 105928 40828
rect 105984 40826 106008 40828
rect 106064 40826 106088 40828
rect 106144 40826 106168 40828
rect 106224 40826 106230 40828
rect 105984 40774 105986 40826
rect 106166 40774 106168 40826
rect 105922 40772 105928 40774
rect 105984 40772 106008 40774
rect 106064 40772 106088 40774
rect 106144 40772 106168 40774
rect 106224 40772 106230 40774
rect 105922 40763 106230 40772
rect 106658 40284 106966 40293
rect 106658 40282 106664 40284
rect 106720 40282 106744 40284
rect 106800 40282 106824 40284
rect 106880 40282 106904 40284
rect 106960 40282 106966 40284
rect 106720 40230 106722 40282
rect 106902 40230 106904 40282
rect 106658 40228 106664 40230
rect 106720 40228 106744 40230
rect 106800 40228 106824 40230
rect 106880 40228 106904 40230
rect 106960 40228 106966 40230
rect 106658 40219 106966 40228
rect 105922 39740 106230 39749
rect 105922 39738 105928 39740
rect 105984 39738 106008 39740
rect 106064 39738 106088 39740
rect 106144 39738 106168 39740
rect 106224 39738 106230 39740
rect 105984 39686 105986 39738
rect 106166 39686 106168 39738
rect 105922 39684 105928 39686
rect 105984 39684 106008 39686
rect 106064 39684 106088 39686
rect 106144 39684 106168 39686
rect 106224 39684 106230 39686
rect 105922 39675 106230 39684
rect 106658 39196 106966 39205
rect 106658 39194 106664 39196
rect 106720 39194 106744 39196
rect 106800 39194 106824 39196
rect 106880 39194 106904 39196
rect 106960 39194 106966 39196
rect 106720 39142 106722 39194
rect 106902 39142 106904 39194
rect 106658 39140 106664 39142
rect 106720 39140 106744 39142
rect 106800 39140 106824 39142
rect 106880 39140 106904 39142
rect 106960 39140 106966 39142
rect 106658 39131 106966 39140
rect 105922 38652 106230 38661
rect 105922 38650 105928 38652
rect 105984 38650 106008 38652
rect 106064 38650 106088 38652
rect 106144 38650 106168 38652
rect 106224 38650 106230 38652
rect 105984 38598 105986 38650
rect 106166 38598 106168 38650
rect 105922 38596 105928 38598
rect 105984 38596 106008 38598
rect 106064 38596 106088 38598
rect 106144 38596 106168 38598
rect 106224 38596 106230 38598
rect 105922 38587 106230 38596
rect 106658 38108 106966 38117
rect 106658 38106 106664 38108
rect 106720 38106 106744 38108
rect 106800 38106 106824 38108
rect 106880 38106 106904 38108
rect 106960 38106 106966 38108
rect 106720 38054 106722 38106
rect 106902 38054 106904 38106
rect 106658 38052 106664 38054
rect 106720 38052 106744 38054
rect 106800 38052 106824 38054
rect 106880 38052 106904 38054
rect 106960 38052 106966 38054
rect 106658 38043 106966 38052
rect 105922 37564 106230 37573
rect 105922 37562 105928 37564
rect 105984 37562 106008 37564
rect 106064 37562 106088 37564
rect 106144 37562 106168 37564
rect 106224 37562 106230 37564
rect 105984 37510 105986 37562
rect 106166 37510 106168 37562
rect 105922 37508 105928 37510
rect 105984 37508 106008 37510
rect 106064 37508 106088 37510
rect 106144 37508 106168 37510
rect 106224 37508 106230 37510
rect 105922 37499 106230 37508
rect 106658 37020 106966 37029
rect 106658 37018 106664 37020
rect 106720 37018 106744 37020
rect 106800 37018 106824 37020
rect 106880 37018 106904 37020
rect 106960 37018 106966 37020
rect 106720 36966 106722 37018
rect 106902 36966 106904 37018
rect 106658 36964 106664 36966
rect 106720 36964 106744 36966
rect 106800 36964 106824 36966
rect 106880 36964 106904 36966
rect 106960 36964 106966 36966
rect 106658 36955 106966 36964
rect 105922 36476 106230 36485
rect 105922 36474 105928 36476
rect 105984 36474 106008 36476
rect 106064 36474 106088 36476
rect 106144 36474 106168 36476
rect 106224 36474 106230 36476
rect 105984 36422 105986 36474
rect 106166 36422 106168 36474
rect 105922 36420 105928 36422
rect 105984 36420 106008 36422
rect 106064 36420 106088 36422
rect 106144 36420 106168 36422
rect 106224 36420 106230 36422
rect 105922 36411 106230 36420
rect 106658 35932 106966 35941
rect 106658 35930 106664 35932
rect 106720 35930 106744 35932
rect 106800 35930 106824 35932
rect 106880 35930 106904 35932
rect 106960 35930 106966 35932
rect 106720 35878 106722 35930
rect 106902 35878 106904 35930
rect 106658 35876 106664 35878
rect 106720 35876 106744 35878
rect 106800 35876 106824 35878
rect 106880 35876 106904 35878
rect 106960 35876 106966 35878
rect 106658 35867 106966 35876
rect 105922 35388 106230 35397
rect 105922 35386 105928 35388
rect 105984 35386 106008 35388
rect 106064 35386 106088 35388
rect 106144 35386 106168 35388
rect 106224 35386 106230 35388
rect 105984 35334 105986 35386
rect 106166 35334 106168 35386
rect 105922 35332 105928 35334
rect 105984 35332 106008 35334
rect 106064 35332 106088 35334
rect 106144 35332 106168 35334
rect 106224 35332 106230 35334
rect 105922 35323 106230 35332
rect 106658 34844 106966 34853
rect 106658 34842 106664 34844
rect 106720 34842 106744 34844
rect 106800 34842 106824 34844
rect 106880 34842 106904 34844
rect 106960 34842 106966 34844
rect 106720 34790 106722 34842
rect 106902 34790 106904 34842
rect 106658 34788 106664 34790
rect 106720 34788 106744 34790
rect 106800 34788 106824 34790
rect 106880 34788 106904 34790
rect 106960 34788 106966 34790
rect 106658 34779 106966 34788
rect 105922 34300 106230 34309
rect 105922 34298 105928 34300
rect 105984 34298 106008 34300
rect 106064 34298 106088 34300
rect 106144 34298 106168 34300
rect 106224 34298 106230 34300
rect 105984 34246 105986 34298
rect 106166 34246 106168 34298
rect 105922 34244 105928 34246
rect 105984 34244 106008 34246
rect 106064 34244 106088 34246
rect 106144 34244 106168 34246
rect 106224 34244 106230 34246
rect 105922 34235 106230 34244
rect 106658 33756 106966 33765
rect 106658 33754 106664 33756
rect 106720 33754 106744 33756
rect 106800 33754 106824 33756
rect 106880 33754 106904 33756
rect 106960 33754 106966 33756
rect 106720 33702 106722 33754
rect 106902 33702 106904 33754
rect 106658 33700 106664 33702
rect 106720 33700 106744 33702
rect 106800 33700 106824 33702
rect 106880 33700 106904 33702
rect 106960 33700 106966 33702
rect 106658 33691 106966 33700
rect 105922 33212 106230 33221
rect 105922 33210 105928 33212
rect 105984 33210 106008 33212
rect 106064 33210 106088 33212
rect 106144 33210 106168 33212
rect 106224 33210 106230 33212
rect 105984 33158 105986 33210
rect 106166 33158 106168 33210
rect 105922 33156 105928 33158
rect 105984 33156 106008 33158
rect 106064 33156 106088 33158
rect 106144 33156 106168 33158
rect 106224 33156 106230 33158
rect 105922 33147 106230 33156
rect 106658 32668 106966 32677
rect 106658 32666 106664 32668
rect 106720 32666 106744 32668
rect 106800 32666 106824 32668
rect 106880 32666 106904 32668
rect 106960 32666 106966 32668
rect 106720 32614 106722 32666
rect 106902 32614 106904 32666
rect 106658 32612 106664 32614
rect 106720 32612 106744 32614
rect 106800 32612 106824 32614
rect 106880 32612 106904 32614
rect 106960 32612 106966 32614
rect 106658 32603 106966 32612
rect 105922 32124 106230 32133
rect 105922 32122 105928 32124
rect 105984 32122 106008 32124
rect 106064 32122 106088 32124
rect 106144 32122 106168 32124
rect 106224 32122 106230 32124
rect 105984 32070 105986 32122
rect 106166 32070 106168 32122
rect 105922 32068 105928 32070
rect 105984 32068 106008 32070
rect 106064 32068 106088 32070
rect 106144 32068 106168 32070
rect 106224 32068 106230 32070
rect 105922 32059 106230 32068
rect 106658 31580 106966 31589
rect 106658 31578 106664 31580
rect 106720 31578 106744 31580
rect 106800 31578 106824 31580
rect 106880 31578 106904 31580
rect 106960 31578 106966 31580
rect 106720 31526 106722 31578
rect 106902 31526 106904 31578
rect 106658 31524 106664 31526
rect 106720 31524 106744 31526
rect 106800 31524 106824 31526
rect 106880 31524 106904 31526
rect 106960 31524 106966 31526
rect 106658 31515 106966 31524
rect 105922 31036 106230 31045
rect 105922 31034 105928 31036
rect 105984 31034 106008 31036
rect 106064 31034 106088 31036
rect 106144 31034 106168 31036
rect 106224 31034 106230 31036
rect 105984 30982 105986 31034
rect 106166 30982 106168 31034
rect 105922 30980 105928 30982
rect 105984 30980 106008 30982
rect 106064 30980 106088 30982
rect 106144 30980 106168 30982
rect 106224 30980 106230 30982
rect 105922 30971 106230 30980
rect 106658 30492 106966 30501
rect 106658 30490 106664 30492
rect 106720 30490 106744 30492
rect 106800 30490 106824 30492
rect 106880 30490 106904 30492
rect 106960 30490 106966 30492
rect 106720 30438 106722 30490
rect 106902 30438 106904 30490
rect 106658 30436 106664 30438
rect 106720 30436 106744 30438
rect 106800 30436 106824 30438
rect 106880 30436 106904 30438
rect 106960 30436 106966 30438
rect 106658 30427 106966 30436
rect 105922 29948 106230 29957
rect 105922 29946 105928 29948
rect 105984 29946 106008 29948
rect 106064 29946 106088 29948
rect 106144 29946 106168 29948
rect 106224 29946 106230 29948
rect 105984 29894 105986 29946
rect 106166 29894 106168 29946
rect 105922 29892 105928 29894
rect 105984 29892 106008 29894
rect 106064 29892 106088 29894
rect 106144 29892 106168 29894
rect 106224 29892 106230 29894
rect 105922 29883 106230 29892
rect 106658 29404 106966 29413
rect 106658 29402 106664 29404
rect 106720 29402 106744 29404
rect 106800 29402 106824 29404
rect 106880 29402 106904 29404
rect 106960 29402 106966 29404
rect 106720 29350 106722 29402
rect 106902 29350 106904 29402
rect 106658 29348 106664 29350
rect 106720 29348 106744 29350
rect 106800 29348 106824 29350
rect 106880 29348 106904 29350
rect 106960 29348 106966 29350
rect 106658 29339 106966 29348
rect 105922 28860 106230 28869
rect 105922 28858 105928 28860
rect 105984 28858 106008 28860
rect 106064 28858 106088 28860
rect 106144 28858 106168 28860
rect 106224 28858 106230 28860
rect 105984 28806 105986 28858
rect 106166 28806 106168 28858
rect 105922 28804 105928 28806
rect 105984 28804 106008 28806
rect 106064 28804 106088 28806
rect 106144 28804 106168 28806
rect 106224 28804 106230 28806
rect 105922 28795 106230 28804
rect 106658 28316 106966 28325
rect 106658 28314 106664 28316
rect 106720 28314 106744 28316
rect 106800 28314 106824 28316
rect 106880 28314 106904 28316
rect 106960 28314 106966 28316
rect 106720 28262 106722 28314
rect 106902 28262 106904 28314
rect 106658 28260 106664 28262
rect 106720 28260 106744 28262
rect 106800 28260 106824 28262
rect 106880 28260 106904 28262
rect 106960 28260 106966 28262
rect 106658 28251 106966 28260
rect 105922 27772 106230 27781
rect 105922 27770 105928 27772
rect 105984 27770 106008 27772
rect 106064 27770 106088 27772
rect 106144 27770 106168 27772
rect 106224 27770 106230 27772
rect 105984 27718 105986 27770
rect 106166 27718 106168 27770
rect 105922 27716 105928 27718
rect 105984 27716 106008 27718
rect 106064 27716 106088 27718
rect 106144 27716 106168 27718
rect 106224 27716 106230 27718
rect 105922 27707 106230 27716
rect 106658 27228 106966 27237
rect 106658 27226 106664 27228
rect 106720 27226 106744 27228
rect 106800 27226 106824 27228
rect 106880 27226 106904 27228
rect 106960 27226 106966 27228
rect 106720 27174 106722 27226
rect 106902 27174 106904 27226
rect 106658 27172 106664 27174
rect 106720 27172 106744 27174
rect 106800 27172 106824 27174
rect 106880 27172 106904 27174
rect 106960 27172 106966 27174
rect 106658 27163 106966 27172
rect 105922 26684 106230 26693
rect 105922 26682 105928 26684
rect 105984 26682 106008 26684
rect 106064 26682 106088 26684
rect 106144 26682 106168 26684
rect 106224 26682 106230 26684
rect 105984 26630 105986 26682
rect 106166 26630 106168 26682
rect 105922 26628 105928 26630
rect 105984 26628 106008 26630
rect 106064 26628 106088 26630
rect 106144 26628 106168 26630
rect 106224 26628 106230 26630
rect 105922 26619 106230 26628
rect 106658 26140 106966 26149
rect 106658 26138 106664 26140
rect 106720 26138 106744 26140
rect 106800 26138 106824 26140
rect 106880 26138 106904 26140
rect 106960 26138 106966 26140
rect 106720 26086 106722 26138
rect 106902 26086 106904 26138
rect 106658 26084 106664 26086
rect 106720 26084 106744 26086
rect 106800 26084 106824 26086
rect 106880 26084 106904 26086
rect 106960 26084 106966 26086
rect 106658 26075 106966 26084
rect 105922 25596 106230 25605
rect 105922 25594 105928 25596
rect 105984 25594 106008 25596
rect 106064 25594 106088 25596
rect 106144 25594 106168 25596
rect 106224 25594 106230 25596
rect 105984 25542 105986 25594
rect 106166 25542 106168 25594
rect 105922 25540 105928 25542
rect 105984 25540 106008 25542
rect 106064 25540 106088 25542
rect 106144 25540 106168 25542
rect 106224 25540 106230 25542
rect 105922 25531 106230 25540
rect 106658 25052 106966 25061
rect 106658 25050 106664 25052
rect 106720 25050 106744 25052
rect 106800 25050 106824 25052
rect 106880 25050 106904 25052
rect 106960 25050 106966 25052
rect 106720 24998 106722 25050
rect 106902 24998 106904 25050
rect 106658 24996 106664 24998
rect 106720 24996 106744 24998
rect 106800 24996 106824 24998
rect 106880 24996 106904 24998
rect 106960 24996 106966 24998
rect 106658 24987 106966 24996
rect 105922 24508 106230 24517
rect 105922 24506 105928 24508
rect 105984 24506 106008 24508
rect 106064 24506 106088 24508
rect 106144 24506 106168 24508
rect 106224 24506 106230 24508
rect 105984 24454 105986 24506
rect 106166 24454 106168 24506
rect 105922 24452 105928 24454
rect 105984 24452 106008 24454
rect 106064 24452 106088 24454
rect 106144 24452 106168 24454
rect 106224 24452 106230 24454
rect 105922 24443 106230 24452
rect 106658 23964 106966 23973
rect 106658 23962 106664 23964
rect 106720 23962 106744 23964
rect 106800 23962 106824 23964
rect 106880 23962 106904 23964
rect 106960 23962 106966 23964
rect 106720 23910 106722 23962
rect 106902 23910 106904 23962
rect 106658 23908 106664 23910
rect 106720 23908 106744 23910
rect 106800 23908 106824 23910
rect 106880 23908 106904 23910
rect 106960 23908 106966 23910
rect 106658 23899 106966 23908
rect 105922 23420 106230 23429
rect 105922 23418 105928 23420
rect 105984 23418 106008 23420
rect 106064 23418 106088 23420
rect 106144 23418 106168 23420
rect 106224 23418 106230 23420
rect 105984 23366 105986 23418
rect 106166 23366 106168 23418
rect 105922 23364 105928 23366
rect 105984 23364 106008 23366
rect 106064 23364 106088 23366
rect 106144 23364 106168 23366
rect 106224 23364 106230 23366
rect 105922 23355 106230 23364
rect 106658 22876 106966 22885
rect 106658 22874 106664 22876
rect 106720 22874 106744 22876
rect 106800 22874 106824 22876
rect 106880 22874 106904 22876
rect 106960 22874 106966 22876
rect 106720 22822 106722 22874
rect 106902 22822 106904 22874
rect 106658 22820 106664 22822
rect 106720 22820 106744 22822
rect 106800 22820 106824 22822
rect 106880 22820 106904 22822
rect 106960 22820 106966 22822
rect 106658 22811 106966 22820
rect 105922 22332 106230 22341
rect 105922 22330 105928 22332
rect 105984 22330 106008 22332
rect 106064 22330 106088 22332
rect 106144 22330 106168 22332
rect 106224 22330 106230 22332
rect 105984 22278 105986 22330
rect 106166 22278 106168 22330
rect 105922 22276 105928 22278
rect 105984 22276 106008 22278
rect 106064 22276 106088 22278
rect 106144 22276 106168 22278
rect 106224 22276 106230 22278
rect 105922 22267 106230 22276
rect 106658 21788 106966 21797
rect 106658 21786 106664 21788
rect 106720 21786 106744 21788
rect 106800 21786 106824 21788
rect 106880 21786 106904 21788
rect 106960 21786 106966 21788
rect 106720 21734 106722 21786
rect 106902 21734 106904 21786
rect 106658 21732 106664 21734
rect 106720 21732 106744 21734
rect 106800 21732 106824 21734
rect 106880 21732 106904 21734
rect 106960 21732 106966 21734
rect 106658 21723 106966 21732
rect 105922 21244 106230 21253
rect 105922 21242 105928 21244
rect 105984 21242 106008 21244
rect 106064 21242 106088 21244
rect 106144 21242 106168 21244
rect 106224 21242 106230 21244
rect 105984 21190 105986 21242
rect 106166 21190 106168 21242
rect 105922 21188 105928 21190
rect 105984 21188 106008 21190
rect 106064 21188 106088 21190
rect 106144 21188 106168 21190
rect 106224 21188 106230 21190
rect 105922 21179 106230 21188
rect 106658 20700 106966 20709
rect 106658 20698 106664 20700
rect 106720 20698 106744 20700
rect 106800 20698 106824 20700
rect 106880 20698 106904 20700
rect 106960 20698 106966 20700
rect 106720 20646 106722 20698
rect 106902 20646 106904 20698
rect 106658 20644 106664 20646
rect 106720 20644 106744 20646
rect 106800 20644 106824 20646
rect 106880 20644 106904 20646
rect 106960 20644 106966 20646
rect 106658 20635 106966 20644
rect 105922 20156 106230 20165
rect 105922 20154 105928 20156
rect 105984 20154 106008 20156
rect 106064 20154 106088 20156
rect 106144 20154 106168 20156
rect 106224 20154 106230 20156
rect 105984 20102 105986 20154
rect 106166 20102 106168 20154
rect 105922 20100 105928 20102
rect 105984 20100 106008 20102
rect 106064 20100 106088 20102
rect 106144 20100 106168 20102
rect 106224 20100 106230 20102
rect 105922 20091 106230 20100
rect 106658 19612 106966 19621
rect 106658 19610 106664 19612
rect 106720 19610 106744 19612
rect 106800 19610 106824 19612
rect 106880 19610 106904 19612
rect 106960 19610 106966 19612
rect 106720 19558 106722 19610
rect 106902 19558 106904 19610
rect 106658 19556 106664 19558
rect 106720 19556 106744 19558
rect 106800 19556 106824 19558
rect 106880 19556 106904 19558
rect 106960 19556 106966 19558
rect 106658 19547 106966 19556
rect 105922 19068 106230 19077
rect 105922 19066 105928 19068
rect 105984 19066 106008 19068
rect 106064 19066 106088 19068
rect 106144 19066 106168 19068
rect 106224 19066 106230 19068
rect 105984 19014 105986 19066
rect 106166 19014 106168 19066
rect 105922 19012 105928 19014
rect 105984 19012 106008 19014
rect 106064 19012 106088 19014
rect 106144 19012 106168 19014
rect 106224 19012 106230 19014
rect 105922 19003 106230 19012
rect 106658 18524 106966 18533
rect 106658 18522 106664 18524
rect 106720 18522 106744 18524
rect 106800 18522 106824 18524
rect 106880 18522 106904 18524
rect 106960 18522 106966 18524
rect 106720 18470 106722 18522
rect 106902 18470 106904 18522
rect 106658 18468 106664 18470
rect 106720 18468 106744 18470
rect 106800 18468 106824 18470
rect 106880 18468 106904 18470
rect 106960 18468 106966 18470
rect 106658 18459 106966 18468
rect 105922 17980 106230 17989
rect 105922 17978 105928 17980
rect 105984 17978 106008 17980
rect 106064 17978 106088 17980
rect 106144 17978 106168 17980
rect 106224 17978 106230 17980
rect 105984 17926 105986 17978
rect 106166 17926 106168 17978
rect 105922 17924 105928 17926
rect 105984 17924 106008 17926
rect 106064 17924 106088 17926
rect 106144 17924 106168 17926
rect 106224 17924 106230 17926
rect 105922 17915 106230 17924
rect 106658 17436 106966 17445
rect 106658 17434 106664 17436
rect 106720 17434 106744 17436
rect 106800 17434 106824 17436
rect 106880 17434 106904 17436
rect 106960 17434 106966 17436
rect 106720 17382 106722 17434
rect 106902 17382 106904 17434
rect 106658 17380 106664 17382
rect 106720 17380 106744 17382
rect 106800 17380 106824 17382
rect 106880 17380 106904 17382
rect 106960 17380 106966 17382
rect 106658 17371 106966 17380
rect 105922 16892 106230 16901
rect 105922 16890 105928 16892
rect 105984 16890 106008 16892
rect 106064 16890 106088 16892
rect 106144 16890 106168 16892
rect 106224 16890 106230 16892
rect 105984 16838 105986 16890
rect 106166 16838 106168 16890
rect 105922 16836 105928 16838
rect 105984 16836 106008 16838
rect 106064 16836 106088 16838
rect 106144 16836 106168 16838
rect 106224 16836 106230 16838
rect 105922 16827 106230 16836
rect 106658 16348 106966 16357
rect 106658 16346 106664 16348
rect 106720 16346 106744 16348
rect 106800 16346 106824 16348
rect 106880 16346 106904 16348
rect 106960 16346 106966 16348
rect 106720 16294 106722 16346
rect 106902 16294 106904 16346
rect 106658 16292 106664 16294
rect 106720 16292 106744 16294
rect 106800 16292 106824 16294
rect 106880 16292 106904 16294
rect 106960 16292 106966 16294
rect 106658 16283 106966 16292
rect 105922 15804 106230 15813
rect 105922 15802 105928 15804
rect 105984 15802 106008 15804
rect 106064 15802 106088 15804
rect 106144 15802 106168 15804
rect 106224 15802 106230 15804
rect 105984 15750 105986 15802
rect 106166 15750 106168 15802
rect 105922 15748 105928 15750
rect 105984 15748 106008 15750
rect 106064 15748 106088 15750
rect 106144 15748 106168 15750
rect 106224 15748 106230 15750
rect 105922 15739 106230 15748
rect 106658 15260 106966 15269
rect 106658 15258 106664 15260
rect 106720 15258 106744 15260
rect 106800 15258 106824 15260
rect 106880 15258 106904 15260
rect 106960 15258 106966 15260
rect 106720 15206 106722 15258
rect 106902 15206 106904 15258
rect 106658 15204 106664 15206
rect 106720 15204 106744 15206
rect 106800 15204 106824 15206
rect 106880 15204 106904 15206
rect 106960 15204 106966 15206
rect 106658 15195 106966 15204
rect 105922 14716 106230 14725
rect 105922 14714 105928 14716
rect 105984 14714 106008 14716
rect 106064 14714 106088 14716
rect 106144 14714 106168 14716
rect 106224 14714 106230 14716
rect 105984 14662 105986 14714
rect 106166 14662 106168 14714
rect 105922 14660 105928 14662
rect 105984 14660 106008 14662
rect 106064 14660 106088 14662
rect 106144 14660 106168 14662
rect 106224 14660 106230 14662
rect 105922 14651 106230 14660
rect 106658 14172 106966 14181
rect 106658 14170 106664 14172
rect 106720 14170 106744 14172
rect 106800 14170 106824 14172
rect 106880 14170 106904 14172
rect 106960 14170 106966 14172
rect 106720 14118 106722 14170
rect 106902 14118 106904 14170
rect 106658 14116 106664 14118
rect 106720 14116 106744 14118
rect 106800 14116 106824 14118
rect 106880 14116 106904 14118
rect 106960 14116 106966 14118
rect 106658 14107 106966 14116
rect 105922 13628 106230 13637
rect 105922 13626 105928 13628
rect 105984 13626 106008 13628
rect 106064 13626 106088 13628
rect 106144 13626 106168 13628
rect 106224 13626 106230 13628
rect 105984 13574 105986 13626
rect 106166 13574 106168 13626
rect 105922 13572 105928 13574
rect 105984 13572 106008 13574
rect 106064 13572 106088 13574
rect 106144 13572 106168 13574
rect 106224 13572 106230 13574
rect 105922 13563 106230 13572
rect 106658 13084 106966 13093
rect 106658 13082 106664 13084
rect 106720 13082 106744 13084
rect 106800 13082 106824 13084
rect 106880 13082 106904 13084
rect 106960 13082 106966 13084
rect 106720 13030 106722 13082
rect 106902 13030 106904 13082
rect 106658 13028 106664 13030
rect 106720 13028 106744 13030
rect 106800 13028 106824 13030
rect 106880 13028 106904 13030
rect 106960 13028 106966 13030
rect 106658 13019 106966 13028
rect 105922 12540 106230 12549
rect 105922 12538 105928 12540
rect 105984 12538 106008 12540
rect 106064 12538 106088 12540
rect 106144 12538 106168 12540
rect 106224 12538 106230 12540
rect 105984 12486 105986 12538
rect 106166 12486 106168 12538
rect 105922 12484 105928 12486
rect 105984 12484 106008 12486
rect 106064 12484 106088 12486
rect 106144 12484 106168 12486
rect 106224 12484 106230 12486
rect 105922 12475 106230 12484
rect 106658 11996 106966 12005
rect 106658 11994 106664 11996
rect 106720 11994 106744 11996
rect 106800 11994 106824 11996
rect 106880 11994 106904 11996
rect 106960 11994 106966 11996
rect 106720 11942 106722 11994
rect 106902 11942 106904 11994
rect 106658 11940 106664 11942
rect 106720 11940 106744 11942
rect 106800 11940 106824 11942
rect 106880 11940 106904 11942
rect 106960 11940 106966 11942
rect 106658 11931 106966 11940
rect 105922 11452 106230 11461
rect 105922 11450 105928 11452
rect 105984 11450 106008 11452
rect 106064 11450 106088 11452
rect 106144 11450 106168 11452
rect 106224 11450 106230 11452
rect 105984 11398 105986 11450
rect 106166 11398 106168 11450
rect 105922 11396 105928 11398
rect 105984 11396 106008 11398
rect 106064 11396 106088 11398
rect 106144 11396 106168 11398
rect 106224 11396 106230 11398
rect 105922 11387 106230 11396
rect 106658 10908 106966 10917
rect 106658 10906 106664 10908
rect 106720 10906 106744 10908
rect 106800 10906 106824 10908
rect 106880 10906 106904 10908
rect 106960 10906 106966 10908
rect 106720 10854 106722 10906
rect 106902 10854 106904 10906
rect 106658 10852 106664 10854
rect 106720 10852 106744 10854
rect 106800 10852 106824 10854
rect 106880 10852 106904 10854
rect 106960 10852 106966 10854
rect 106658 10843 106966 10852
rect 105922 10364 106230 10373
rect 105922 10362 105928 10364
rect 105984 10362 106008 10364
rect 106064 10362 106088 10364
rect 106144 10362 106168 10364
rect 106224 10362 106230 10364
rect 105984 10310 105986 10362
rect 106166 10310 106168 10362
rect 105922 10308 105928 10310
rect 105984 10308 106008 10310
rect 106064 10308 106088 10310
rect 106144 10308 106168 10310
rect 106224 10308 106230 10310
rect 105922 10299 106230 10308
rect 106658 9820 106966 9829
rect 106658 9818 106664 9820
rect 106720 9818 106744 9820
rect 106800 9818 106824 9820
rect 106880 9818 106904 9820
rect 106960 9818 106966 9820
rect 106720 9766 106722 9818
rect 106902 9766 106904 9818
rect 106658 9764 106664 9766
rect 106720 9764 106744 9766
rect 106800 9764 106824 9766
rect 106880 9764 106904 9766
rect 106960 9764 106966 9766
rect 106658 9755 106966 9764
rect 105922 9276 106230 9285
rect 105922 9274 105928 9276
rect 105984 9274 106008 9276
rect 106064 9274 106088 9276
rect 106144 9274 106168 9276
rect 106224 9274 106230 9276
rect 105984 9222 105986 9274
rect 106166 9222 106168 9274
rect 105922 9220 105928 9222
rect 105984 9220 106008 9222
rect 106064 9220 106088 9222
rect 106144 9220 106168 9222
rect 106224 9220 106230 9222
rect 105922 9211 106230 9220
rect 103980 9104 104032 9110
rect 103980 9046 104032 9052
rect 103704 9036 103756 9042
rect 103704 8978 103756 8984
rect 103612 8968 103664 8974
rect 103612 8910 103664 8916
rect 106658 8732 106966 8741
rect 106658 8730 106664 8732
rect 106720 8730 106744 8732
rect 106800 8730 106824 8732
rect 106880 8730 106904 8732
rect 106960 8730 106966 8732
rect 106720 8678 106722 8730
rect 106902 8678 106904 8730
rect 106658 8676 106664 8678
rect 106720 8676 106744 8678
rect 106800 8676 106824 8678
rect 106880 8676 106904 8678
rect 106960 8676 106966 8678
rect 106658 8667 106966 8676
rect 105922 8188 106230 8197
rect 105922 8186 105928 8188
rect 105984 8186 106008 8188
rect 106064 8186 106088 8188
rect 106144 8186 106168 8188
rect 106224 8186 106230 8188
rect 105984 8134 105986 8186
rect 106166 8134 106168 8186
rect 105922 8132 105928 8134
rect 105984 8132 106008 8134
rect 106064 8132 106088 8134
rect 106144 8132 106168 8134
rect 106224 8132 106230 8134
rect 105922 8123 106230 8132
rect 97034 7644 97342 7653
rect 97034 7642 97040 7644
rect 97096 7642 97120 7644
rect 97176 7642 97200 7644
rect 97256 7642 97280 7644
rect 97336 7642 97342 7644
rect 97096 7590 97098 7642
rect 97278 7590 97280 7642
rect 97034 7588 97040 7590
rect 97096 7588 97120 7590
rect 97176 7588 97200 7590
rect 97256 7588 97280 7590
rect 97336 7588 97342 7590
rect 97034 7579 97342 7588
rect 106658 7644 106966 7653
rect 106658 7642 106664 7644
rect 106720 7642 106744 7644
rect 106800 7642 106824 7644
rect 106880 7642 106904 7644
rect 106960 7642 106966 7644
rect 106720 7590 106722 7642
rect 106902 7590 106904 7642
rect 106658 7588 106664 7590
rect 106720 7588 106744 7590
rect 106800 7588 106824 7590
rect 106880 7588 106904 7590
rect 106960 7588 106966 7590
rect 106658 7579 106966 7588
rect 90548 7540 90600 7546
rect 90548 7482 90600 7488
rect 90640 7540 90692 7546
rect 90640 7482 90692 7488
rect 90824 7540 90876 7546
rect 90824 7482 90876 7488
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 96374 7100 96682 7109
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7035 96682 7044
rect 105922 7100 106230 7109
rect 105922 7098 105928 7100
rect 105984 7098 106008 7100
rect 106064 7098 106088 7100
rect 106144 7098 106168 7100
rect 106224 7098 106230 7100
rect 105984 7046 105986 7098
rect 106166 7046 106168 7098
rect 105922 7044 105928 7046
rect 105984 7044 106008 7046
rect 106064 7044 106088 7046
rect 106144 7044 106168 7046
rect 106224 7044 106230 7046
rect 105922 7035 106230 7044
rect 66314 6556 66622 6565
rect 66314 6554 66320 6556
rect 66376 6554 66400 6556
rect 66456 6554 66480 6556
rect 66536 6554 66560 6556
rect 66616 6554 66622 6556
rect 66376 6502 66378 6554
rect 66558 6502 66560 6554
rect 66314 6500 66320 6502
rect 66376 6500 66400 6502
rect 66456 6500 66480 6502
rect 66536 6500 66560 6502
rect 66616 6500 66622 6502
rect 66314 6491 66622 6500
rect 97034 6556 97342 6565
rect 97034 6554 97040 6556
rect 97096 6554 97120 6556
rect 97176 6554 97200 6556
rect 97256 6554 97280 6556
rect 97336 6554 97342 6556
rect 97096 6502 97098 6554
rect 97278 6502 97280 6554
rect 97034 6500 97040 6502
rect 97096 6500 97120 6502
rect 97176 6500 97200 6502
rect 97256 6500 97280 6502
rect 97336 6500 97342 6502
rect 97034 6491 97342 6500
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 96374 6012 96682 6021
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5947 96682 5956
rect 66314 5468 66622 5477
rect 66314 5466 66320 5468
rect 66376 5466 66400 5468
rect 66456 5466 66480 5468
rect 66536 5466 66560 5468
rect 66616 5466 66622 5468
rect 66376 5414 66378 5466
rect 66558 5414 66560 5466
rect 66314 5412 66320 5414
rect 66376 5412 66400 5414
rect 66456 5412 66480 5414
rect 66536 5412 66560 5414
rect 66616 5412 66622 5414
rect 66314 5403 66622 5412
rect 97034 5468 97342 5477
rect 97034 5466 97040 5468
rect 97096 5466 97120 5468
rect 97176 5466 97200 5468
rect 97256 5466 97280 5468
rect 97336 5466 97342 5468
rect 97096 5414 97098 5466
rect 97278 5414 97280 5466
rect 97034 5412 97040 5414
rect 97096 5412 97120 5414
rect 97176 5412 97200 5414
rect 97256 5412 97280 5414
rect 97336 5412 97342 5414
rect 97034 5403 97342 5412
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 96374 4924 96682 4933
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4859 96682 4868
rect 66314 4380 66622 4389
rect 66314 4378 66320 4380
rect 66376 4378 66400 4380
rect 66456 4378 66480 4380
rect 66536 4378 66560 4380
rect 66616 4378 66622 4380
rect 66376 4326 66378 4378
rect 66558 4326 66560 4378
rect 66314 4324 66320 4326
rect 66376 4324 66400 4326
rect 66456 4324 66480 4326
rect 66536 4324 66560 4326
rect 66616 4324 66622 4326
rect 66314 4315 66622 4324
rect 97034 4380 97342 4389
rect 97034 4378 97040 4380
rect 97096 4378 97120 4380
rect 97176 4378 97200 4380
rect 97256 4378 97280 4380
rect 97336 4378 97342 4380
rect 97096 4326 97098 4378
rect 97278 4326 97280 4378
rect 97034 4324 97040 4326
rect 97096 4324 97120 4326
rect 97176 4324 97200 4326
rect 97256 4324 97280 4326
rect 97336 4324 97342 4326
rect 97034 4315 97342 4324
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 96374 3836 96682 3845
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3771 96682 3780
rect 66314 3292 66622 3301
rect 66314 3290 66320 3292
rect 66376 3290 66400 3292
rect 66456 3290 66480 3292
rect 66536 3290 66560 3292
rect 66616 3290 66622 3292
rect 66376 3238 66378 3290
rect 66558 3238 66560 3290
rect 66314 3236 66320 3238
rect 66376 3236 66400 3238
rect 66456 3236 66480 3238
rect 66536 3236 66560 3238
rect 66616 3236 66622 3238
rect 66314 3227 66622 3236
rect 97034 3292 97342 3301
rect 97034 3290 97040 3292
rect 97096 3290 97120 3292
rect 97176 3290 97200 3292
rect 97256 3290 97280 3292
rect 97336 3290 97342 3292
rect 97096 3238 97098 3290
rect 97278 3238 97280 3290
rect 97034 3236 97040 3238
rect 97096 3236 97120 3238
rect 97176 3236 97200 3238
rect 97256 3236 97280 3238
rect 97336 3236 97342 3238
rect 97034 3227 97342 3236
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 96374 2748 96682 2757
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2683 96682 2692
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 32956 2644 33008 2650
rect 32956 2586 33008 2592
rect 34244 2644 34296 2650
rect 34244 2586 34296 2592
rect 35440 2644 35492 2650
rect 35440 2586 35492 2592
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 38752 2644 38804 2650
rect 38752 2586 38804 2592
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 41328 2644 41380 2650
rect 41328 2586 41380 2592
rect 42156 2644 42208 2650
rect 42156 2586 42208 2592
rect 43444 2644 43496 2650
rect 43444 2586 43496 2592
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 39948 2304 40000 2310
rect 39948 2246 40000 2252
rect 41236 2304 41288 2310
rect 41236 2246 41288 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 31588 800 31616 2246
rect 32876 800 32904 2246
rect 34164 800 34192 2246
rect 35452 800 35480 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36096 800 36124 2246
rect 37384 800 37412 2246
rect 38672 800 38700 2246
rect 39960 800 39988 2246
rect 41248 800 41276 2246
rect 41892 800 41920 2246
rect 43180 800 43208 2246
rect 66314 2204 66622 2213
rect 66314 2202 66320 2204
rect 66376 2202 66400 2204
rect 66456 2202 66480 2204
rect 66536 2202 66560 2204
rect 66616 2202 66622 2204
rect 66376 2150 66378 2202
rect 66558 2150 66560 2202
rect 66314 2148 66320 2150
rect 66376 2148 66400 2150
rect 66456 2148 66480 2150
rect 66536 2148 66560 2150
rect 66616 2148 66622 2150
rect 66314 2139 66622 2148
rect 97034 2204 97342 2213
rect 97034 2202 97040 2204
rect 97096 2202 97120 2204
rect 97176 2202 97200 2204
rect 97256 2202 97280 2204
rect 97336 2202 97342 2204
rect 97096 2150 97098 2202
rect 97278 2150 97280 2202
rect 97034 2148 97040 2150
rect 97096 2148 97120 2150
rect 97176 2148 97200 2150
rect 97256 2148 97280 2150
rect 97336 2148 97342 2150
rect 97034 2139 97342 2148
rect 16118 0 16174 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 43166 0 43222 800
<< via2 >>
rect 4220 147450 4276 147452
rect 4300 147450 4356 147452
rect 4380 147450 4436 147452
rect 4460 147450 4516 147452
rect 4220 147398 4266 147450
rect 4266 147398 4276 147450
rect 4300 147398 4330 147450
rect 4330 147398 4342 147450
rect 4342 147398 4356 147450
rect 4380 147398 4394 147450
rect 4394 147398 4406 147450
rect 4406 147398 4436 147450
rect 4460 147398 4470 147450
rect 4470 147398 4516 147450
rect 4220 147396 4276 147398
rect 4300 147396 4356 147398
rect 4380 147396 4436 147398
rect 4460 147396 4516 147398
rect 34940 147450 34996 147452
rect 35020 147450 35076 147452
rect 35100 147450 35156 147452
rect 35180 147450 35236 147452
rect 34940 147398 34986 147450
rect 34986 147398 34996 147450
rect 35020 147398 35050 147450
rect 35050 147398 35062 147450
rect 35062 147398 35076 147450
rect 35100 147398 35114 147450
rect 35114 147398 35126 147450
rect 35126 147398 35156 147450
rect 35180 147398 35190 147450
rect 35190 147398 35236 147450
rect 34940 147396 34996 147398
rect 35020 147396 35076 147398
rect 35100 147396 35156 147398
rect 35180 147396 35236 147398
rect 65660 147450 65716 147452
rect 65740 147450 65796 147452
rect 65820 147450 65876 147452
rect 65900 147450 65956 147452
rect 65660 147398 65706 147450
rect 65706 147398 65716 147450
rect 65740 147398 65770 147450
rect 65770 147398 65782 147450
rect 65782 147398 65796 147450
rect 65820 147398 65834 147450
rect 65834 147398 65846 147450
rect 65846 147398 65876 147450
rect 65900 147398 65910 147450
rect 65910 147398 65956 147450
rect 65660 147396 65716 147398
rect 65740 147396 65796 147398
rect 65820 147396 65876 147398
rect 65900 147396 65956 147398
rect 96380 147450 96436 147452
rect 96460 147450 96516 147452
rect 96540 147450 96596 147452
rect 96620 147450 96676 147452
rect 96380 147398 96426 147450
rect 96426 147398 96436 147450
rect 96460 147398 96490 147450
rect 96490 147398 96502 147450
rect 96502 147398 96516 147450
rect 96540 147398 96554 147450
rect 96554 147398 96566 147450
rect 96566 147398 96596 147450
rect 96620 147398 96630 147450
rect 96630 147398 96676 147450
rect 96380 147396 96436 147398
rect 96460 147396 96516 147398
rect 96540 147396 96596 147398
rect 96620 147396 96676 147398
rect 4880 146906 4936 146908
rect 4960 146906 5016 146908
rect 5040 146906 5096 146908
rect 5120 146906 5176 146908
rect 4880 146854 4926 146906
rect 4926 146854 4936 146906
rect 4960 146854 4990 146906
rect 4990 146854 5002 146906
rect 5002 146854 5016 146906
rect 5040 146854 5054 146906
rect 5054 146854 5066 146906
rect 5066 146854 5096 146906
rect 5120 146854 5130 146906
rect 5130 146854 5176 146906
rect 4880 146852 4936 146854
rect 4960 146852 5016 146854
rect 5040 146852 5096 146854
rect 5120 146852 5176 146854
rect 35600 146906 35656 146908
rect 35680 146906 35736 146908
rect 35760 146906 35816 146908
rect 35840 146906 35896 146908
rect 35600 146854 35646 146906
rect 35646 146854 35656 146906
rect 35680 146854 35710 146906
rect 35710 146854 35722 146906
rect 35722 146854 35736 146906
rect 35760 146854 35774 146906
rect 35774 146854 35786 146906
rect 35786 146854 35816 146906
rect 35840 146854 35850 146906
rect 35850 146854 35896 146906
rect 35600 146852 35656 146854
rect 35680 146852 35736 146854
rect 35760 146852 35816 146854
rect 35840 146852 35896 146854
rect 66320 146906 66376 146908
rect 66400 146906 66456 146908
rect 66480 146906 66536 146908
rect 66560 146906 66616 146908
rect 66320 146854 66366 146906
rect 66366 146854 66376 146906
rect 66400 146854 66430 146906
rect 66430 146854 66442 146906
rect 66442 146854 66456 146906
rect 66480 146854 66494 146906
rect 66494 146854 66506 146906
rect 66506 146854 66536 146906
rect 66560 146854 66570 146906
rect 66570 146854 66616 146906
rect 66320 146852 66376 146854
rect 66400 146852 66456 146854
rect 66480 146852 66536 146854
rect 66560 146852 66616 146854
rect 97040 146906 97096 146908
rect 97120 146906 97176 146908
rect 97200 146906 97256 146908
rect 97280 146906 97336 146908
rect 97040 146854 97086 146906
rect 97086 146854 97096 146906
rect 97120 146854 97150 146906
rect 97150 146854 97162 146906
rect 97162 146854 97176 146906
rect 97200 146854 97214 146906
rect 97214 146854 97226 146906
rect 97226 146854 97256 146906
rect 97280 146854 97290 146906
rect 97290 146854 97336 146906
rect 97040 146852 97096 146854
rect 97120 146852 97176 146854
rect 97200 146852 97256 146854
rect 97280 146852 97336 146854
rect 4220 146362 4276 146364
rect 4300 146362 4356 146364
rect 4380 146362 4436 146364
rect 4460 146362 4516 146364
rect 4220 146310 4266 146362
rect 4266 146310 4276 146362
rect 4300 146310 4330 146362
rect 4330 146310 4342 146362
rect 4342 146310 4356 146362
rect 4380 146310 4394 146362
rect 4394 146310 4406 146362
rect 4406 146310 4436 146362
rect 4460 146310 4470 146362
rect 4470 146310 4516 146362
rect 4220 146308 4276 146310
rect 4300 146308 4356 146310
rect 4380 146308 4436 146310
rect 4460 146308 4516 146310
rect 34940 146362 34996 146364
rect 35020 146362 35076 146364
rect 35100 146362 35156 146364
rect 35180 146362 35236 146364
rect 34940 146310 34986 146362
rect 34986 146310 34996 146362
rect 35020 146310 35050 146362
rect 35050 146310 35062 146362
rect 35062 146310 35076 146362
rect 35100 146310 35114 146362
rect 35114 146310 35126 146362
rect 35126 146310 35156 146362
rect 35180 146310 35190 146362
rect 35190 146310 35236 146362
rect 34940 146308 34996 146310
rect 35020 146308 35076 146310
rect 35100 146308 35156 146310
rect 35180 146308 35236 146310
rect 65660 146362 65716 146364
rect 65740 146362 65796 146364
rect 65820 146362 65876 146364
rect 65900 146362 65956 146364
rect 65660 146310 65706 146362
rect 65706 146310 65716 146362
rect 65740 146310 65770 146362
rect 65770 146310 65782 146362
rect 65782 146310 65796 146362
rect 65820 146310 65834 146362
rect 65834 146310 65846 146362
rect 65846 146310 65876 146362
rect 65900 146310 65910 146362
rect 65910 146310 65956 146362
rect 65660 146308 65716 146310
rect 65740 146308 65796 146310
rect 65820 146308 65876 146310
rect 65900 146308 65956 146310
rect 96380 146362 96436 146364
rect 96460 146362 96516 146364
rect 96540 146362 96596 146364
rect 96620 146362 96676 146364
rect 96380 146310 96426 146362
rect 96426 146310 96436 146362
rect 96460 146310 96490 146362
rect 96490 146310 96502 146362
rect 96502 146310 96516 146362
rect 96540 146310 96554 146362
rect 96554 146310 96566 146362
rect 96566 146310 96596 146362
rect 96620 146310 96630 146362
rect 96630 146310 96676 146362
rect 96380 146308 96436 146310
rect 96460 146308 96516 146310
rect 96540 146308 96596 146310
rect 96620 146308 96676 146310
rect 4880 145818 4936 145820
rect 4960 145818 5016 145820
rect 5040 145818 5096 145820
rect 5120 145818 5176 145820
rect 4880 145766 4926 145818
rect 4926 145766 4936 145818
rect 4960 145766 4990 145818
rect 4990 145766 5002 145818
rect 5002 145766 5016 145818
rect 5040 145766 5054 145818
rect 5054 145766 5066 145818
rect 5066 145766 5096 145818
rect 5120 145766 5130 145818
rect 5130 145766 5176 145818
rect 4880 145764 4936 145766
rect 4960 145764 5016 145766
rect 5040 145764 5096 145766
rect 5120 145764 5176 145766
rect 35600 145818 35656 145820
rect 35680 145818 35736 145820
rect 35760 145818 35816 145820
rect 35840 145818 35896 145820
rect 35600 145766 35646 145818
rect 35646 145766 35656 145818
rect 35680 145766 35710 145818
rect 35710 145766 35722 145818
rect 35722 145766 35736 145818
rect 35760 145766 35774 145818
rect 35774 145766 35786 145818
rect 35786 145766 35816 145818
rect 35840 145766 35850 145818
rect 35850 145766 35896 145818
rect 35600 145764 35656 145766
rect 35680 145764 35736 145766
rect 35760 145764 35816 145766
rect 35840 145764 35896 145766
rect 66320 145818 66376 145820
rect 66400 145818 66456 145820
rect 66480 145818 66536 145820
rect 66560 145818 66616 145820
rect 66320 145766 66366 145818
rect 66366 145766 66376 145818
rect 66400 145766 66430 145818
rect 66430 145766 66442 145818
rect 66442 145766 66456 145818
rect 66480 145766 66494 145818
rect 66494 145766 66506 145818
rect 66506 145766 66536 145818
rect 66560 145766 66570 145818
rect 66570 145766 66616 145818
rect 66320 145764 66376 145766
rect 66400 145764 66456 145766
rect 66480 145764 66536 145766
rect 66560 145764 66616 145766
rect 97040 145818 97096 145820
rect 97120 145818 97176 145820
rect 97200 145818 97256 145820
rect 97280 145818 97336 145820
rect 97040 145766 97086 145818
rect 97086 145766 97096 145818
rect 97120 145766 97150 145818
rect 97150 145766 97162 145818
rect 97162 145766 97176 145818
rect 97200 145766 97214 145818
rect 97214 145766 97226 145818
rect 97226 145766 97256 145818
rect 97280 145766 97290 145818
rect 97290 145766 97336 145818
rect 97040 145764 97096 145766
rect 97120 145764 97176 145766
rect 97200 145764 97256 145766
rect 97280 145764 97336 145766
rect 4220 145274 4276 145276
rect 4300 145274 4356 145276
rect 4380 145274 4436 145276
rect 4460 145274 4516 145276
rect 4220 145222 4266 145274
rect 4266 145222 4276 145274
rect 4300 145222 4330 145274
rect 4330 145222 4342 145274
rect 4342 145222 4356 145274
rect 4380 145222 4394 145274
rect 4394 145222 4406 145274
rect 4406 145222 4436 145274
rect 4460 145222 4470 145274
rect 4470 145222 4516 145274
rect 4220 145220 4276 145222
rect 4300 145220 4356 145222
rect 4380 145220 4436 145222
rect 4460 145220 4516 145222
rect 34940 145274 34996 145276
rect 35020 145274 35076 145276
rect 35100 145274 35156 145276
rect 35180 145274 35236 145276
rect 34940 145222 34986 145274
rect 34986 145222 34996 145274
rect 35020 145222 35050 145274
rect 35050 145222 35062 145274
rect 35062 145222 35076 145274
rect 35100 145222 35114 145274
rect 35114 145222 35126 145274
rect 35126 145222 35156 145274
rect 35180 145222 35190 145274
rect 35190 145222 35236 145274
rect 34940 145220 34996 145222
rect 35020 145220 35076 145222
rect 35100 145220 35156 145222
rect 35180 145220 35236 145222
rect 65660 145274 65716 145276
rect 65740 145274 65796 145276
rect 65820 145274 65876 145276
rect 65900 145274 65956 145276
rect 65660 145222 65706 145274
rect 65706 145222 65716 145274
rect 65740 145222 65770 145274
rect 65770 145222 65782 145274
rect 65782 145222 65796 145274
rect 65820 145222 65834 145274
rect 65834 145222 65846 145274
rect 65846 145222 65876 145274
rect 65900 145222 65910 145274
rect 65910 145222 65956 145274
rect 65660 145220 65716 145222
rect 65740 145220 65796 145222
rect 65820 145220 65876 145222
rect 65900 145220 65956 145222
rect 96380 145274 96436 145276
rect 96460 145274 96516 145276
rect 96540 145274 96596 145276
rect 96620 145274 96676 145276
rect 96380 145222 96426 145274
rect 96426 145222 96436 145274
rect 96460 145222 96490 145274
rect 96490 145222 96502 145274
rect 96502 145222 96516 145274
rect 96540 145222 96554 145274
rect 96554 145222 96566 145274
rect 96566 145222 96596 145274
rect 96620 145222 96630 145274
rect 96630 145222 96676 145274
rect 96380 145220 96436 145222
rect 96460 145220 96516 145222
rect 96540 145220 96596 145222
rect 96620 145220 96676 145222
rect 4880 144730 4936 144732
rect 4960 144730 5016 144732
rect 5040 144730 5096 144732
rect 5120 144730 5176 144732
rect 4880 144678 4926 144730
rect 4926 144678 4936 144730
rect 4960 144678 4990 144730
rect 4990 144678 5002 144730
rect 5002 144678 5016 144730
rect 5040 144678 5054 144730
rect 5054 144678 5066 144730
rect 5066 144678 5096 144730
rect 5120 144678 5130 144730
rect 5130 144678 5176 144730
rect 4880 144676 4936 144678
rect 4960 144676 5016 144678
rect 5040 144676 5096 144678
rect 5120 144676 5176 144678
rect 35600 144730 35656 144732
rect 35680 144730 35736 144732
rect 35760 144730 35816 144732
rect 35840 144730 35896 144732
rect 35600 144678 35646 144730
rect 35646 144678 35656 144730
rect 35680 144678 35710 144730
rect 35710 144678 35722 144730
rect 35722 144678 35736 144730
rect 35760 144678 35774 144730
rect 35774 144678 35786 144730
rect 35786 144678 35816 144730
rect 35840 144678 35850 144730
rect 35850 144678 35896 144730
rect 35600 144676 35656 144678
rect 35680 144676 35736 144678
rect 35760 144676 35816 144678
rect 35840 144676 35896 144678
rect 66320 144730 66376 144732
rect 66400 144730 66456 144732
rect 66480 144730 66536 144732
rect 66560 144730 66616 144732
rect 66320 144678 66366 144730
rect 66366 144678 66376 144730
rect 66400 144678 66430 144730
rect 66430 144678 66442 144730
rect 66442 144678 66456 144730
rect 66480 144678 66494 144730
rect 66494 144678 66506 144730
rect 66506 144678 66536 144730
rect 66560 144678 66570 144730
rect 66570 144678 66616 144730
rect 66320 144676 66376 144678
rect 66400 144676 66456 144678
rect 66480 144676 66536 144678
rect 66560 144676 66616 144678
rect 97040 144730 97096 144732
rect 97120 144730 97176 144732
rect 97200 144730 97256 144732
rect 97280 144730 97336 144732
rect 97040 144678 97086 144730
rect 97086 144678 97096 144730
rect 97120 144678 97150 144730
rect 97150 144678 97162 144730
rect 97162 144678 97176 144730
rect 97200 144678 97214 144730
rect 97214 144678 97226 144730
rect 97226 144678 97256 144730
rect 97280 144678 97290 144730
rect 97290 144678 97336 144730
rect 97040 144676 97096 144678
rect 97120 144676 97176 144678
rect 97200 144676 97256 144678
rect 97280 144676 97336 144678
rect 4220 144186 4276 144188
rect 4300 144186 4356 144188
rect 4380 144186 4436 144188
rect 4460 144186 4516 144188
rect 4220 144134 4266 144186
rect 4266 144134 4276 144186
rect 4300 144134 4330 144186
rect 4330 144134 4342 144186
rect 4342 144134 4356 144186
rect 4380 144134 4394 144186
rect 4394 144134 4406 144186
rect 4406 144134 4436 144186
rect 4460 144134 4470 144186
rect 4470 144134 4516 144186
rect 4220 144132 4276 144134
rect 4300 144132 4356 144134
rect 4380 144132 4436 144134
rect 4460 144132 4516 144134
rect 34940 144186 34996 144188
rect 35020 144186 35076 144188
rect 35100 144186 35156 144188
rect 35180 144186 35236 144188
rect 34940 144134 34986 144186
rect 34986 144134 34996 144186
rect 35020 144134 35050 144186
rect 35050 144134 35062 144186
rect 35062 144134 35076 144186
rect 35100 144134 35114 144186
rect 35114 144134 35126 144186
rect 35126 144134 35156 144186
rect 35180 144134 35190 144186
rect 35190 144134 35236 144186
rect 34940 144132 34996 144134
rect 35020 144132 35076 144134
rect 35100 144132 35156 144134
rect 35180 144132 35236 144134
rect 65660 144186 65716 144188
rect 65740 144186 65796 144188
rect 65820 144186 65876 144188
rect 65900 144186 65956 144188
rect 65660 144134 65706 144186
rect 65706 144134 65716 144186
rect 65740 144134 65770 144186
rect 65770 144134 65782 144186
rect 65782 144134 65796 144186
rect 65820 144134 65834 144186
rect 65834 144134 65846 144186
rect 65846 144134 65876 144186
rect 65900 144134 65910 144186
rect 65910 144134 65956 144186
rect 65660 144132 65716 144134
rect 65740 144132 65796 144134
rect 65820 144132 65876 144134
rect 65900 144132 65956 144134
rect 96380 144186 96436 144188
rect 96460 144186 96516 144188
rect 96540 144186 96596 144188
rect 96620 144186 96676 144188
rect 96380 144134 96426 144186
rect 96426 144134 96436 144186
rect 96460 144134 96490 144186
rect 96490 144134 96502 144186
rect 96502 144134 96516 144186
rect 96540 144134 96554 144186
rect 96554 144134 96566 144186
rect 96566 144134 96596 144186
rect 96620 144134 96630 144186
rect 96630 144134 96676 144186
rect 96380 144132 96436 144134
rect 96460 144132 96516 144134
rect 96540 144132 96596 144134
rect 96620 144132 96676 144134
rect 4880 143642 4936 143644
rect 4960 143642 5016 143644
rect 5040 143642 5096 143644
rect 5120 143642 5176 143644
rect 4880 143590 4926 143642
rect 4926 143590 4936 143642
rect 4960 143590 4990 143642
rect 4990 143590 5002 143642
rect 5002 143590 5016 143642
rect 5040 143590 5054 143642
rect 5054 143590 5066 143642
rect 5066 143590 5096 143642
rect 5120 143590 5130 143642
rect 5130 143590 5176 143642
rect 4880 143588 4936 143590
rect 4960 143588 5016 143590
rect 5040 143588 5096 143590
rect 5120 143588 5176 143590
rect 35600 143642 35656 143644
rect 35680 143642 35736 143644
rect 35760 143642 35816 143644
rect 35840 143642 35896 143644
rect 35600 143590 35646 143642
rect 35646 143590 35656 143642
rect 35680 143590 35710 143642
rect 35710 143590 35722 143642
rect 35722 143590 35736 143642
rect 35760 143590 35774 143642
rect 35774 143590 35786 143642
rect 35786 143590 35816 143642
rect 35840 143590 35850 143642
rect 35850 143590 35896 143642
rect 35600 143588 35656 143590
rect 35680 143588 35736 143590
rect 35760 143588 35816 143590
rect 35840 143588 35896 143590
rect 66320 143642 66376 143644
rect 66400 143642 66456 143644
rect 66480 143642 66536 143644
rect 66560 143642 66616 143644
rect 66320 143590 66366 143642
rect 66366 143590 66376 143642
rect 66400 143590 66430 143642
rect 66430 143590 66442 143642
rect 66442 143590 66456 143642
rect 66480 143590 66494 143642
rect 66494 143590 66506 143642
rect 66506 143590 66536 143642
rect 66560 143590 66570 143642
rect 66570 143590 66616 143642
rect 66320 143588 66376 143590
rect 66400 143588 66456 143590
rect 66480 143588 66536 143590
rect 66560 143588 66616 143590
rect 97040 143642 97096 143644
rect 97120 143642 97176 143644
rect 97200 143642 97256 143644
rect 97280 143642 97336 143644
rect 97040 143590 97086 143642
rect 97086 143590 97096 143642
rect 97120 143590 97150 143642
rect 97150 143590 97162 143642
rect 97162 143590 97176 143642
rect 97200 143590 97214 143642
rect 97214 143590 97226 143642
rect 97226 143590 97256 143642
rect 97280 143590 97290 143642
rect 97290 143590 97336 143642
rect 97040 143588 97096 143590
rect 97120 143588 97176 143590
rect 97200 143588 97256 143590
rect 97280 143588 97336 143590
rect 4220 143098 4276 143100
rect 4300 143098 4356 143100
rect 4380 143098 4436 143100
rect 4460 143098 4516 143100
rect 4220 143046 4266 143098
rect 4266 143046 4276 143098
rect 4300 143046 4330 143098
rect 4330 143046 4342 143098
rect 4342 143046 4356 143098
rect 4380 143046 4394 143098
rect 4394 143046 4406 143098
rect 4406 143046 4436 143098
rect 4460 143046 4470 143098
rect 4470 143046 4516 143098
rect 4220 143044 4276 143046
rect 4300 143044 4356 143046
rect 4380 143044 4436 143046
rect 4460 143044 4516 143046
rect 34940 143098 34996 143100
rect 35020 143098 35076 143100
rect 35100 143098 35156 143100
rect 35180 143098 35236 143100
rect 34940 143046 34986 143098
rect 34986 143046 34996 143098
rect 35020 143046 35050 143098
rect 35050 143046 35062 143098
rect 35062 143046 35076 143098
rect 35100 143046 35114 143098
rect 35114 143046 35126 143098
rect 35126 143046 35156 143098
rect 35180 143046 35190 143098
rect 35190 143046 35236 143098
rect 34940 143044 34996 143046
rect 35020 143044 35076 143046
rect 35100 143044 35156 143046
rect 35180 143044 35236 143046
rect 65660 143098 65716 143100
rect 65740 143098 65796 143100
rect 65820 143098 65876 143100
rect 65900 143098 65956 143100
rect 65660 143046 65706 143098
rect 65706 143046 65716 143098
rect 65740 143046 65770 143098
rect 65770 143046 65782 143098
rect 65782 143046 65796 143098
rect 65820 143046 65834 143098
rect 65834 143046 65846 143098
rect 65846 143046 65876 143098
rect 65900 143046 65910 143098
rect 65910 143046 65956 143098
rect 65660 143044 65716 143046
rect 65740 143044 65796 143046
rect 65820 143044 65876 143046
rect 65900 143044 65956 143046
rect 96380 143098 96436 143100
rect 96460 143098 96516 143100
rect 96540 143098 96596 143100
rect 96620 143098 96676 143100
rect 96380 143046 96426 143098
rect 96426 143046 96436 143098
rect 96460 143046 96490 143098
rect 96490 143046 96502 143098
rect 96502 143046 96516 143098
rect 96540 143046 96554 143098
rect 96554 143046 96566 143098
rect 96566 143046 96596 143098
rect 96620 143046 96630 143098
rect 96630 143046 96676 143098
rect 96380 143044 96436 143046
rect 96460 143044 96516 143046
rect 96540 143044 96596 143046
rect 96620 143044 96676 143046
rect 4880 142554 4936 142556
rect 4960 142554 5016 142556
rect 5040 142554 5096 142556
rect 5120 142554 5176 142556
rect 4880 142502 4926 142554
rect 4926 142502 4936 142554
rect 4960 142502 4990 142554
rect 4990 142502 5002 142554
rect 5002 142502 5016 142554
rect 5040 142502 5054 142554
rect 5054 142502 5066 142554
rect 5066 142502 5096 142554
rect 5120 142502 5130 142554
rect 5130 142502 5176 142554
rect 4880 142500 4936 142502
rect 4960 142500 5016 142502
rect 5040 142500 5096 142502
rect 5120 142500 5176 142502
rect 35600 142554 35656 142556
rect 35680 142554 35736 142556
rect 35760 142554 35816 142556
rect 35840 142554 35896 142556
rect 35600 142502 35646 142554
rect 35646 142502 35656 142554
rect 35680 142502 35710 142554
rect 35710 142502 35722 142554
rect 35722 142502 35736 142554
rect 35760 142502 35774 142554
rect 35774 142502 35786 142554
rect 35786 142502 35816 142554
rect 35840 142502 35850 142554
rect 35850 142502 35896 142554
rect 35600 142500 35656 142502
rect 35680 142500 35736 142502
rect 35760 142500 35816 142502
rect 35840 142500 35896 142502
rect 66320 142554 66376 142556
rect 66400 142554 66456 142556
rect 66480 142554 66536 142556
rect 66560 142554 66616 142556
rect 66320 142502 66366 142554
rect 66366 142502 66376 142554
rect 66400 142502 66430 142554
rect 66430 142502 66442 142554
rect 66442 142502 66456 142554
rect 66480 142502 66494 142554
rect 66494 142502 66506 142554
rect 66506 142502 66536 142554
rect 66560 142502 66570 142554
rect 66570 142502 66616 142554
rect 66320 142500 66376 142502
rect 66400 142500 66456 142502
rect 66480 142500 66536 142502
rect 66560 142500 66616 142502
rect 97040 142554 97096 142556
rect 97120 142554 97176 142556
rect 97200 142554 97256 142556
rect 97280 142554 97336 142556
rect 97040 142502 97086 142554
rect 97086 142502 97096 142554
rect 97120 142502 97150 142554
rect 97150 142502 97162 142554
rect 97162 142502 97176 142554
rect 97200 142502 97214 142554
rect 97214 142502 97226 142554
rect 97226 142502 97256 142554
rect 97280 142502 97290 142554
rect 97290 142502 97336 142554
rect 97040 142500 97096 142502
rect 97120 142500 97176 142502
rect 97200 142500 97256 142502
rect 97280 142500 97336 142502
rect 4220 142010 4276 142012
rect 4300 142010 4356 142012
rect 4380 142010 4436 142012
rect 4460 142010 4516 142012
rect 4220 141958 4266 142010
rect 4266 141958 4276 142010
rect 4300 141958 4330 142010
rect 4330 141958 4342 142010
rect 4342 141958 4356 142010
rect 4380 141958 4394 142010
rect 4394 141958 4406 142010
rect 4406 141958 4436 142010
rect 4460 141958 4470 142010
rect 4470 141958 4516 142010
rect 4220 141956 4276 141958
rect 4300 141956 4356 141958
rect 4380 141956 4436 141958
rect 4460 141956 4516 141958
rect 34940 142010 34996 142012
rect 35020 142010 35076 142012
rect 35100 142010 35156 142012
rect 35180 142010 35236 142012
rect 34940 141958 34986 142010
rect 34986 141958 34996 142010
rect 35020 141958 35050 142010
rect 35050 141958 35062 142010
rect 35062 141958 35076 142010
rect 35100 141958 35114 142010
rect 35114 141958 35126 142010
rect 35126 141958 35156 142010
rect 35180 141958 35190 142010
rect 35190 141958 35236 142010
rect 34940 141956 34996 141958
rect 35020 141956 35076 141958
rect 35100 141956 35156 141958
rect 35180 141956 35236 141958
rect 65660 142010 65716 142012
rect 65740 142010 65796 142012
rect 65820 142010 65876 142012
rect 65900 142010 65956 142012
rect 65660 141958 65706 142010
rect 65706 141958 65716 142010
rect 65740 141958 65770 142010
rect 65770 141958 65782 142010
rect 65782 141958 65796 142010
rect 65820 141958 65834 142010
rect 65834 141958 65846 142010
rect 65846 141958 65876 142010
rect 65900 141958 65910 142010
rect 65910 141958 65956 142010
rect 65660 141956 65716 141958
rect 65740 141956 65796 141958
rect 65820 141956 65876 141958
rect 65900 141956 65956 141958
rect 96380 142010 96436 142012
rect 96460 142010 96516 142012
rect 96540 142010 96596 142012
rect 96620 142010 96676 142012
rect 96380 141958 96426 142010
rect 96426 141958 96436 142010
rect 96460 141958 96490 142010
rect 96490 141958 96502 142010
rect 96502 141958 96516 142010
rect 96540 141958 96554 142010
rect 96554 141958 96566 142010
rect 96566 141958 96596 142010
rect 96620 141958 96630 142010
rect 96630 141958 96676 142010
rect 96380 141956 96436 141958
rect 96460 141956 96516 141958
rect 96540 141956 96596 141958
rect 96620 141956 96676 141958
rect 4880 141466 4936 141468
rect 4960 141466 5016 141468
rect 5040 141466 5096 141468
rect 5120 141466 5176 141468
rect 4880 141414 4926 141466
rect 4926 141414 4936 141466
rect 4960 141414 4990 141466
rect 4990 141414 5002 141466
rect 5002 141414 5016 141466
rect 5040 141414 5054 141466
rect 5054 141414 5066 141466
rect 5066 141414 5096 141466
rect 5120 141414 5130 141466
rect 5130 141414 5176 141466
rect 4880 141412 4936 141414
rect 4960 141412 5016 141414
rect 5040 141412 5096 141414
rect 5120 141412 5176 141414
rect 35600 141466 35656 141468
rect 35680 141466 35736 141468
rect 35760 141466 35816 141468
rect 35840 141466 35896 141468
rect 35600 141414 35646 141466
rect 35646 141414 35656 141466
rect 35680 141414 35710 141466
rect 35710 141414 35722 141466
rect 35722 141414 35736 141466
rect 35760 141414 35774 141466
rect 35774 141414 35786 141466
rect 35786 141414 35816 141466
rect 35840 141414 35850 141466
rect 35850 141414 35896 141466
rect 35600 141412 35656 141414
rect 35680 141412 35736 141414
rect 35760 141412 35816 141414
rect 35840 141412 35896 141414
rect 66320 141466 66376 141468
rect 66400 141466 66456 141468
rect 66480 141466 66536 141468
rect 66560 141466 66616 141468
rect 66320 141414 66366 141466
rect 66366 141414 66376 141466
rect 66400 141414 66430 141466
rect 66430 141414 66442 141466
rect 66442 141414 66456 141466
rect 66480 141414 66494 141466
rect 66494 141414 66506 141466
rect 66506 141414 66536 141466
rect 66560 141414 66570 141466
rect 66570 141414 66616 141466
rect 66320 141412 66376 141414
rect 66400 141412 66456 141414
rect 66480 141412 66536 141414
rect 66560 141412 66616 141414
rect 97040 141466 97096 141468
rect 97120 141466 97176 141468
rect 97200 141466 97256 141468
rect 97280 141466 97336 141468
rect 97040 141414 97086 141466
rect 97086 141414 97096 141466
rect 97120 141414 97150 141466
rect 97150 141414 97162 141466
rect 97162 141414 97176 141466
rect 97200 141414 97214 141466
rect 97214 141414 97226 141466
rect 97226 141414 97256 141466
rect 97280 141414 97290 141466
rect 97290 141414 97336 141466
rect 97040 141412 97096 141414
rect 97120 141412 97176 141414
rect 97200 141412 97256 141414
rect 97280 141412 97336 141414
rect 4220 140922 4276 140924
rect 4300 140922 4356 140924
rect 4380 140922 4436 140924
rect 4460 140922 4516 140924
rect 4220 140870 4266 140922
rect 4266 140870 4276 140922
rect 4300 140870 4330 140922
rect 4330 140870 4342 140922
rect 4342 140870 4356 140922
rect 4380 140870 4394 140922
rect 4394 140870 4406 140922
rect 4406 140870 4436 140922
rect 4460 140870 4470 140922
rect 4470 140870 4516 140922
rect 4220 140868 4276 140870
rect 4300 140868 4356 140870
rect 4380 140868 4436 140870
rect 4460 140868 4516 140870
rect 34940 140922 34996 140924
rect 35020 140922 35076 140924
rect 35100 140922 35156 140924
rect 35180 140922 35236 140924
rect 34940 140870 34986 140922
rect 34986 140870 34996 140922
rect 35020 140870 35050 140922
rect 35050 140870 35062 140922
rect 35062 140870 35076 140922
rect 35100 140870 35114 140922
rect 35114 140870 35126 140922
rect 35126 140870 35156 140922
rect 35180 140870 35190 140922
rect 35190 140870 35236 140922
rect 34940 140868 34996 140870
rect 35020 140868 35076 140870
rect 35100 140868 35156 140870
rect 35180 140868 35236 140870
rect 65660 140922 65716 140924
rect 65740 140922 65796 140924
rect 65820 140922 65876 140924
rect 65900 140922 65956 140924
rect 65660 140870 65706 140922
rect 65706 140870 65716 140922
rect 65740 140870 65770 140922
rect 65770 140870 65782 140922
rect 65782 140870 65796 140922
rect 65820 140870 65834 140922
rect 65834 140870 65846 140922
rect 65846 140870 65876 140922
rect 65900 140870 65910 140922
rect 65910 140870 65956 140922
rect 65660 140868 65716 140870
rect 65740 140868 65796 140870
rect 65820 140868 65876 140870
rect 65900 140868 65956 140870
rect 96380 140922 96436 140924
rect 96460 140922 96516 140924
rect 96540 140922 96596 140924
rect 96620 140922 96676 140924
rect 96380 140870 96426 140922
rect 96426 140870 96436 140922
rect 96460 140870 96490 140922
rect 96490 140870 96502 140922
rect 96502 140870 96516 140922
rect 96540 140870 96554 140922
rect 96554 140870 96566 140922
rect 96566 140870 96596 140922
rect 96620 140870 96630 140922
rect 96630 140870 96676 140922
rect 96380 140868 96436 140870
rect 96460 140868 96516 140870
rect 96540 140868 96596 140870
rect 96620 140868 96676 140870
rect 4880 140378 4936 140380
rect 4960 140378 5016 140380
rect 5040 140378 5096 140380
rect 5120 140378 5176 140380
rect 4880 140326 4926 140378
rect 4926 140326 4936 140378
rect 4960 140326 4990 140378
rect 4990 140326 5002 140378
rect 5002 140326 5016 140378
rect 5040 140326 5054 140378
rect 5054 140326 5066 140378
rect 5066 140326 5096 140378
rect 5120 140326 5130 140378
rect 5130 140326 5176 140378
rect 4880 140324 4936 140326
rect 4960 140324 5016 140326
rect 5040 140324 5096 140326
rect 5120 140324 5176 140326
rect 35600 140378 35656 140380
rect 35680 140378 35736 140380
rect 35760 140378 35816 140380
rect 35840 140378 35896 140380
rect 35600 140326 35646 140378
rect 35646 140326 35656 140378
rect 35680 140326 35710 140378
rect 35710 140326 35722 140378
rect 35722 140326 35736 140378
rect 35760 140326 35774 140378
rect 35774 140326 35786 140378
rect 35786 140326 35816 140378
rect 35840 140326 35850 140378
rect 35850 140326 35896 140378
rect 35600 140324 35656 140326
rect 35680 140324 35736 140326
rect 35760 140324 35816 140326
rect 35840 140324 35896 140326
rect 66320 140378 66376 140380
rect 66400 140378 66456 140380
rect 66480 140378 66536 140380
rect 66560 140378 66616 140380
rect 66320 140326 66366 140378
rect 66366 140326 66376 140378
rect 66400 140326 66430 140378
rect 66430 140326 66442 140378
rect 66442 140326 66456 140378
rect 66480 140326 66494 140378
rect 66494 140326 66506 140378
rect 66506 140326 66536 140378
rect 66560 140326 66570 140378
rect 66570 140326 66616 140378
rect 66320 140324 66376 140326
rect 66400 140324 66456 140326
rect 66480 140324 66536 140326
rect 66560 140324 66616 140326
rect 97040 140378 97096 140380
rect 97120 140378 97176 140380
rect 97200 140378 97256 140380
rect 97280 140378 97336 140380
rect 97040 140326 97086 140378
rect 97086 140326 97096 140378
rect 97120 140326 97150 140378
rect 97150 140326 97162 140378
rect 97162 140326 97176 140378
rect 97200 140326 97214 140378
rect 97214 140326 97226 140378
rect 97226 140326 97256 140378
rect 97280 140326 97290 140378
rect 97290 140326 97336 140378
rect 97040 140324 97096 140326
rect 97120 140324 97176 140326
rect 97200 140324 97256 140326
rect 97280 140324 97336 140326
rect 4220 139834 4276 139836
rect 4300 139834 4356 139836
rect 4380 139834 4436 139836
rect 4460 139834 4516 139836
rect 4220 139782 4266 139834
rect 4266 139782 4276 139834
rect 4300 139782 4330 139834
rect 4330 139782 4342 139834
rect 4342 139782 4356 139834
rect 4380 139782 4394 139834
rect 4394 139782 4406 139834
rect 4406 139782 4436 139834
rect 4460 139782 4470 139834
rect 4470 139782 4516 139834
rect 4220 139780 4276 139782
rect 4300 139780 4356 139782
rect 4380 139780 4436 139782
rect 4460 139780 4516 139782
rect 34940 139834 34996 139836
rect 35020 139834 35076 139836
rect 35100 139834 35156 139836
rect 35180 139834 35236 139836
rect 34940 139782 34986 139834
rect 34986 139782 34996 139834
rect 35020 139782 35050 139834
rect 35050 139782 35062 139834
rect 35062 139782 35076 139834
rect 35100 139782 35114 139834
rect 35114 139782 35126 139834
rect 35126 139782 35156 139834
rect 35180 139782 35190 139834
rect 35190 139782 35236 139834
rect 34940 139780 34996 139782
rect 35020 139780 35076 139782
rect 35100 139780 35156 139782
rect 35180 139780 35236 139782
rect 65660 139834 65716 139836
rect 65740 139834 65796 139836
rect 65820 139834 65876 139836
rect 65900 139834 65956 139836
rect 65660 139782 65706 139834
rect 65706 139782 65716 139834
rect 65740 139782 65770 139834
rect 65770 139782 65782 139834
rect 65782 139782 65796 139834
rect 65820 139782 65834 139834
rect 65834 139782 65846 139834
rect 65846 139782 65876 139834
rect 65900 139782 65910 139834
rect 65910 139782 65956 139834
rect 65660 139780 65716 139782
rect 65740 139780 65796 139782
rect 65820 139780 65876 139782
rect 65900 139780 65956 139782
rect 96380 139834 96436 139836
rect 96460 139834 96516 139836
rect 96540 139834 96596 139836
rect 96620 139834 96676 139836
rect 96380 139782 96426 139834
rect 96426 139782 96436 139834
rect 96460 139782 96490 139834
rect 96490 139782 96502 139834
rect 96502 139782 96516 139834
rect 96540 139782 96554 139834
rect 96554 139782 96566 139834
rect 96566 139782 96596 139834
rect 96620 139782 96630 139834
rect 96630 139782 96676 139834
rect 96380 139780 96436 139782
rect 96460 139780 96516 139782
rect 96540 139780 96596 139782
rect 96620 139780 96676 139782
rect 4880 139290 4936 139292
rect 4960 139290 5016 139292
rect 5040 139290 5096 139292
rect 5120 139290 5176 139292
rect 4880 139238 4926 139290
rect 4926 139238 4936 139290
rect 4960 139238 4990 139290
rect 4990 139238 5002 139290
rect 5002 139238 5016 139290
rect 5040 139238 5054 139290
rect 5054 139238 5066 139290
rect 5066 139238 5096 139290
rect 5120 139238 5130 139290
rect 5130 139238 5176 139290
rect 4880 139236 4936 139238
rect 4960 139236 5016 139238
rect 5040 139236 5096 139238
rect 5120 139236 5176 139238
rect 35600 139290 35656 139292
rect 35680 139290 35736 139292
rect 35760 139290 35816 139292
rect 35840 139290 35896 139292
rect 35600 139238 35646 139290
rect 35646 139238 35656 139290
rect 35680 139238 35710 139290
rect 35710 139238 35722 139290
rect 35722 139238 35736 139290
rect 35760 139238 35774 139290
rect 35774 139238 35786 139290
rect 35786 139238 35816 139290
rect 35840 139238 35850 139290
rect 35850 139238 35896 139290
rect 35600 139236 35656 139238
rect 35680 139236 35736 139238
rect 35760 139236 35816 139238
rect 35840 139236 35896 139238
rect 66320 139290 66376 139292
rect 66400 139290 66456 139292
rect 66480 139290 66536 139292
rect 66560 139290 66616 139292
rect 66320 139238 66366 139290
rect 66366 139238 66376 139290
rect 66400 139238 66430 139290
rect 66430 139238 66442 139290
rect 66442 139238 66456 139290
rect 66480 139238 66494 139290
rect 66494 139238 66506 139290
rect 66506 139238 66536 139290
rect 66560 139238 66570 139290
rect 66570 139238 66616 139290
rect 66320 139236 66376 139238
rect 66400 139236 66456 139238
rect 66480 139236 66536 139238
rect 66560 139236 66616 139238
rect 97040 139290 97096 139292
rect 97120 139290 97176 139292
rect 97200 139290 97256 139292
rect 97280 139290 97336 139292
rect 97040 139238 97086 139290
rect 97086 139238 97096 139290
rect 97120 139238 97150 139290
rect 97150 139238 97162 139290
rect 97162 139238 97176 139290
rect 97200 139238 97214 139290
rect 97214 139238 97226 139290
rect 97226 139238 97256 139290
rect 97280 139238 97290 139290
rect 97290 139238 97336 139290
rect 97040 139236 97096 139238
rect 97120 139236 97176 139238
rect 97200 139236 97256 139238
rect 97280 139236 97336 139238
rect 4220 138746 4276 138748
rect 4300 138746 4356 138748
rect 4380 138746 4436 138748
rect 4460 138746 4516 138748
rect 4220 138694 4266 138746
rect 4266 138694 4276 138746
rect 4300 138694 4330 138746
rect 4330 138694 4342 138746
rect 4342 138694 4356 138746
rect 4380 138694 4394 138746
rect 4394 138694 4406 138746
rect 4406 138694 4436 138746
rect 4460 138694 4470 138746
rect 4470 138694 4516 138746
rect 4220 138692 4276 138694
rect 4300 138692 4356 138694
rect 4380 138692 4436 138694
rect 4460 138692 4516 138694
rect 34940 138746 34996 138748
rect 35020 138746 35076 138748
rect 35100 138746 35156 138748
rect 35180 138746 35236 138748
rect 34940 138694 34986 138746
rect 34986 138694 34996 138746
rect 35020 138694 35050 138746
rect 35050 138694 35062 138746
rect 35062 138694 35076 138746
rect 35100 138694 35114 138746
rect 35114 138694 35126 138746
rect 35126 138694 35156 138746
rect 35180 138694 35190 138746
rect 35190 138694 35236 138746
rect 34940 138692 34996 138694
rect 35020 138692 35076 138694
rect 35100 138692 35156 138694
rect 35180 138692 35236 138694
rect 65660 138746 65716 138748
rect 65740 138746 65796 138748
rect 65820 138746 65876 138748
rect 65900 138746 65956 138748
rect 65660 138694 65706 138746
rect 65706 138694 65716 138746
rect 65740 138694 65770 138746
rect 65770 138694 65782 138746
rect 65782 138694 65796 138746
rect 65820 138694 65834 138746
rect 65834 138694 65846 138746
rect 65846 138694 65876 138746
rect 65900 138694 65910 138746
rect 65910 138694 65956 138746
rect 65660 138692 65716 138694
rect 65740 138692 65796 138694
rect 65820 138692 65876 138694
rect 65900 138692 65956 138694
rect 96380 138746 96436 138748
rect 96460 138746 96516 138748
rect 96540 138746 96596 138748
rect 96620 138746 96676 138748
rect 96380 138694 96426 138746
rect 96426 138694 96436 138746
rect 96460 138694 96490 138746
rect 96490 138694 96502 138746
rect 96502 138694 96516 138746
rect 96540 138694 96554 138746
rect 96554 138694 96566 138746
rect 96566 138694 96596 138746
rect 96620 138694 96630 138746
rect 96630 138694 96676 138746
rect 96380 138692 96436 138694
rect 96460 138692 96516 138694
rect 96540 138692 96596 138694
rect 96620 138692 96676 138694
rect 4880 138202 4936 138204
rect 4960 138202 5016 138204
rect 5040 138202 5096 138204
rect 5120 138202 5176 138204
rect 4880 138150 4926 138202
rect 4926 138150 4936 138202
rect 4960 138150 4990 138202
rect 4990 138150 5002 138202
rect 5002 138150 5016 138202
rect 5040 138150 5054 138202
rect 5054 138150 5066 138202
rect 5066 138150 5096 138202
rect 5120 138150 5130 138202
rect 5130 138150 5176 138202
rect 4880 138148 4936 138150
rect 4960 138148 5016 138150
rect 5040 138148 5096 138150
rect 5120 138148 5176 138150
rect 35600 138202 35656 138204
rect 35680 138202 35736 138204
rect 35760 138202 35816 138204
rect 35840 138202 35896 138204
rect 35600 138150 35646 138202
rect 35646 138150 35656 138202
rect 35680 138150 35710 138202
rect 35710 138150 35722 138202
rect 35722 138150 35736 138202
rect 35760 138150 35774 138202
rect 35774 138150 35786 138202
rect 35786 138150 35816 138202
rect 35840 138150 35850 138202
rect 35850 138150 35896 138202
rect 35600 138148 35656 138150
rect 35680 138148 35736 138150
rect 35760 138148 35816 138150
rect 35840 138148 35896 138150
rect 66320 138202 66376 138204
rect 66400 138202 66456 138204
rect 66480 138202 66536 138204
rect 66560 138202 66616 138204
rect 66320 138150 66366 138202
rect 66366 138150 66376 138202
rect 66400 138150 66430 138202
rect 66430 138150 66442 138202
rect 66442 138150 66456 138202
rect 66480 138150 66494 138202
rect 66494 138150 66506 138202
rect 66506 138150 66536 138202
rect 66560 138150 66570 138202
rect 66570 138150 66616 138202
rect 66320 138148 66376 138150
rect 66400 138148 66456 138150
rect 66480 138148 66536 138150
rect 66560 138148 66616 138150
rect 97040 138202 97096 138204
rect 97120 138202 97176 138204
rect 97200 138202 97256 138204
rect 97280 138202 97336 138204
rect 97040 138150 97086 138202
rect 97086 138150 97096 138202
rect 97120 138150 97150 138202
rect 97150 138150 97162 138202
rect 97162 138150 97176 138202
rect 97200 138150 97214 138202
rect 97214 138150 97226 138202
rect 97226 138150 97256 138202
rect 97280 138150 97290 138202
rect 97290 138150 97336 138202
rect 97040 138148 97096 138150
rect 97120 138148 97176 138150
rect 97200 138148 97256 138150
rect 97280 138148 97336 138150
rect 4220 137658 4276 137660
rect 4300 137658 4356 137660
rect 4380 137658 4436 137660
rect 4460 137658 4516 137660
rect 4220 137606 4266 137658
rect 4266 137606 4276 137658
rect 4300 137606 4330 137658
rect 4330 137606 4342 137658
rect 4342 137606 4356 137658
rect 4380 137606 4394 137658
rect 4394 137606 4406 137658
rect 4406 137606 4436 137658
rect 4460 137606 4470 137658
rect 4470 137606 4516 137658
rect 4220 137604 4276 137606
rect 4300 137604 4356 137606
rect 4380 137604 4436 137606
rect 4460 137604 4516 137606
rect 34940 137658 34996 137660
rect 35020 137658 35076 137660
rect 35100 137658 35156 137660
rect 35180 137658 35236 137660
rect 34940 137606 34986 137658
rect 34986 137606 34996 137658
rect 35020 137606 35050 137658
rect 35050 137606 35062 137658
rect 35062 137606 35076 137658
rect 35100 137606 35114 137658
rect 35114 137606 35126 137658
rect 35126 137606 35156 137658
rect 35180 137606 35190 137658
rect 35190 137606 35236 137658
rect 34940 137604 34996 137606
rect 35020 137604 35076 137606
rect 35100 137604 35156 137606
rect 35180 137604 35236 137606
rect 65660 137658 65716 137660
rect 65740 137658 65796 137660
rect 65820 137658 65876 137660
rect 65900 137658 65956 137660
rect 65660 137606 65706 137658
rect 65706 137606 65716 137658
rect 65740 137606 65770 137658
rect 65770 137606 65782 137658
rect 65782 137606 65796 137658
rect 65820 137606 65834 137658
rect 65834 137606 65846 137658
rect 65846 137606 65876 137658
rect 65900 137606 65910 137658
rect 65910 137606 65956 137658
rect 65660 137604 65716 137606
rect 65740 137604 65796 137606
rect 65820 137604 65876 137606
rect 65900 137604 65956 137606
rect 96380 137658 96436 137660
rect 96460 137658 96516 137660
rect 96540 137658 96596 137660
rect 96620 137658 96676 137660
rect 96380 137606 96426 137658
rect 96426 137606 96436 137658
rect 96460 137606 96490 137658
rect 96490 137606 96502 137658
rect 96502 137606 96516 137658
rect 96540 137606 96554 137658
rect 96554 137606 96566 137658
rect 96566 137606 96596 137658
rect 96620 137606 96630 137658
rect 96630 137606 96676 137658
rect 96380 137604 96436 137606
rect 96460 137604 96516 137606
rect 96540 137604 96596 137606
rect 96620 137604 96676 137606
rect 4880 137114 4936 137116
rect 4960 137114 5016 137116
rect 5040 137114 5096 137116
rect 5120 137114 5176 137116
rect 4880 137062 4926 137114
rect 4926 137062 4936 137114
rect 4960 137062 4990 137114
rect 4990 137062 5002 137114
rect 5002 137062 5016 137114
rect 5040 137062 5054 137114
rect 5054 137062 5066 137114
rect 5066 137062 5096 137114
rect 5120 137062 5130 137114
rect 5130 137062 5176 137114
rect 4880 137060 4936 137062
rect 4960 137060 5016 137062
rect 5040 137060 5096 137062
rect 5120 137060 5176 137062
rect 35600 137114 35656 137116
rect 35680 137114 35736 137116
rect 35760 137114 35816 137116
rect 35840 137114 35896 137116
rect 35600 137062 35646 137114
rect 35646 137062 35656 137114
rect 35680 137062 35710 137114
rect 35710 137062 35722 137114
rect 35722 137062 35736 137114
rect 35760 137062 35774 137114
rect 35774 137062 35786 137114
rect 35786 137062 35816 137114
rect 35840 137062 35850 137114
rect 35850 137062 35896 137114
rect 35600 137060 35656 137062
rect 35680 137060 35736 137062
rect 35760 137060 35816 137062
rect 35840 137060 35896 137062
rect 66320 137114 66376 137116
rect 66400 137114 66456 137116
rect 66480 137114 66536 137116
rect 66560 137114 66616 137116
rect 66320 137062 66366 137114
rect 66366 137062 66376 137114
rect 66400 137062 66430 137114
rect 66430 137062 66442 137114
rect 66442 137062 66456 137114
rect 66480 137062 66494 137114
rect 66494 137062 66506 137114
rect 66506 137062 66536 137114
rect 66560 137062 66570 137114
rect 66570 137062 66616 137114
rect 66320 137060 66376 137062
rect 66400 137060 66456 137062
rect 66480 137060 66536 137062
rect 66560 137060 66616 137062
rect 97040 137114 97096 137116
rect 97120 137114 97176 137116
rect 97200 137114 97256 137116
rect 97280 137114 97336 137116
rect 97040 137062 97086 137114
rect 97086 137062 97096 137114
rect 97120 137062 97150 137114
rect 97150 137062 97162 137114
rect 97162 137062 97176 137114
rect 97200 137062 97214 137114
rect 97214 137062 97226 137114
rect 97226 137062 97256 137114
rect 97280 137062 97290 137114
rect 97290 137062 97336 137114
rect 97040 137060 97096 137062
rect 97120 137060 97176 137062
rect 97200 137060 97256 137062
rect 97280 137060 97336 137062
rect 4220 136570 4276 136572
rect 4300 136570 4356 136572
rect 4380 136570 4436 136572
rect 4460 136570 4516 136572
rect 4220 136518 4266 136570
rect 4266 136518 4276 136570
rect 4300 136518 4330 136570
rect 4330 136518 4342 136570
rect 4342 136518 4356 136570
rect 4380 136518 4394 136570
rect 4394 136518 4406 136570
rect 4406 136518 4436 136570
rect 4460 136518 4470 136570
rect 4470 136518 4516 136570
rect 4220 136516 4276 136518
rect 4300 136516 4356 136518
rect 4380 136516 4436 136518
rect 4460 136516 4516 136518
rect 34940 136570 34996 136572
rect 35020 136570 35076 136572
rect 35100 136570 35156 136572
rect 35180 136570 35236 136572
rect 34940 136518 34986 136570
rect 34986 136518 34996 136570
rect 35020 136518 35050 136570
rect 35050 136518 35062 136570
rect 35062 136518 35076 136570
rect 35100 136518 35114 136570
rect 35114 136518 35126 136570
rect 35126 136518 35156 136570
rect 35180 136518 35190 136570
rect 35190 136518 35236 136570
rect 34940 136516 34996 136518
rect 35020 136516 35076 136518
rect 35100 136516 35156 136518
rect 35180 136516 35236 136518
rect 4880 136026 4936 136028
rect 4960 136026 5016 136028
rect 5040 136026 5096 136028
rect 5120 136026 5176 136028
rect 4880 135974 4926 136026
rect 4926 135974 4936 136026
rect 4960 135974 4990 136026
rect 4990 135974 5002 136026
rect 5002 135974 5016 136026
rect 5040 135974 5054 136026
rect 5054 135974 5066 136026
rect 5066 135974 5096 136026
rect 5120 135974 5130 136026
rect 5130 135974 5176 136026
rect 4880 135972 4936 135974
rect 4960 135972 5016 135974
rect 5040 135972 5096 135974
rect 5120 135972 5176 135974
rect 4220 135482 4276 135484
rect 4300 135482 4356 135484
rect 4380 135482 4436 135484
rect 4460 135482 4516 135484
rect 4220 135430 4266 135482
rect 4266 135430 4276 135482
rect 4300 135430 4330 135482
rect 4330 135430 4342 135482
rect 4342 135430 4356 135482
rect 4380 135430 4394 135482
rect 4394 135430 4406 135482
rect 4406 135430 4436 135482
rect 4460 135430 4470 135482
rect 4470 135430 4516 135482
rect 4220 135428 4276 135430
rect 4300 135428 4356 135430
rect 4380 135428 4436 135430
rect 4460 135428 4516 135430
rect 4880 134938 4936 134940
rect 4960 134938 5016 134940
rect 5040 134938 5096 134940
rect 5120 134938 5176 134940
rect 4880 134886 4926 134938
rect 4926 134886 4936 134938
rect 4960 134886 4990 134938
rect 4990 134886 5002 134938
rect 5002 134886 5016 134938
rect 5040 134886 5054 134938
rect 5054 134886 5066 134938
rect 5066 134886 5096 134938
rect 5120 134886 5130 134938
rect 5130 134886 5176 134938
rect 4880 134884 4936 134886
rect 4960 134884 5016 134886
rect 5040 134884 5096 134886
rect 5120 134884 5176 134886
rect 4220 134394 4276 134396
rect 4300 134394 4356 134396
rect 4380 134394 4436 134396
rect 4460 134394 4516 134396
rect 4220 134342 4266 134394
rect 4266 134342 4276 134394
rect 4300 134342 4330 134394
rect 4330 134342 4342 134394
rect 4342 134342 4356 134394
rect 4380 134342 4394 134394
rect 4394 134342 4406 134394
rect 4406 134342 4436 134394
rect 4460 134342 4470 134394
rect 4470 134342 4516 134394
rect 4220 134340 4276 134342
rect 4300 134340 4356 134342
rect 4380 134340 4436 134342
rect 4460 134340 4516 134342
rect 4880 133850 4936 133852
rect 4960 133850 5016 133852
rect 5040 133850 5096 133852
rect 5120 133850 5176 133852
rect 4880 133798 4926 133850
rect 4926 133798 4936 133850
rect 4960 133798 4990 133850
rect 4990 133798 5002 133850
rect 5002 133798 5016 133850
rect 5040 133798 5054 133850
rect 5054 133798 5066 133850
rect 5066 133798 5096 133850
rect 5120 133798 5130 133850
rect 5130 133798 5176 133850
rect 4880 133796 4936 133798
rect 4960 133796 5016 133798
rect 5040 133796 5096 133798
rect 5120 133796 5176 133798
rect 4220 133306 4276 133308
rect 4300 133306 4356 133308
rect 4380 133306 4436 133308
rect 4460 133306 4516 133308
rect 4220 133254 4266 133306
rect 4266 133254 4276 133306
rect 4300 133254 4330 133306
rect 4330 133254 4342 133306
rect 4342 133254 4356 133306
rect 4380 133254 4394 133306
rect 4394 133254 4406 133306
rect 4406 133254 4436 133306
rect 4460 133254 4470 133306
rect 4470 133254 4516 133306
rect 4220 133252 4276 133254
rect 4300 133252 4356 133254
rect 4380 133252 4436 133254
rect 4460 133252 4516 133254
rect 4880 132762 4936 132764
rect 4960 132762 5016 132764
rect 5040 132762 5096 132764
rect 5120 132762 5176 132764
rect 4880 132710 4926 132762
rect 4926 132710 4936 132762
rect 4960 132710 4990 132762
rect 4990 132710 5002 132762
rect 5002 132710 5016 132762
rect 5040 132710 5054 132762
rect 5054 132710 5066 132762
rect 5066 132710 5096 132762
rect 5120 132710 5130 132762
rect 5130 132710 5176 132762
rect 4880 132708 4936 132710
rect 4960 132708 5016 132710
rect 5040 132708 5096 132710
rect 5120 132708 5176 132710
rect 4220 132218 4276 132220
rect 4300 132218 4356 132220
rect 4380 132218 4436 132220
rect 4460 132218 4516 132220
rect 4220 132166 4266 132218
rect 4266 132166 4276 132218
rect 4300 132166 4330 132218
rect 4330 132166 4342 132218
rect 4342 132166 4356 132218
rect 4380 132166 4394 132218
rect 4394 132166 4406 132218
rect 4406 132166 4436 132218
rect 4460 132166 4470 132218
rect 4470 132166 4516 132218
rect 4220 132164 4276 132166
rect 4300 132164 4356 132166
rect 4380 132164 4436 132166
rect 4460 132164 4516 132166
rect 4880 131674 4936 131676
rect 4960 131674 5016 131676
rect 5040 131674 5096 131676
rect 5120 131674 5176 131676
rect 4880 131622 4926 131674
rect 4926 131622 4936 131674
rect 4960 131622 4990 131674
rect 4990 131622 5002 131674
rect 5002 131622 5016 131674
rect 5040 131622 5054 131674
rect 5054 131622 5066 131674
rect 5066 131622 5096 131674
rect 5120 131622 5130 131674
rect 5130 131622 5176 131674
rect 4880 131620 4936 131622
rect 4960 131620 5016 131622
rect 5040 131620 5096 131622
rect 5120 131620 5176 131622
rect 4220 131130 4276 131132
rect 4300 131130 4356 131132
rect 4380 131130 4436 131132
rect 4460 131130 4516 131132
rect 4220 131078 4266 131130
rect 4266 131078 4276 131130
rect 4300 131078 4330 131130
rect 4330 131078 4342 131130
rect 4342 131078 4356 131130
rect 4380 131078 4394 131130
rect 4394 131078 4406 131130
rect 4406 131078 4436 131130
rect 4460 131078 4470 131130
rect 4470 131078 4516 131130
rect 4220 131076 4276 131078
rect 4300 131076 4356 131078
rect 4380 131076 4436 131078
rect 4460 131076 4516 131078
rect 4880 130586 4936 130588
rect 4960 130586 5016 130588
rect 5040 130586 5096 130588
rect 5120 130586 5176 130588
rect 4880 130534 4926 130586
rect 4926 130534 4936 130586
rect 4960 130534 4990 130586
rect 4990 130534 5002 130586
rect 5002 130534 5016 130586
rect 5040 130534 5054 130586
rect 5054 130534 5066 130586
rect 5066 130534 5096 130586
rect 5120 130534 5130 130586
rect 5130 130534 5176 130586
rect 4880 130532 4936 130534
rect 4960 130532 5016 130534
rect 5040 130532 5096 130534
rect 5120 130532 5176 130534
rect 4220 130042 4276 130044
rect 4300 130042 4356 130044
rect 4380 130042 4436 130044
rect 4460 130042 4516 130044
rect 4220 129990 4266 130042
rect 4266 129990 4276 130042
rect 4300 129990 4330 130042
rect 4330 129990 4342 130042
rect 4342 129990 4356 130042
rect 4380 129990 4394 130042
rect 4394 129990 4406 130042
rect 4406 129990 4436 130042
rect 4460 129990 4470 130042
rect 4470 129990 4516 130042
rect 4220 129988 4276 129990
rect 4300 129988 4356 129990
rect 4380 129988 4436 129990
rect 4460 129988 4516 129990
rect 4880 129498 4936 129500
rect 4960 129498 5016 129500
rect 5040 129498 5096 129500
rect 5120 129498 5176 129500
rect 4880 129446 4926 129498
rect 4926 129446 4936 129498
rect 4960 129446 4990 129498
rect 4990 129446 5002 129498
rect 5002 129446 5016 129498
rect 5040 129446 5054 129498
rect 5054 129446 5066 129498
rect 5066 129446 5096 129498
rect 5120 129446 5130 129498
rect 5130 129446 5176 129498
rect 4880 129444 4936 129446
rect 4960 129444 5016 129446
rect 5040 129444 5096 129446
rect 5120 129444 5176 129446
rect 4220 128954 4276 128956
rect 4300 128954 4356 128956
rect 4380 128954 4436 128956
rect 4460 128954 4516 128956
rect 4220 128902 4266 128954
rect 4266 128902 4276 128954
rect 4300 128902 4330 128954
rect 4330 128902 4342 128954
rect 4342 128902 4356 128954
rect 4380 128902 4394 128954
rect 4394 128902 4406 128954
rect 4406 128902 4436 128954
rect 4460 128902 4470 128954
rect 4470 128902 4516 128954
rect 4220 128900 4276 128902
rect 4300 128900 4356 128902
rect 4380 128900 4436 128902
rect 4460 128900 4516 128902
rect 4880 128410 4936 128412
rect 4960 128410 5016 128412
rect 5040 128410 5096 128412
rect 5120 128410 5176 128412
rect 4880 128358 4926 128410
rect 4926 128358 4936 128410
rect 4960 128358 4990 128410
rect 4990 128358 5002 128410
rect 5002 128358 5016 128410
rect 5040 128358 5054 128410
rect 5054 128358 5066 128410
rect 5066 128358 5096 128410
rect 5120 128358 5130 128410
rect 5130 128358 5176 128410
rect 4880 128356 4936 128358
rect 4960 128356 5016 128358
rect 5040 128356 5096 128358
rect 5120 128356 5176 128358
rect 4220 127866 4276 127868
rect 4300 127866 4356 127868
rect 4380 127866 4436 127868
rect 4460 127866 4516 127868
rect 4220 127814 4266 127866
rect 4266 127814 4276 127866
rect 4300 127814 4330 127866
rect 4330 127814 4342 127866
rect 4342 127814 4356 127866
rect 4380 127814 4394 127866
rect 4394 127814 4406 127866
rect 4406 127814 4436 127866
rect 4460 127814 4470 127866
rect 4470 127814 4516 127866
rect 4220 127812 4276 127814
rect 4300 127812 4356 127814
rect 4380 127812 4436 127814
rect 4460 127812 4516 127814
rect 4880 127322 4936 127324
rect 4960 127322 5016 127324
rect 5040 127322 5096 127324
rect 5120 127322 5176 127324
rect 4880 127270 4926 127322
rect 4926 127270 4936 127322
rect 4960 127270 4990 127322
rect 4990 127270 5002 127322
rect 5002 127270 5016 127322
rect 5040 127270 5054 127322
rect 5054 127270 5066 127322
rect 5066 127270 5096 127322
rect 5120 127270 5130 127322
rect 5130 127270 5176 127322
rect 4880 127268 4936 127270
rect 4960 127268 5016 127270
rect 5040 127268 5096 127270
rect 5120 127268 5176 127270
rect 4220 126778 4276 126780
rect 4300 126778 4356 126780
rect 4380 126778 4436 126780
rect 4460 126778 4516 126780
rect 4220 126726 4266 126778
rect 4266 126726 4276 126778
rect 4300 126726 4330 126778
rect 4330 126726 4342 126778
rect 4342 126726 4356 126778
rect 4380 126726 4394 126778
rect 4394 126726 4406 126778
rect 4406 126726 4436 126778
rect 4460 126726 4470 126778
rect 4470 126726 4516 126778
rect 4220 126724 4276 126726
rect 4300 126724 4356 126726
rect 4380 126724 4436 126726
rect 4460 126724 4516 126726
rect 4880 126234 4936 126236
rect 4960 126234 5016 126236
rect 5040 126234 5096 126236
rect 5120 126234 5176 126236
rect 4880 126182 4926 126234
rect 4926 126182 4936 126234
rect 4960 126182 4990 126234
rect 4990 126182 5002 126234
rect 5002 126182 5016 126234
rect 5040 126182 5054 126234
rect 5054 126182 5066 126234
rect 5066 126182 5096 126234
rect 5120 126182 5130 126234
rect 5130 126182 5176 126234
rect 4880 126180 4936 126182
rect 4960 126180 5016 126182
rect 5040 126180 5096 126182
rect 5120 126180 5176 126182
rect 4220 125690 4276 125692
rect 4300 125690 4356 125692
rect 4380 125690 4436 125692
rect 4460 125690 4516 125692
rect 4220 125638 4266 125690
rect 4266 125638 4276 125690
rect 4300 125638 4330 125690
rect 4330 125638 4342 125690
rect 4342 125638 4356 125690
rect 4380 125638 4394 125690
rect 4394 125638 4406 125690
rect 4406 125638 4436 125690
rect 4460 125638 4470 125690
rect 4470 125638 4516 125690
rect 4220 125636 4276 125638
rect 4300 125636 4356 125638
rect 4380 125636 4436 125638
rect 4460 125636 4516 125638
rect 4880 125146 4936 125148
rect 4960 125146 5016 125148
rect 5040 125146 5096 125148
rect 5120 125146 5176 125148
rect 4880 125094 4926 125146
rect 4926 125094 4936 125146
rect 4960 125094 4990 125146
rect 4990 125094 5002 125146
rect 5002 125094 5016 125146
rect 5040 125094 5054 125146
rect 5054 125094 5066 125146
rect 5066 125094 5096 125146
rect 5120 125094 5130 125146
rect 5130 125094 5176 125146
rect 4880 125092 4936 125094
rect 4960 125092 5016 125094
rect 5040 125092 5096 125094
rect 5120 125092 5176 125094
rect 4220 124602 4276 124604
rect 4300 124602 4356 124604
rect 4380 124602 4436 124604
rect 4460 124602 4516 124604
rect 4220 124550 4266 124602
rect 4266 124550 4276 124602
rect 4300 124550 4330 124602
rect 4330 124550 4342 124602
rect 4342 124550 4356 124602
rect 4380 124550 4394 124602
rect 4394 124550 4406 124602
rect 4406 124550 4436 124602
rect 4460 124550 4470 124602
rect 4470 124550 4516 124602
rect 4220 124548 4276 124550
rect 4300 124548 4356 124550
rect 4380 124548 4436 124550
rect 4460 124548 4516 124550
rect 4880 124058 4936 124060
rect 4960 124058 5016 124060
rect 5040 124058 5096 124060
rect 5120 124058 5176 124060
rect 4880 124006 4926 124058
rect 4926 124006 4936 124058
rect 4960 124006 4990 124058
rect 4990 124006 5002 124058
rect 5002 124006 5016 124058
rect 5040 124006 5054 124058
rect 5054 124006 5066 124058
rect 5066 124006 5096 124058
rect 5120 124006 5130 124058
rect 5130 124006 5176 124058
rect 4880 124004 4936 124006
rect 4960 124004 5016 124006
rect 5040 124004 5096 124006
rect 5120 124004 5176 124006
rect 4220 123514 4276 123516
rect 4300 123514 4356 123516
rect 4380 123514 4436 123516
rect 4460 123514 4516 123516
rect 4220 123462 4266 123514
rect 4266 123462 4276 123514
rect 4300 123462 4330 123514
rect 4330 123462 4342 123514
rect 4342 123462 4356 123514
rect 4380 123462 4394 123514
rect 4394 123462 4406 123514
rect 4406 123462 4436 123514
rect 4460 123462 4470 123514
rect 4470 123462 4516 123514
rect 4220 123460 4276 123462
rect 4300 123460 4356 123462
rect 4380 123460 4436 123462
rect 4460 123460 4516 123462
rect 4880 122970 4936 122972
rect 4960 122970 5016 122972
rect 5040 122970 5096 122972
rect 5120 122970 5176 122972
rect 4880 122918 4926 122970
rect 4926 122918 4936 122970
rect 4960 122918 4990 122970
rect 4990 122918 5002 122970
rect 5002 122918 5016 122970
rect 5040 122918 5054 122970
rect 5054 122918 5066 122970
rect 5066 122918 5096 122970
rect 5120 122918 5130 122970
rect 5130 122918 5176 122970
rect 4880 122916 4936 122918
rect 4960 122916 5016 122918
rect 5040 122916 5096 122918
rect 5120 122916 5176 122918
rect 4220 122426 4276 122428
rect 4300 122426 4356 122428
rect 4380 122426 4436 122428
rect 4460 122426 4516 122428
rect 4220 122374 4266 122426
rect 4266 122374 4276 122426
rect 4300 122374 4330 122426
rect 4330 122374 4342 122426
rect 4342 122374 4356 122426
rect 4380 122374 4394 122426
rect 4394 122374 4406 122426
rect 4406 122374 4436 122426
rect 4460 122374 4470 122426
rect 4470 122374 4516 122426
rect 4220 122372 4276 122374
rect 4300 122372 4356 122374
rect 4380 122372 4436 122374
rect 4460 122372 4516 122374
rect 4880 121882 4936 121884
rect 4960 121882 5016 121884
rect 5040 121882 5096 121884
rect 5120 121882 5176 121884
rect 4880 121830 4926 121882
rect 4926 121830 4936 121882
rect 4960 121830 4990 121882
rect 4990 121830 5002 121882
rect 5002 121830 5016 121882
rect 5040 121830 5054 121882
rect 5054 121830 5066 121882
rect 5066 121830 5096 121882
rect 5120 121830 5130 121882
rect 5130 121830 5176 121882
rect 4880 121828 4936 121830
rect 4960 121828 5016 121830
rect 5040 121828 5096 121830
rect 5120 121828 5176 121830
rect 4220 121338 4276 121340
rect 4300 121338 4356 121340
rect 4380 121338 4436 121340
rect 4460 121338 4516 121340
rect 4220 121286 4266 121338
rect 4266 121286 4276 121338
rect 4300 121286 4330 121338
rect 4330 121286 4342 121338
rect 4342 121286 4356 121338
rect 4380 121286 4394 121338
rect 4394 121286 4406 121338
rect 4406 121286 4436 121338
rect 4460 121286 4470 121338
rect 4470 121286 4516 121338
rect 4220 121284 4276 121286
rect 4300 121284 4356 121286
rect 4380 121284 4436 121286
rect 4460 121284 4516 121286
rect 4880 120794 4936 120796
rect 4960 120794 5016 120796
rect 5040 120794 5096 120796
rect 5120 120794 5176 120796
rect 4880 120742 4926 120794
rect 4926 120742 4936 120794
rect 4960 120742 4990 120794
rect 4990 120742 5002 120794
rect 5002 120742 5016 120794
rect 5040 120742 5054 120794
rect 5054 120742 5066 120794
rect 5066 120742 5096 120794
rect 5120 120742 5130 120794
rect 5130 120742 5176 120794
rect 4880 120740 4936 120742
rect 4960 120740 5016 120742
rect 5040 120740 5096 120742
rect 5120 120740 5176 120742
rect 4220 120250 4276 120252
rect 4300 120250 4356 120252
rect 4380 120250 4436 120252
rect 4460 120250 4516 120252
rect 4220 120198 4266 120250
rect 4266 120198 4276 120250
rect 4300 120198 4330 120250
rect 4330 120198 4342 120250
rect 4342 120198 4356 120250
rect 4380 120198 4394 120250
rect 4394 120198 4406 120250
rect 4406 120198 4436 120250
rect 4460 120198 4470 120250
rect 4470 120198 4516 120250
rect 4220 120196 4276 120198
rect 4300 120196 4356 120198
rect 4380 120196 4436 120198
rect 4460 120196 4516 120198
rect 4880 119706 4936 119708
rect 4960 119706 5016 119708
rect 5040 119706 5096 119708
rect 5120 119706 5176 119708
rect 4880 119654 4926 119706
rect 4926 119654 4936 119706
rect 4960 119654 4990 119706
rect 4990 119654 5002 119706
rect 5002 119654 5016 119706
rect 5040 119654 5054 119706
rect 5054 119654 5066 119706
rect 5066 119654 5096 119706
rect 5120 119654 5130 119706
rect 5130 119654 5176 119706
rect 4880 119652 4936 119654
rect 4960 119652 5016 119654
rect 5040 119652 5096 119654
rect 5120 119652 5176 119654
rect 4220 119162 4276 119164
rect 4300 119162 4356 119164
rect 4380 119162 4436 119164
rect 4460 119162 4516 119164
rect 4220 119110 4266 119162
rect 4266 119110 4276 119162
rect 4300 119110 4330 119162
rect 4330 119110 4342 119162
rect 4342 119110 4356 119162
rect 4380 119110 4394 119162
rect 4394 119110 4406 119162
rect 4406 119110 4436 119162
rect 4460 119110 4470 119162
rect 4470 119110 4516 119162
rect 4220 119108 4276 119110
rect 4300 119108 4356 119110
rect 4380 119108 4436 119110
rect 4460 119108 4516 119110
rect 4880 118618 4936 118620
rect 4960 118618 5016 118620
rect 5040 118618 5096 118620
rect 5120 118618 5176 118620
rect 4880 118566 4926 118618
rect 4926 118566 4936 118618
rect 4960 118566 4990 118618
rect 4990 118566 5002 118618
rect 5002 118566 5016 118618
rect 5040 118566 5054 118618
rect 5054 118566 5066 118618
rect 5066 118566 5096 118618
rect 5120 118566 5130 118618
rect 5130 118566 5176 118618
rect 4880 118564 4936 118566
rect 4960 118564 5016 118566
rect 5040 118564 5096 118566
rect 5120 118564 5176 118566
rect 4220 118074 4276 118076
rect 4300 118074 4356 118076
rect 4380 118074 4436 118076
rect 4460 118074 4516 118076
rect 4220 118022 4266 118074
rect 4266 118022 4276 118074
rect 4300 118022 4330 118074
rect 4330 118022 4342 118074
rect 4342 118022 4356 118074
rect 4380 118022 4394 118074
rect 4394 118022 4406 118074
rect 4406 118022 4436 118074
rect 4460 118022 4470 118074
rect 4470 118022 4516 118074
rect 4220 118020 4276 118022
rect 4300 118020 4356 118022
rect 4380 118020 4436 118022
rect 4460 118020 4516 118022
rect 4880 117530 4936 117532
rect 4960 117530 5016 117532
rect 5040 117530 5096 117532
rect 5120 117530 5176 117532
rect 4880 117478 4926 117530
rect 4926 117478 4936 117530
rect 4960 117478 4990 117530
rect 4990 117478 5002 117530
rect 5002 117478 5016 117530
rect 5040 117478 5054 117530
rect 5054 117478 5066 117530
rect 5066 117478 5096 117530
rect 5120 117478 5130 117530
rect 5130 117478 5176 117530
rect 4880 117476 4936 117478
rect 4960 117476 5016 117478
rect 5040 117476 5096 117478
rect 5120 117476 5176 117478
rect 4220 116986 4276 116988
rect 4300 116986 4356 116988
rect 4380 116986 4436 116988
rect 4460 116986 4516 116988
rect 4220 116934 4266 116986
rect 4266 116934 4276 116986
rect 4300 116934 4330 116986
rect 4330 116934 4342 116986
rect 4342 116934 4356 116986
rect 4380 116934 4394 116986
rect 4394 116934 4406 116986
rect 4406 116934 4436 116986
rect 4460 116934 4470 116986
rect 4470 116934 4516 116986
rect 4220 116932 4276 116934
rect 4300 116932 4356 116934
rect 4380 116932 4436 116934
rect 4460 116932 4516 116934
rect 4880 116442 4936 116444
rect 4960 116442 5016 116444
rect 5040 116442 5096 116444
rect 5120 116442 5176 116444
rect 4880 116390 4926 116442
rect 4926 116390 4936 116442
rect 4960 116390 4990 116442
rect 4990 116390 5002 116442
rect 5002 116390 5016 116442
rect 5040 116390 5054 116442
rect 5054 116390 5066 116442
rect 5066 116390 5096 116442
rect 5120 116390 5130 116442
rect 5130 116390 5176 116442
rect 4880 116388 4936 116390
rect 4960 116388 5016 116390
rect 5040 116388 5096 116390
rect 5120 116388 5176 116390
rect 4220 115898 4276 115900
rect 4300 115898 4356 115900
rect 4380 115898 4436 115900
rect 4460 115898 4516 115900
rect 4220 115846 4266 115898
rect 4266 115846 4276 115898
rect 4300 115846 4330 115898
rect 4330 115846 4342 115898
rect 4342 115846 4356 115898
rect 4380 115846 4394 115898
rect 4394 115846 4406 115898
rect 4406 115846 4436 115898
rect 4460 115846 4470 115898
rect 4470 115846 4516 115898
rect 4220 115844 4276 115846
rect 4300 115844 4356 115846
rect 4380 115844 4436 115846
rect 4460 115844 4516 115846
rect 4880 115354 4936 115356
rect 4960 115354 5016 115356
rect 5040 115354 5096 115356
rect 5120 115354 5176 115356
rect 4880 115302 4926 115354
rect 4926 115302 4936 115354
rect 4960 115302 4990 115354
rect 4990 115302 5002 115354
rect 5002 115302 5016 115354
rect 5040 115302 5054 115354
rect 5054 115302 5066 115354
rect 5066 115302 5096 115354
rect 5120 115302 5130 115354
rect 5130 115302 5176 115354
rect 4880 115300 4936 115302
rect 4960 115300 5016 115302
rect 5040 115300 5096 115302
rect 5120 115300 5176 115302
rect 4220 114810 4276 114812
rect 4300 114810 4356 114812
rect 4380 114810 4436 114812
rect 4460 114810 4516 114812
rect 4220 114758 4266 114810
rect 4266 114758 4276 114810
rect 4300 114758 4330 114810
rect 4330 114758 4342 114810
rect 4342 114758 4356 114810
rect 4380 114758 4394 114810
rect 4394 114758 4406 114810
rect 4406 114758 4436 114810
rect 4460 114758 4470 114810
rect 4470 114758 4516 114810
rect 4220 114756 4276 114758
rect 4300 114756 4356 114758
rect 4380 114756 4436 114758
rect 4460 114756 4516 114758
rect 4880 114266 4936 114268
rect 4960 114266 5016 114268
rect 5040 114266 5096 114268
rect 5120 114266 5176 114268
rect 4880 114214 4926 114266
rect 4926 114214 4936 114266
rect 4960 114214 4990 114266
rect 4990 114214 5002 114266
rect 5002 114214 5016 114266
rect 5040 114214 5054 114266
rect 5054 114214 5066 114266
rect 5066 114214 5096 114266
rect 5120 114214 5130 114266
rect 5130 114214 5176 114266
rect 4880 114212 4936 114214
rect 4960 114212 5016 114214
rect 5040 114212 5096 114214
rect 5120 114212 5176 114214
rect 4220 113722 4276 113724
rect 4300 113722 4356 113724
rect 4380 113722 4436 113724
rect 4460 113722 4516 113724
rect 4220 113670 4266 113722
rect 4266 113670 4276 113722
rect 4300 113670 4330 113722
rect 4330 113670 4342 113722
rect 4342 113670 4356 113722
rect 4380 113670 4394 113722
rect 4394 113670 4406 113722
rect 4406 113670 4436 113722
rect 4460 113670 4470 113722
rect 4470 113670 4516 113722
rect 4220 113668 4276 113670
rect 4300 113668 4356 113670
rect 4380 113668 4436 113670
rect 4460 113668 4516 113670
rect 4880 113178 4936 113180
rect 4960 113178 5016 113180
rect 5040 113178 5096 113180
rect 5120 113178 5176 113180
rect 4880 113126 4926 113178
rect 4926 113126 4936 113178
rect 4960 113126 4990 113178
rect 4990 113126 5002 113178
rect 5002 113126 5016 113178
rect 5040 113126 5054 113178
rect 5054 113126 5066 113178
rect 5066 113126 5096 113178
rect 5120 113126 5130 113178
rect 5130 113126 5176 113178
rect 4880 113124 4936 113126
rect 4960 113124 5016 113126
rect 5040 113124 5096 113126
rect 5120 113124 5176 113126
rect 4220 112634 4276 112636
rect 4300 112634 4356 112636
rect 4380 112634 4436 112636
rect 4460 112634 4516 112636
rect 4220 112582 4266 112634
rect 4266 112582 4276 112634
rect 4300 112582 4330 112634
rect 4330 112582 4342 112634
rect 4342 112582 4356 112634
rect 4380 112582 4394 112634
rect 4394 112582 4406 112634
rect 4406 112582 4436 112634
rect 4460 112582 4470 112634
rect 4470 112582 4516 112634
rect 4220 112580 4276 112582
rect 4300 112580 4356 112582
rect 4380 112580 4436 112582
rect 4460 112580 4516 112582
rect 4880 112090 4936 112092
rect 4960 112090 5016 112092
rect 5040 112090 5096 112092
rect 5120 112090 5176 112092
rect 4880 112038 4926 112090
rect 4926 112038 4936 112090
rect 4960 112038 4990 112090
rect 4990 112038 5002 112090
rect 5002 112038 5016 112090
rect 5040 112038 5054 112090
rect 5054 112038 5066 112090
rect 5066 112038 5096 112090
rect 5120 112038 5130 112090
rect 5130 112038 5176 112090
rect 4880 112036 4936 112038
rect 4960 112036 5016 112038
rect 5040 112036 5096 112038
rect 5120 112036 5176 112038
rect 4220 111546 4276 111548
rect 4300 111546 4356 111548
rect 4380 111546 4436 111548
rect 4460 111546 4516 111548
rect 4220 111494 4266 111546
rect 4266 111494 4276 111546
rect 4300 111494 4330 111546
rect 4330 111494 4342 111546
rect 4342 111494 4356 111546
rect 4380 111494 4394 111546
rect 4394 111494 4406 111546
rect 4406 111494 4436 111546
rect 4460 111494 4470 111546
rect 4470 111494 4516 111546
rect 4220 111492 4276 111494
rect 4300 111492 4356 111494
rect 4380 111492 4436 111494
rect 4460 111492 4516 111494
rect 4880 111002 4936 111004
rect 4960 111002 5016 111004
rect 5040 111002 5096 111004
rect 5120 111002 5176 111004
rect 4880 110950 4926 111002
rect 4926 110950 4936 111002
rect 4960 110950 4990 111002
rect 4990 110950 5002 111002
rect 5002 110950 5016 111002
rect 5040 110950 5054 111002
rect 5054 110950 5066 111002
rect 5066 110950 5096 111002
rect 5120 110950 5130 111002
rect 5130 110950 5176 111002
rect 4880 110948 4936 110950
rect 4960 110948 5016 110950
rect 5040 110948 5096 110950
rect 5120 110948 5176 110950
rect 1306 110880 1362 110936
rect 4220 110458 4276 110460
rect 4300 110458 4356 110460
rect 4380 110458 4436 110460
rect 4460 110458 4516 110460
rect 4220 110406 4266 110458
rect 4266 110406 4276 110458
rect 4300 110406 4330 110458
rect 4330 110406 4342 110458
rect 4342 110406 4356 110458
rect 4380 110406 4394 110458
rect 4394 110406 4406 110458
rect 4406 110406 4436 110458
rect 4460 110406 4470 110458
rect 4470 110406 4516 110458
rect 4220 110404 4276 110406
rect 4300 110404 4356 110406
rect 4380 110404 4436 110406
rect 4460 110404 4516 110406
rect 4880 109914 4936 109916
rect 4960 109914 5016 109916
rect 5040 109914 5096 109916
rect 5120 109914 5176 109916
rect 4880 109862 4926 109914
rect 4926 109862 4936 109914
rect 4960 109862 4990 109914
rect 4990 109862 5002 109914
rect 5002 109862 5016 109914
rect 5040 109862 5054 109914
rect 5054 109862 5066 109914
rect 5066 109862 5096 109914
rect 5120 109862 5130 109914
rect 5130 109862 5176 109914
rect 4880 109860 4936 109862
rect 4960 109860 5016 109862
rect 5040 109860 5096 109862
rect 5120 109860 5176 109862
rect 1306 109520 1362 109576
rect 4220 109370 4276 109372
rect 4300 109370 4356 109372
rect 4380 109370 4436 109372
rect 4460 109370 4516 109372
rect 4220 109318 4266 109370
rect 4266 109318 4276 109370
rect 4300 109318 4330 109370
rect 4330 109318 4342 109370
rect 4342 109318 4356 109370
rect 4380 109318 4394 109370
rect 4394 109318 4406 109370
rect 4406 109318 4436 109370
rect 4460 109318 4470 109370
rect 4470 109318 4516 109370
rect 4220 109316 4276 109318
rect 4300 109316 4356 109318
rect 4380 109316 4436 109318
rect 4460 109316 4516 109318
rect 4880 108826 4936 108828
rect 4960 108826 5016 108828
rect 5040 108826 5096 108828
rect 5120 108826 5176 108828
rect 4880 108774 4926 108826
rect 4926 108774 4936 108826
rect 4960 108774 4990 108826
rect 4990 108774 5002 108826
rect 5002 108774 5016 108826
rect 5040 108774 5054 108826
rect 5054 108774 5066 108826
rect 5066 108774 5096 108826
rect 5120 108774 5130 108826
rect 5130 108774 5176 108826
rect 4880 108772 4936 108774
rect 4960 108772 5016 108774
rect 5040 108772 5096 108774
rect 5120 108772 5176 108774
rect 4220 108282 4276 108284
rect 4300 108282 4356 108284
rect 4380 108282 4436 108284
rect 4460 108282 4516 108284
rect 4220 108230 4266 108282
rect 4266 108230 4276 108282
rect 4300 108230 4330 108282
rect 4330 108230 4342 108282
rect 4342 108230 4356 108282
rect 4380 108230 4394 108282
rect 4394 108230 4406 108282
rect 4406 108230 4436 108282
rect 4460 108230 4470 108282
rect 4470 108230 4516 108282
rect 4220 108228 4276 108230
rect 4300 108228 4356 108230
rect 4380 108228 4436 108230
rect 4460 108228 4516 108230
rect 1306 108160 1362 108216
rect 4880 107738 4936 107740
rect 4960 107738 5016 107740
rect 5040 107738 5096 107740
rect 5120 107738 5176 107740
rect 4880 107686 4926 107738
rect 4926 107686 4936 107738
rect 4960 107686 4990 107738
rect 4990 107686 5002 107738
rect 5002 107686 5016 107738
rect 5040 107686 5054 107738
rect 5054 107686 5066 107738
rect 5066 107686 5096 107738
rect 5120 107686 5130 107738
rect 5130 107686 5176 107738
rect 4880 107684 4936 107686
rect 4960 107684 5016 107686
rect 5040 107684 5096 107686
rect 5120 107684 5176 107686
rect 4220 107194 4276 107196
rect 4300 107194 4356 107196
rect 4380 107194 4436 107196
rect 4460 107194 4516 107196
rect 4220 107142 4266 107194
rect 4266 107142 4276 107194
rect 4300 107142 4330 107194
rect 4330 107142 4342 107194
rect 4342 107142 4356 107194
rect 4380 107142 4394 107194
rect 4394 107142 4406 107194
rect 4406 107142 4436 107194
rect 4460 107142 4470 107194
rect 4470 107142 4516 107194
rect 4220 107140 4276 107142
rect 4300 107140 4356 107142
rect 4380 107140 4436 107142
rect 4460 107140 4516 107142
rect 1214 106836 1216 106856
rect 1216 106836 1268 106856
rect 1268 106836 1270 106856
rect 1214 106800 1270 106836
rect 4880 106650 4936 106652
rect 4960 106650 5016 106652
rect 5040 106650 5096 106652
rect 5120 106650 5176 106652
rect 4880 106598 4926 106650
rect 4926 106598 4936 106650
rect 4960 106598 4990 106650
rect 4990 106598 5002 106650
rect 5002 106598 5016 106650
rect 5040 106598 5054 106650
rect 5054 106598 5066 106650
rect 5066 106598 5096 106650
rect 5120 106598 5130 106650
rect 5130 106598 5176 106650
rect 4880 106596 4936 106598
rect 4960 106596 5016 106598
rect 5040 106596 5096 106598
rect 5120 106596 5176 106598
rect 4220 106106 4276 106108
rect 4300 106106 4356 106108
rect 4380 106106 4436 106108
rect 4460 106106 4516 106108
rect 4220 106054 4266 106106
rect 4266 106054 4276 106106
rect 4300 106054 4330 106106
rect 4330 106054 4342 106106
rect 4342 106054 4356 106106
rect 4380 106054 4394 106106
rect 4394 106054 4406 106106
rect 4406 106054 4436 106106
rect 4460 106054 4470 106106
rect 4470 106054 4516 106106
rect 4220 106052 4276 106054
rect 4300 106052 4356 106054
rect 4380 106052 4436 106054
rect 4460 106052 4516 106054
rect 4880 105562 4936 105564
rect 4960 105562 5016 105564
rect 5040 105562 5096 105564
rect 5120 105562 5176 105564
rect 4880 105510 4926 105562
rect 4926 105510 4936 105562
rect 4960 105510 4990 105562
rect 4990 105510 5002 105562
rect 5002 105510 5016 105562
rect 5040 105510 5054 105562
rect 5054 105510 5066 105562
rect 5066 105510 5096 105562
rect 5120 105510 5130 105562
rect 5130 105510 5176 105562
rect 4880 105508 4936 105510
rect 4960 105508 5016 105510
rect 5040 105508 5096 105510
rect 5120 105508 5176 105510
rect 1306 105440 1362 105496
rect 4220 105018 4276 105020
rect 4300 105018 4356 105020
rect 4380 105018 4436 105020
rect 4460 105018 4516 105020
rect 4220 104966 4266 105018
rect 4266 104966 4276 105018
rect 4300 104966 4330 105018
rect 4330 104966 4342 105018
rect 4342 104966 4356 105018
rect 4380 104966 4394 105018
rect 4394 104966 4406 105018
rect 4406 104966 4436 105018
rect 4460 104966 4470 105018
rect 4470 104966 4516 105018
rect 4220 104964 4276 104966
rect 4300 104964 4356 104966
rect 4380 104964 4436 104966
rect 4460 104964 4516 104966
rect 4880 104474 4936 104476
rect 4960 104474 5016 104476
rect 5040 104474 5096 104476
rect 5120 104474 5176 104476
rect 4880 104422 4926 104474
rect 4926 104422 4936 104474
rect 4960 104422 4990 104474
rect 4990 104422 5002 104474
rect 5002 104422 5016 104474
rect 5040 104422 5054 104474
rect 5054 104422 5066 104474
rect 5066 104422 5096 104474
rect 5120 104422 5130 104474
rect 5130 104422 5176 104474
rect 4880 104420 4936 104422
rect 4960 104420 5016 104422
rect 5040 104420 5096 104422
rect 5120 104420 5176 104422
rect 1306 104080 1362 104136
rect 4220 103930 4276 103932
rect 4300 103930 4356 103932
rect 4380 103930 4436 103932
rect 4460 103930 4516 103932
rect 4220 103878 4266 103930
rect 4266 103878 4276 103930
rect 4300 103878 4330 103930
rect 4330 103878 4342 103930
rect 4342 103878 4356 103930
rect 4380 103878 4394 103930
rect 4394 103878 4406 103930
rect 4406 103878 4436 103930
rect 4460 103878 4470 103930
rect 4470 103878 4516 103930
rect 4220 103876 4276 103878
rect 4300 103876 4356 103878
rect 4380 103876 4436 103878
rect 4460 103876 4516 103878
rect 4880 103386 4936 103388
rect 4960 103386 5016 103388
rect 5040 103386 5096 103388
rect 5120 103386 5176 103388
rect 4880 103334 4926 103386
rect 4926 103334 4936 103386
rect 4960 103334 4990 103386
rect 4990 103334 5002 103386
rect 5002 103334 5016 103386
rect 5040 103334 5054 103386
rect 5054 103334 5066 103386
rect 5066 103334 5096 103386
rect 5120 103334 5130 103386
rect 5130 103334 5176 103386
rect 4880 103332 4936 103334
rect 4960 103332 5016 103334
rect 5040 103332 5096 103334
rect 5120 103332 5176 103334
rect 4220 102842 4276 102844
rect 4300 102842 4356 102844
rect 4380 102842 4436 102844
rect 4460 102842 4516 102844
rect 4220 102790 4266 102842
rect 4266 102790 4276 102842
rect 4300 102790 4330 102842
rect 4330 102790 4342 102842
rect 4342 102790 4356 102842
rect 4380 102790 4394 102842
rect 4394 102790 4406 102842
rect 4406 102790 4436 102842
rect 4460 102790 4470 102842
rect 4470 102790 4516 102842
rect 4220 102788 4276 102790
rect 4300 102788 4356 102790
rect 4380 102788 4436 102790
rect 4460 102788 4516 102790
rect 4880 102298 4936 102300
rect 4960 102298 5016 102300
rect 5040 102298 5096 102300
rect 5120 102298 5176 102300
rect 4880 102246 4926 102298
rect 4926 102246 4936 102298
rect 4960 102246 4990 102298
rect 4990 102246 5002 102298
rect 5002 102246 5016 102298
rect 5040 102246 5054 102298
rect 5054 102246 5066 102298
rect 5066 102246 5096 102298
rect 5120 102246 5130 102298
rect 5130 102246 5176 102298
rect 4880 102244 4936 102246
rect 4960 102244 5016 102246
rect 5040 102244 5096 102246
rect 5120 102244 5176 102246
rect 4220 101754 4276 101756
rect 4300 101754 4356 101756
rect 4380 101754 4436 101756
rect 4460 101754 4516 101756
rect 4220 101702 4266 101754
rect 4266 101702 4276 101754
rect 4300 101702 4330 101754
rect 4330 101702 4342 101754
rect 4342 101702 4356 101754
rect 4380 101702 4394 101754
rect 4394 101702 4406 101754
rect 4406 101702 4436 101754
rect 4460 101702 4470 101754
rect 4470 101702 4516 101754
rect 4220 101700 4276 101702
rect 4300 101700 4356 101702
rect 4380 101700 4436 101702
rect 4460 101700 4516 101702
rect 4880 101210 4936 101212
rect 4960 101210 5016 101212
rect 5040 101210 5096 101212
rect 5120 101210 5176 101212
rect 4880 101158 4926 101210
rect 4926 101158 4936 101210
rect 4960 101158 4990 101210
rect 4990 101158 5002 101210
rect 5002 101158 5016 101210
rect 5040 101158 5054 101210
rect 5054 101158 5066 101210
rect 5066 101158 5096 101210
rect 5120 101158 5130 101210
rect 5130 101158 5176 101210
rect 4880 101156 4936 101158
rect 4960 101156 5016 101158
rect 5040 101156 5096 101158
rect 5120 101156 5176 101158
rect 4220 100666 4276 100668
rect 4300 100666 4356 100668
rect 4380 100666 4436 100668
rect 4460 100666 4516 100668
rect 4220 100614 4266 100666
rect 4266 100614 4276 100666
rect 4300 100614 4330 100666
rect 4330 100614 4342 100666
rect 4342 100614 4356 100666
rect 4380 100614 4394 100666
rect 4394 100614 4406 100666
rect 4406 100614 4436 100666
rect 4460 100614 4470 100666
rect 4470 100614 4516 100666
rect 4220 100612 4276 100614
rect 4300 100612 4356 100614
rect 4380 100612 4436 100614
rect 4460 100612 4516 100614
rect 4880 100122 4936 100124
rect 4960 100122 5016 100124
rect 5040 100122 5096 100124
rect 5120 100122 5176 100124
rect 4880 100070 4926 100122
rect 4926 100070 4936 100122
rect 4960 100070 4990 100122
rect 4990 100070 5002 100122
rect 5002 100070 5016 100122
rect 5040 100070 5054 100122
rect 5054 100070 5066 100122
rect 5066 100070 5096 100122
rect 5120 100070 5130 100122
rect 5130 100070 5176 100122
rect 4880 100068 4936 100070
rect 4960 100068 5016 100070
rect 5040 100068 5096 100070
rect 5120 100068 5176 100070
rect 4220 99578 4276 99580
rect 4300 99578 4356 99580
rect 4380 99578 4436 99580
rect 4460 99578 4516 99580
rect 4220 99526 4266 99578
rect 4266 99526 4276 99578
rect 4300 99526 4330 99578
rect 4330 99526 4342 99578
rect 4342 99526 4356 99578
rect 4380 99526 4394 99578
rect 4394 99526 4406 99578
rect 4406 99526 4436 99578
rect 4460 99526 4470 99578
rect 4470 99526 4516 99578
rect 4220 99524 4276 99526
rect 4300 99524 4356 99526
rect 4380 99524 4436 99526
rect 4460 99524 4516 99526
rect 4880 99034 4936 99036
rect 4960 99034 5016 99036
rect 5040 99034 5096 99036
rect 5120 99034 5176 99036
rect 4880 98982 4926 99034
rect 4926 98982 4936 99034
rect 4960 98982 4990 99034
rect 4990 98982 5002 99034
rect 5002 98982 5016 99034
rect 5040 98982 5054 99034
rect 5054 98982 5066 99034
rect 5066 98982 5096 99034
rect 5120 98982 5130 99034
rect 5130 98982 5176 99034
rect 4880 98980 4936 98982
rect 4960 98980 5016 98982
rect 5040 98980 5096 98982
rect 5120 98980 5176 98982
rect 4220 98490 4276 98492
rect 4300 98490 4356 98492
rect 4380 98490 4436 98492
rect 4460 98490 4516 98492
rect 4220 98438 4266 98490
rect 4266 98438 4276 98490
rect 4300 98438 4330 98490
rect 4330 98438 4342 98490
rect 4342 98438 4356 98490
rect 4380 98438 4394 98490
rect 4394 98438 4406 98490
rect 4406 98438 4436 98490
rect 4460 98438 4470 98490
rect 4470 98438 4516 98490
rect 4220 98436 4276 98438
rect 4300 98436 4356 98438
rect 4380 98436 4436 98438
rect 4460 98436 4516 98438
rect 4880 97946 4936 97948
rect 4960 97946 5016 97948
rect 5040 97946 5096 97948
rect 5120 97946 5176 97948
rect 4880 97894 4926 97946
rect 4926 97894 4936 97946
rect 4960 97894 4990 97946
rect 4990 97894 5002 97946
rect 5002 97894 5016 97946
rect 5040 97894 5054 97946
rect 5054 97894 5066 97946
rect 5066 97894 5096 97946
rect 5120 97894 5130 97946
rect 5130 97894 5176 97946
rect 4880 97892 4936 97894
rect 4960 97892 5016 97894
rect 5040 97892 5096 97894
rect 5120 97892 5176 97894
rect 4220 97402 4276 97404
rect 4300 97402 4356 97404
rect 4380 97402 4436 97404
rect 4460 97402 4516 97404
rect 4220 97350 4266 97402
rect 4266 97350 4276 97402
rect 4300 97350 4330 97402
rect 4330 97350 4342 97402
rect 4342 97350 4356 97402
rect 4380 97350 4394 97402
rect 4394 97350 4406 97402
rect 4406 97350 4436 97402
rect 4460 97350 4470 97402
rect 4470 97350 4516 97402
rect 4220 97348 4276 97350
rect 4300 97348 4356 97350
rect 4380 97348 4436 97350
rect 4460 97348 4516 97350
rect 4880 96858 4936 96860
rect 4960 96858 5016 96860
rect 5040 96858 5096 96860
rect 5120 96858 5176 96860
rect 4880 96806 4926 96858
rect 4926 96806 4936 96858
rect 4960 96806 4990 96858
rect 4990 96806 5002 96858
rect 5002 96806 5016 96858
rect 5040 96806 5054 96858
rect 5054 96806 5066 96858
rect 5066 96806 5096 96858
rect 5120 96806 5130 96858
rect 5130 96806 5176 96858
rect 4880 96804 4936 96806
rect 4960 96804 5016 96806
rect 5040 96804 5096 96806
rect 5120 96804 5176 96806
rect 4220 96314 4276 96316
rect 4300 96314 4356 96316
rect 4380 96314 4436 96316
rect 4460 96314 4516 96316
rect 4220 96262 4266 96314
rect 4266 96262 4276 96314
rect 4300 96262 4330 96314
rect 4330 96262 4342 96314
rect 4342 96262 4356 96314
rect 4380 96262 4394 96314
rect 4394 96262 4406 96314
rect 4406 96262 4436 96314
rect 4460 96262 4470 96314
rect 4470 96262 4516 96314
rect 4220 96260 4276 96262
rect 4300 96260 4356 96262
rect 4380 96260 4436 96262
rect 4460 96260 4516 96262
rect 4880 95770 4936 95772
rect 4960 95770 5016 95772
rect 5040 95770 5096 95772
rect 5120 95770 5176 95772
rect 4880 95718 4926 95770
rect 4926 95718 4936 95770
rect 4960 95718 4990 95770
rect 4990 95718 5002 95770
rect 5002 95718 5016 95770
rect 5040 95718 5054 95770
rect 5054 95718 5066 95770
rect 5066 95718 5096 95770
rect 5120 95718 5130 95770
rect 5130 95718 5176 95770
rect 4880 95716 4936 95718
rect 4960 95716 5016 95718
rect 5040 95716 5096 95718
rect 5120 95716 5176 95718
rect 4220 95226 4276 95228
rect 4300 95226 4356 95228
rect 4380 95226 4436 95228
rect 4460 95226 4516 95228
rect 4220 95174 4266 95226
rect 4266 95174 4276 95226
rect 4300 95174 4330 95226
rect 4330 95174 4342 95226
rect 4342 95174 4356 95226
rect 4380 95174 4394 95226
rect 4394 95174 4406 95226
rect 4406 95174 4436 95226
rect 4460 95174 4470 95226
rect 4470 95174 4516 95226
rect 4220 95172 4276 95174
rect 4300 95172 4356 95174
rect 4380 95172 4436 95174
rect 4460 95172 4516 95174
rect 4880 94682 4936 94684
rect 4960 94682 5016 94684
rect 5040 94682 5096 94684
rect 5120 94682 5176 94684
rect 4880 94630 4926 94682
rect 4926 94630 4936 94682
rect 4960 94630 4990 94682
rect 4990 94630 5002 94682
rect 5002 94630 5016 94682
rect 5040 94630 5054 94682
rect 5054 94630 5066 94682
rect 5066 94630 5096 94682
rect 5120 94630 5130 94682
rect 5130 94630 5176 94682
rect 4880 94628 4936 94630
rect 4960 94628 5016 94630
rect 5040 94628 5096 94630
rect 5120 94628 5176 94630
rect 4220 94138 4276 94140
rect 4300 94138 4356 94140
rect 4380 94138 4436 94140
rect 4460 94138 4516 94140
rect 4220 94086 4266 94138
rect 4266 94086 4276 94138
rect 4300 94086 4330 94138
rect 4330 94086 4342 94138
rect 4342 94086 4356 94138
rect 4380 94086 4394 94138
rect 4394 94086 4406 94138
rect 4406 94086 4436 94138
rect 4460 94086 4470 94138
rect 4470 94086 4516 94138
rect 4220 94084 4276 94086
rect 4300 94084 4356 94086
rect 4380 94084 4436 94086
rect 4460 94084 4516 94086
rect 4880 93594 4936 93596
rect 4960 93594 5016 93596
rect 5040 93594 5096 93596
rect 5120 93594 5176 93596
rect 4880 93542 4926 93594
rect 4926 93542 4936 93594
rect 4960 93542 4990 93594
rect 4990 93542 5002 93594
rect 5002 93542 5016 93594
rect 5040 93542 5054 93594
rect 5054 93542 5066 93594
rect 5066 93542 5096 93594
rect 5120 93542 5130 93594
rect 5130 93542 5176 93594
rect 4880 93540 4936 93542
rect 4960 93540 5016 93542
rect 5040 93540 5096 93542
rect 5120 93540 5176 93542
rect 4220 93050 4276 93052
rect 4300 93050 4356 93052
rect 4380 93050 4436 93052
rect 4460 93050 4516 93052
rect 4220 92998 4266 93050
rect 4266 92998 4276 93050
rect 4300 92998 4330 93050
rect 4330 92998 4342 93050
rect 4342 92998 4356 93050
rect 4380 92998 4394 93050
rect 4394 92998 4406 93050
rect 4406 92998 4436 93050
rect 4460 92998 4470 93050
rect 4470 92998 4516 93050
rect 4220 92996 4276 92998
rect 4300 92996 4356 92998
rect 4380 92996 4436 92998
rect 4460 92996 4516 92998
rect 4880 92506 4936 92508
rect 4960 92506 5016 92508
rect 5040 92506 5096 92508
rect 5120 92506 5176 92508
rect 4880 92454 4926 92506
rect 4926 92454 4936 92506
rect 4960 92454 4990 92506
rect 4990 92454 5002 92506
rect 5002 92454 5016 92506
rect 5040 92454 5054 92506
rect 5054 92454 5066 92506
rect 5066 92454 5096 92506
rect 5120 92454 5130 92506
rect 5130 92454 5176 92506
rect 4880 92452 4936 92454
rect 4960 92452 5016 92454
rect 5040 92452 5096 92454
rect 5120 92452 5176 92454
rect 4220 91962 4276 91964
rect 4300 91962 4356 91964
rect 4380 91962 4436 91964
rect 4460 91962 4516 91964
rect 4220 91910 4266 91962
rect 4266 91910 4276 91962
rect 4300 91910 4330 91962
rect 4330 91910 4342 91962
rect 4342 91910 4356 91962
rect 4380 91910 4394 91962
rect 4394 91910 4406 91962
rect 4406 91910 4436 91962
rect 4460 91910 4470 91962
rect 4470 91910 4516 91962
rect 4220 91908 4276 91910
rect 4300 91908 4356 91910
rect 4380 91908 4436 91910
rect 4460 91908 4516 91910
rect 4880 91418 4936 91420
rect 4960 91418 5016 91420
rect 5040 91418 5096 91420
rect 5120 91418 5176 91420
rect 4880 91366 4926 91418
rect 4926 91366 4936 91418
rect 4960 91366 4990 91418
rect 4990 91366 5002 91418
rect 5002 91366 5016 91418
rect 5040 91366 5054 91418
rect 5054 91366 5066 91418
rect 5066 91366 5096 91418
rect 5120 91366 5130 91418
rect 5130 91366 5176 91418
rect 4880 91364 4936 91366
rect 4960 91364 5016 91366
rect 5040 91364 5096 91366
rect 5120 91364 5176 91366
rect 4220 90874 4276 90876
rect 4300 90874 4356 90876
rect 4380 90874 4436 90876
rect 4460 90874 4516 90876
rect 4220 90822 4266 90874
rect 4266 90822 4276 90874
rect 4300 90822 4330 90874
rect 4330 90822 4342 90874
rect 4342 90822 4356 90874
rect 4380 90822 4394 90874
rect 4394 90822 4406 90874
rect 4406 90822 4436 90874
rect 4460 90822 4470 90874
rect 4470 90822 4516 90874
rect 4220 90820 4276 90822
rect 4300 90820 4356 90822
rect 4380 90820 4436 90822
rect 4460 90820 4516 90822
rect 4880 90330 4936 90332
rect 4960 90330 5016 90332
rect 5040 90330 5096 90332
rect 5120 90330 5176 90332
rect 4880 90278 4926 90330
rect 4926 90278 4936 90330
rect 4960 90278 4990 90330
rect 4990 90278 5002 90330
rect 5002 90278 5016 90330
rect 5040 90278 5054 90330
rect 5054 90278 5066 90330
rect 5066 90278 5096 90330
rect 5120 90278 5130 90330
rect 5130 90278 5176 90330
rect 4880 90276 4936 90278
rect 4960 90276 5016 90278
rect 5040 90276 5096 90278
rect 5120 90276 5176 90278
rect 4220 89786 4276 89788
rect 4300 89786 4356 89788
rect 4380 89786 4436 89788
rect 4460 89786 4516 89788
rect 4220 89734 4266 89786
rect 4266 89734 4276 89786
rect 4300 89734 4330 89786
rect 4330 89734 4342 89786
rect 4342 89734 4356 89786
rect 4380 89734 4394 89786
rect 4394 89734 4406 89786
rect 4406 89734 4436 89786
rect 4460 89734 4470 89786
rect 4470 89734 4516 89786
rect 4220 89732 4276 89734
rect 4300 89732 4356 89734
rect 4380 89732 4436 89734
rect 4460 89732 4516 89734
rect 4880 89242 4936 89244
rect 4960 89242 5016 89244
rect 5040 89242 5096 89244
rect 5120 89242 5176 89244
rect 4880 89190 4926 89242
rect 4926 89190 4936 89242
rect 4960 89190 4990 89242
rect 4990 89190 5002 89242
rect 5002 89190 5016 89242
rect 5040 89190 5054 89242
rect 5054 89190 5066 89242
rect 5066 89190 5096 89242
rect 5120 89190 5130 89242
rect 5130 89190 5176 89242
rect 4880 89188 4936 89190
rect 4960 89188 5016 89190
rect 5040 89188 5096 89190
rect 5120 89188 5176 89190
rect 4220 88698 4276 88700
rect 4300 88698 4356 88700
rect 4380 88698 4436 88700
rect 4460 88698 4516 88700
rect 4220 88646 4266 88698
rect 4266 88646 4276 88698
rect 4300 88646 4330 88698
rect 4330 88646 4342 88698
rect 4342 88646 4356 88698
rect 4380 88646 4394 88698
rect 4394 88646 4406 88698
rect 4406 88646 4436 88698
rect 4460 88646 4470 88698
rect 4470 88646 4516 88698
rect 4220 88644 4276 88646
rect 4300 88644 4356 88646
rect 4380 88644 4436 88646
rect 4460 88644 4516 88646
rect 1306 88440 1362 88496
rect 4880 88154 4936 88156
rect 4960 88154 5016 88156
rect 5040 88154 5096 88156
rect 5120 88154 5176 88156
rect 4880 88102 4926 88154
rect 4926 88102 4936 88154
rect 4960 88102 4990 88154
rect 4990 88102 5002 88154
rect 5002 88102 5016 88154
rect 5040 88102 5054 88154
rect 5054 88102 5066 88154
rect 5066 88102 5096 88154
rect 5120 88102 5130 88154
rect 5130 88102 5176 88154
rect 4880 88100 4936 88102
rect 4960 88100 5016 88102
rect 5040 88100 5096 88102
rect 5120 88100 5176 88102
rect 1214 87760 1270 87816
rect 4220 87610 4276 87612
rect 4300 87610 4356 87612
rect 4380 87610 4436 87612
rect 4460 87610 4516 87612
rect 4220 87558 4266 87610
rect 4266 87558 4276 87610
rect 4300 87558 4330 87610
rect 4330 87558 4342 87610
rect 4342 87558 4356 87610
rect 4380 87558 4394 87610
rect 4394 87558 4406 87610
rect 4406 87558 4436 87610
rect 4460 87558 4470 87610
rect 4470 87558 4516 87610
rect 4220 87556 4276 87558
rect 4300 87556 4356 87558
rect 4380 87556 4436 87558
rect 4460 87556 4516 87558
rect 1214 87080 1270 87136
rect 1306 86400 1362 86456
rect 1306 85720 1362 85776
rect 4880 87066 4936 87068
rect 4960 87066 5016 87068
rect 5040 87066 5096 87068
rect 5120 87066 5176 87068
rect 4880 87014 4926 87066
rect 4926 87014 4936 87066
rect 4960 87014 4990 87066
rect 4990 87014 5002 87066
rect 5002 87014 5016 87066
rect 5040 87014 5054 87066
rect 5054 87014 5066 87066
rect 5066 87014 5096 87066
rect 5120 87014 5130 87066
rect 5130 87014 5176 87066
rect 4880 87012 4936 87014
rect 4960 87012 5016 87014
rect 5040 87012 5096 87014
rect 5120 87012 5176 87014
rect 4220 86522 4276 86524
rect 4300 86522 4356 86524
rect 4380 86522 4436 86524
rect 4460 86522 4516 86524
rect 4220 86470 4266 86522
rect 4266 86470 4276 86522
rect 4300 86470 4330 86522
rect 4330 86470 4342 86522
rect 4342 86470 4356 86522
rect 4380 86470 4394 86522
rect 4394 86470 4406 86522
rect 4406 86470 4436 86522
rect 4460 86470 4470 86522
rect 4470 86470 4516 86522
rect 4220 86468 4276 86470
rect 4300 86468 4356 86470
rect 4380 86468 4436 86470
rect 4460 86468 4516 86470
rect 4880 85978 4936 85980
rect 4960 85978 5016 85980
rect 5040 85978 5096 85980
rect 5120 85978 5176 85980
rect 4880 85926 4926 85978
rect 4926 85926 4936 85978
rect 4960 85926 4990 85978
rect 4990 85926 5002 85978
rect 5002 85926 5016 85978
rect 5040 85926 5054 85978
rect 5054 85926 5066 85978
rect 5066 85926 5096 85978
rect 5120 85926 5130 85978
rect 5130 85926 5176 85978
rect 4880 85924 4936 85926
rect 4960 85924 5016 85926
rect 5040 85924 5096 85926
rect 5120 85924 5176 85926
rect 5538 85448 5594 85504
rect 4220 85434 4276 85436
rect 4300 85434 4356 85436
rect 4380 85434 4436 85436
rect 4460 85434 4516 85436
rect 4220 85382 4266 85434
rect 4266 85382 4276 85434
rect 4300 85382 4330 85434
rect 4330 85382 4342 85434
rect 4342 85382 4356 85434
rect 4380 85382 4394 85434
rect 4394 85382 4406 85434
rect 4406 85382 4436 85434
rect 4460 85382 4470 85434
rect 4470 85382 4516 85434
rect 4220 85380 4276 85382
rect 4300 85380 4356 85382
rect 4380 85380 4436 85382
rect 4460 85380 4516 85382
rect 1214 85060 1270 85096
rect 1214 85040 1216 85060
rect 1216 85040 1268 85060
rect 1268 85040 1270 85060
rect 1306 84360 1362 84416
rect 1306 83680 1362 83736
rect 4880 84890 4936 84892
rect 4960 84890 5016 84892
rect 5040 84890 5096 84892
rect 5120 84890 5176 84892
rect 4880 84838 4926 84890
rect 4926 84838 4936 84890
rect 4960 84838 4990 84890
rect 4990 84838 5002 84890
rect 5002 84838 5016 84890
rect 5040 84838 5054 84890
rect 5054 84838 5066 84890
rect 5066 84838 5096 84890
rect 5120 84838 5130 84890
rect 5130 84838 5176 84890
rect 4880 84836 4936 84838
rect 4960 84836 5016 84838
rect 5040 84836 5096 84838
rect 5120 84836 5176 84838
rect 4220 84346 4276 84348
rect 4300 84346 4356 84348
rect 4380 84346 4436 84348
rect 4460 84346 4516 84348
rect 4220 84294 4266 84346
rect 4266 84294 4276 84346
rect 4300 84294 4330 84346
rect 4330 84294 4342 84346
rect 4342 84294 4356 84346
rect 4380 84294 4394 84346
rect 4394 84294 4406 84346
rect 4406 84294 4436 84346
rect 4460 84294 4470 84346
rect 4470 84294 4516 84346
rect 4220 84292 4276 84294
rect 4300 84292 4356 84294
rect 4380 84292 4436 84294
rect 4460 84292 4516 84294
rect 1306 83000 1362 83056
rect 1214 82320 1270 82376
rect 1214 81640 1270 81696
rect 1306 80960 1362 81016
rect 4880 83802 4936 83804
rect 4960 83802 5016 83804
rect 5040 83802 5096 83804
rect 5120 83802 5176 83804
rect 4880 83750 4926 83802
rect 4926 83750 4936 83802
rect 4960 83750 4990 83802
rect 4990 83750 5002 83802
rect 5002 83750 5016 83802
rect 5040 83750 5054 83802
rect 5054 83750 5066 83802
rect 5066 83750 5096 83802
rect 5120 83750 5130 83802
rect 5130 83750 5176 83802
rect 4880 83748 4936 83750
rect 4960 83748 5016 83750
rect 5040 83748 5096 83750
rect 5120 83748 5176 83750
rect 4220 83258 4276 83260
rect 4300 83258 4356 83260
rect 4380 83258 4436 83260
rect 4460 83258 4516 83260
rect 4220 83206 4266 83258
rect 4266 83206 4276 83258
rect 4300 83206 4330 83258
rect 4330 83206 4342 83258
rect 4342 83206 4356 83258
rect 4380 83206 4394 83258
rect 4394 83206 4406 83258
rect 4406 83206 4436 83258
rect 4460 83206 4470 83258
rect 4470 83206 4516 83258
rect 4220 83204 4276 83206
rect 4300 83204 4356 83206
rect 4380 83204 4436 83206
rect 4460 83204 4516 83206
rect 4880 82714 4936 82716
rect 4960 82714 5016 82716
rect 5040 82714 5096 82716
rect 5120 82714 5176 82716
rect 4880 82662 4926 82714
rect 4926 82662 4936 82714
rect 4960 82662 4990 82714
rect 4990 82662 5002 82714
rect 5002 82662 5016 82714
rect 5040 82662 5054 82714
rect 5054 82662 5066 82714
rect 5066 82662 5096 82714
rect 5120 82662 5130 82714
rect 5130 82662 5176 82714
rect 4880 82660 4936 82662
rect 4960 82660 5016 82662
rect 5040 82660 5096 82662
rect 5120 82660 5176 82662
rect 4220 82170 4276 82172
rect 4300 82170 4356 82172
rect 4380 82170 4436 82172
rect 4460 82170 4516 82172
rect 4220 82118 4266 82170
rect 4266 82118 4276 82170
rect 4300 82118 4330 82170
rect 4330 82118 4342 82170
rect 4342 82118 4356 82170
rect 4380 82118 4394 82170
rect 4394 82118 4406 82170
rect 4406 82118 4436 82170
rect 4460 82118 4470 82170
rect 4470 82118 4516 82170
rect 4220 82116 4276 82118
rect 4300 82116 4356 82118
rect 4380 82116 4436 82118
rect 4460 82116 4516 82118
rect 4880 81626 4936 81628
rect 4960 81626 5016 81628
rect 5040 81626 5096 81628
rect 5120 81626 5176 81628
rect 4880 81574 4926 81626
rect 4926 81574 4936 81626
rect 4960 81574 4990 81626
rect 4990 81574 5002 81626
rect 5002 81574 5016 81626
rect 5040 81574 5054 81626
rect 5054 81574 5066 81626
rect 5066 81574 5096 81626
rect 5120 81574 5130 81626
rect 5130 81574 5176 81626
rect 4880 81572 4936 81574
rect 4960 81572 5016 81574
rect 5040 81572 5096 81574
rect 5120 81572 5176 81574
rect 4220 81082 4276 81084
rect 4300 81082 4356 81084
rect 4380 81082 4436 81084
rect 4460 81082 4516 81084
rect 4220 81030 4266 81082
rect 4266 81030 4276 81082
rect 4300 81030 4330 81082
rect 4330 81030 4342 81082
rect 4342 81030 4356 81082
rect 4380 81030 4394 81082
rect 4394 81030 4406 81082
rect 4406 81030 4436 81082
rect 4460 81030 4470 81082
rect 4470 81030 4516 81082
rect 4220 81028 4276 81030
rect 4300 81028 4356 81030
rect 4380 81028 4436 81030
rect 4460 81028 4516 81030
rect 4880 80538 4936 80540
rect 4960 80538 5016 80540
rect 5040 80538 5096 80540
rect 5120 80538 5176 80540
rect 4880 80486 4926 80538
rect 4926 80486 4936 80538
rect 4960 80486 4990 80538
rect 4990 80486 5002 80538
rect 5002 80486 5016 80538
rect 5040 80486 5054 80538
rect 5054 80486 5066 80538
rect 5066 80486 5096 80538
rect 5120 80486 5130 80538
rect 5130 80486 5176 80538
rect 4880 80484 4936 80486
rect 4960 80484 5016 80486
rect 5040 80484 5096 80486
rect 5120 80484 5176 80486
rect 1306 80316 1308 80336
rect 1308 80316 1360 80336
rect 1360 80316 1362 80336
rect 1306 80280 1362 80316
rect 4220 79994 4276 79996
rect 4300 79994 4356 79996
rect 4380 79994 4436 79996
rect 4460 79994 4516 79996
rect 4220 79942 4266 79994
rect 4266 79942 4276 79994
rect 4300 79942 4330 79994
rect 4330 79942 4342 79994
rect 4342 79942 4356 79994
rect 4380 79942 4394 79994
rect 4394 79942 4406 79994
rect 4406 79942 4436 79994
rect 4460 79942 4470 79994
rect 4470 79942 4516 79994
rect 4220 79940 4276 79942
rect 4300 79940 4356 79942
rect 4380 79940 4436 79942
rect 4460 79940 4516 79942
rect 1214 79620 1270 79656
rect 1214 79600 1216 79620
rect 1216 79600 1268 79620
rect 1268 79600 1270 79620
rect 4880 79450 4936 79452
rect 4960 79450 5016 79452
rect 5040 79450 5096 79452
rect 5120 79450 5176 79452
rect 4880 79398 4926 79450
rect 4926 79398 4936 79450
rect 4960 79398 4990 79450
rect 4990 79398 5002 79450
rect 5002 79398 5016 79450
rect 5040 79398 5054 79450
rect 5054 79398 5066 79450
rect 5066 79398 5096 79450
rect 5120 79398 5130 79450
rect 5130 79398 5176 79450
rect 4880 79396 4936 79398
rect 4960 79396 5016 79398
rect 5040 79396 5096 79398
rect 5120 79396 5176 79398
rect 1306 78920 1362 78976
rect 4220 78906 4276 78908
rect 4300 78906 4356 78908
rect 4380 78906 4436 78908
rect 4460 78906 4516 78908
rect 4220 78854 4266 78906
rect 4266 78854 4276 78906
rect 4300 78854 4330 78906
rect 4330 78854 4342 78906
rect 4342 78854 4356 78906
rect 4380 78854 4394 78906
rect 4394 78854 4406 78906
rect 4406 78854 4436 78906
rect 4460 78854 4470 78906
rect 4470 78854 4516 78906
rect 4220 78852 4276 78854
rect 4300 78852 4356 78854
rect 4380 78852 4436 78854
rect 4460 78852 4516 78854
rect 4880 78362 4936 78364
rect 4960 78362 5016 78364
rect 5040 78362 5096 78364
rect 5120 78362 5176 78364
rect 4880 78310 4926 78362
rect 4926 78310 4936 78362
rect 4960 78310 4990 78362
rect 4990 78310 5002 78362
rect 5002 78310 5016 78362
rect 5040 78310 5054 78362
rect 5054 78310 5066 78362
rect 5066 78310 5096 78362
rect 5120 78310 5130 78362
rect 5130 78310 5176 78362
rect 4880 78308 4936 78310
rect 4960 78308 5016 78310
rect 5040 78308 5096 78310
rect 5120 78308 5176 78310
rect 1306 78240 1362 78296
rect 1306 77560 1362 77616
rect 4220 77818 4276 77820
rect 4300 77818 4356 77820
rect 4380 77818 4436 77820
rect 4460 77818 4516 77820
rect 4220 77766 4266 77818
rect 4266 77766 4276 77818
rect 4300 77766 4330 77818
rect 4330 77766 4342 77818
rect 4342 77766 4356 77818
rect 4380 77766 4394 77818
rect 4394 77766 4406 77818
rect 4406 77766 4436 77818
rect 4460 77766 4470 77818
rect 4470 77766 4516 77818
rect 4220 77764 4276 77766
rect 4300 77764 4356 77766
rect 4380 77764 4436 77766
rect 4460 77764 4516 77766
rect 4880 77274 4936 77276
rect 4960 77274 5016 77276
rect 5040 77274 5096 77276
rect 5120 77274 5176 77276
rect 4880 77222 4926 77274
rect 4926 77222 4936 77274
rect 4960 77222 4990 77274
rect 4990 77222 5002 77274
rect 5002 77222 5016 77274
rect 5040 77222 5054 77274
rect 5054 77222 5066 77274
rect 5066 77222 5096 77274
rect 5120 77222 5130 77274
rect 5130 77222 5176 77274
rect 4880 77220 4936 77222
rect 4960 77220 5016 77222
rect 5040 77220 5096 77222
rect 5120 77220 5176 77222
rect 1214 76880 1270 76936
rect 4220 76730 4276 76732
rect 4300 76730 4356 76732
rect 4380 76730 4436 76732
rect 4460 76730 4516 76732
rect 4220 76678 4266 76730
rect 4266 76678 4276 76730
rect 4300 76678 4330 76730
rect 4330 76678 4342 76730
rect 4342 76678 4356 76730
rect 4380 76678 4394 76730
rect 4394 76678 4406 76730
rect 4406 76678 4436 76730
rect 4460 76678 4470 76730
rect 4470 76678 4516 76730
rect 4220 76676 4276 76678
rect 4300 76676 4356 76678
rect 4380 76676 4436 76678
rect 4460 76676 4516 76678
rect 846 76336 902 76392
rect 4880 76186 4936 76188
rect 4960 76186 5016 76188
rect 5040 76186 5096 76188
rect 5120 76186 5176 76188
rect 4880 76134 4926 76186
rect 4926 76134 4936 76186
rect 4960 76134 4990 76186
rect 4990 76134 5002 76186
rect 5002 76134 5016 76186
rect 5040 76134 5054 76186
rect 5054 76134 5066 76186
rect 5066 76134 5096 76186
rect 5120 76134 5130 76186
rect 5130 76134 5176 76186
rect 4880 76132 4936 76134
rect 4960 76132 5016 76134
rect 5040 76132 5096 76134
rect 5120 76132 5176 76134
rect 4220 75642 4276 75644
rect 4300 75642 4356 75644
rect 4380 75642 4436 75644
rect 4460 75642 4516 75644
rect 4220 75590 4266 75642
rect 4266 75590 4276 75642
rect 4300 75590 4330 75642
rect 4330 75590 4342 75642
rect 4342 75590 4356 75642
rect 4380 75590 4394 75642
rect 4394 75590 4406 75642
rect 4406 75590 4436 75642
rect 4460 75590 4470 75642
rect 4470 75590 4516 75642
rect 4220 75588 4276 75590
rect 4300 75588 4356 75590
rect 4380 75588 4436 75590
rect 4460 75588 4516 75590
rect 1490 75520 1546 75576
rect 4880 75098 4936 75100
rect 4960 75098 5016 75100
rect 5040 75098 5096 75100
rect 5120 75098 5176 75100
rect 4880 75046 4926 75098
rect 4926 75046 4936 75098
rect 4960 75046 4990 75098
rect 4990 75046 5002 75098
rect 5002 75046 5016 75098
rect 5040 75046 5054 75098
rect 5054 75046 5066 75098
rect 5066 75046 5096 75098
rect 5120 75046 5130 75098
rect 5130 75046 5176 75098
rect 4880 75044 4936 75046
rect 4960 75044 5016 75046
rect 5040 75044 5096 75046
rect 5120 75044 5176 75046
rect 846 74976 902 75032
rect 4220 74554 4276 74556
rect 4300 74554 4356 74556
rect 4380 74554 4436 74556
rect 4460 74554 4516 74556
rect 4220 74502 4266 74554
rect 4266 74502 4276 74554
rect 4300 74502 4330 74554
rect 4330 74502 4342 74554
rect 4342 74502 4356 74554
rect 4380 74502 4394 74554
rect 4394 74502 4406 74554
rect 4406 74502 4436 74554
rect 4460 74502 4470 74554
rect 4470 74502 4516 74554
rect 4220 74500 4276 74502
rect 4300 74500 4356 74502
rect 4380 74500 4436 74502
rect 4460 74500 4516 74502
rect 846 74332 848 74352
rect 848 74332 900 74352
rect 900 74332 902 74352
rect 846 74296 902 74332
rect 4880 74010 4936 74012
rect 4960 74010 5016 74012
rect 5040 74010 5096 74012
rect 5120 74010 5176 74012
rect 4880 73958 4926 74010
rect 4926 73958 4936 74010
rect 4960 73958 4990 74010
rect 4990 73958 5002 74010
rect 5002 73958 5016 74010
rect 5040 73958 5054 74010
rect 5054 73958 5066 74010
rect 5066 73958 5096 74010
rect 5120 73958 5130 74010
rect 5130 73958 5176 74010
rect 4880 73956 4936 73958
rect 4960 73956 5016 73958
rect 5040 73956 5096 73958
rect 5120 73956 5176 73958
rect 846 73636 902 73672
rect 846 73616 848 73636
rect 848 73616 900 73636
rect 900 73616 902 73636
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 846 72972 848 72992
rect 848 72972 900 72992
rect 900 72972 902 72992
rect 846 72936 902 72972
rect 4880 72922 4936 72924
rect 4960 72922 5016 72924
rect 5040 72922 5096 72924
rect 5120 72922 5176 72924
rect 4880 72870 4926 72922
rect 4926 72870 4936 72922
rect 4960 72870 4990 72922
rect 4990 72870 5002 72922
rect 5002 72870 5016 72922
rect 5040 72870 5054 72922
rect 5054 72870 5066 72922
rect 5066 72870 5096 72922
rect 5120 72870 5130 72922
rect 5130 72870 5176 72922
rect 4880 72868 4936 72870
rect 4960 72868 5016 72870
rect 5040 72868 5096 72870
rect 5120 72868 5176 72870
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 846 72256 902 72312
rect 4880 71834 4936 71836
rect 4960 71834 5016 71836
rect 5040 71834 5096 71836
rect 5120 71834 5176 71836
rect 4880 71782 4926 71834
rect 4926 71782 4936 71834
rect 4960 71782 4990 71834
rect 4990 71782 5002 71834
rect 5002 71782 5016 71834
rect 5040 71782 5054 71834
rect 5054 71782 5066 71834
rect 5066 71782 5096 71834
rect 5120 71782 5130 71834
rect 5130 71782 5176 71834
rect 4880 71780 4936 71782
rect 4960 71780 5016 71782
rect 5040 71780 5096 71782
rect 5120 71780 5176 71782
rect 1214 71440 1270 71496
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 5538 79464 5594 79520
rect 7470 79872 7526 79928
rect 9494 111196 9550 111252
rect 9494 109540 9550 109552
rect 9494 109496 9496 109540
rect 9496 109496 9548 109540
rect 9548 109496 9550 109540
rect 9494 108400 9496 108424
rect 9496 108400 9548 108424
rect 9548 108400 9550 108424
rect 9494 108368 9550 108400
rect 9494 106668 9550 106724
rect 9494 105585 9550 105641
rect 9494 103905 9550 103961
rect 8390 79600 8446 79656
rect 35600 136026 35656 136028
rect 35680 136026 35736 136028
rect 35760 136026 35816 136028
rect 35840 136026 35896 136028
rect 35600 135974 35646 136026
rect 35646 135974 35656 136026
rect 35680 135974 35710 136026
rect 35710 135974 35722 136026
rect 35722 135974 35736 136026
rect 35760 135974 35774 136026
rect 35774 135974 35786 136026
rect 35786 135974 35816 136026
rect 35840 135974 35850 136026
rect 35850 135974 35896 136026
rect 35600 135972 35656 135974
rect 35680 135972 35736 135974
rect 35760 135972 35816 135974
rect 35840 135972 35896 135974
rect 38750 134136 38806 134192
rect 43166 134136 43222 134192
rect 65660 136570 65716 136572
rect 65740 136570 65796 136572
rect 65820 136570 65876 136572
rect 65900 136570 65956 136572
rect 65660 136518 65706 136570
rect 65706 136518 65716 136570
rect 65740 136518 65770 136570
rect 65770 136518 65782 136570
rect 65782 136518 65796 136570
rect 65820 136518 65834 136570
rect 65834 136518 65846 136570
rect 65846 136518 65876 136570
rect 65900 136518 65910 136570
rect 65910 136518 65956 136570
rect 65660 136516 65716 136518
rect 65740 136516 65796 136518
rect 65820 136516 65876 136518
rect 65900 136516 65956 136518
rect 60554 135224 60610 135280
rect 63130 135224 63186 135280
rect 66320 136026 66376 136028
rect 66400 136026 66456 136028
rect 66480 136026 66536 136028
rect 66560 136026 66616 136028
rect 66320 135974 66366 136026
rect 66366 135974 66376 136026
rect 66400 135974 66430 136026
rect 66430 135974 66442 136026
rect 66442 135974 66456 136026
rect 66480 135974 66494 136026
rect 66494 135974 66506 136026
rect 66506 135974 66536 136026
rect 66560 135974 66570 136026
rect 66570 135974 66616 136026
rect 66320 135972 66376 135974
rect 66400 135972 66456 135974
rect 66480 135972 66536 135974
rect 66560 135972 66616 135974
rect 63590 135088 63646 135144
rect 55402 134136 55458 134192
rect 57978 134136 58034 134192
rect 72698 135224 72754 135280
rect 96380 136570 96436 136572
rect 96460 136570 96516 136572
rect 96540 136570 96596 136572
rect 96620 136570 96676 136572
rect 96380 136518 96426 136570
rect 96426 136518 96436 136570
rect 96460 136518 96490 136570
rect 96490 136518 96502 136570
rect 96502 136518 96516 136570
rect 96540 136518 96554 136570
rect 96554 136518 96566 136570
rect 96566 136518 96596 136570
rect 96620 136518 96630 136570
rect 96630 136518 96676 136570
rect 96380 136516 96436 136518
rect 96460 136516 96516 136518
rect 96540 136516 96596 136518
rect 96620 136516 96676 136518
rect 77390 134408 77446 134464
rect 72514 134136 72570 134192
rect 97040 136026 97096 136028
rect 97120 136026 97176 136028
rect 97200 136026 97256 136028
rect 97280 136026 97336 136028
rect 97040 135974 97086 136026
rect 97086 135974 97096 136026
rect 97120 135974 97150 136026
rect 97150 135974 97162 136026
rect 97162 135974 97176 136026
rect 97200 135974 97214 136026
rect 97214 135974 97226 136026
rect 97226 135974 97256 136026
rect 97280 135974 97290 136026
rect 97290 135974 97336 136026
rect 97040 135972 97096 135974
rect 97120 135972 97176 135974
rect 97200 135972 97256 135974
rect 97280 135972 97336 135974
rect 95974 135632 96030 135688
rect 36082 133864 36138 133920
rect 38566 133864 38622 133920
rect 46110 133864 46166 133920
rect 48502 133864 48558 133920
rect 51078 133864 51134 133920
rect 68558 133864 68614 133920
rect 86314 133864 86370 133920
rect 87326 133900 87328 133920
rect 87328 133900 87380 133920
rect 87380 133900 87382 133920
rect 87326 133864 87382 133900
rect 102046 92204 102102 92260
rect 9310 79192 9366 79248
rect 9218 79056 9274 79112
rect 9586 79736 9642 79792
rect 16118 79872 16174 79928
rect 23478 79872 23534 79928
rect 36266 79872 36322 79928
rect 39762 79892 39818 79928
rect 39762 79872 39764 79892
rect 39764 79872 39816 79892
rect 39816 79872 39818 79892
rect 4880 70746 4936 70748
rect 4960 70746 5016 70748
rect 5040 70746 5096 70748
rect 5120 70746 5176 70748
rect 4880 70694 4926 70746
rect 4926 70694 4936 70746
rect 4960 70694 4990 70746
rect 4990 70694 5002 70746
rect 5002 70694 5016 70746
rect 5040 70694 5054 70746
rect 5054 70694 5066 70746
rect 5066 70694 5096 70746
rect 5120 70694 5130 70746
rect 5130 70694 5176 70746
rect 4880 70692 4936 70694
rect 4960 70692 5016 70694
rect 5040 70692 5096 70694
rect 5120 70692 5176 70694
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 4880 69658 4936 69660
rect 4960 69658 5016 69660
rect 5040 69658 5096 69660
rect 5120 69658 5176 69660
rect 4880 69606 4926 69658
rect 4926 69606 4936 69658
rect 4960 69606 4990 69658
rect 4990 69606 5002 69658
rect 5002 69606 5016 69658
rect 5040 69606 5054 69658
rect 5054 69606 5066 69658
rect 5066 69606 5096 69658
rect 5120 69606 5130 69658
rect 5130 69606 5176 69658
rect 4880 69604 4936 69606
rect 4960 69604 5016 69606
rect 5040 69604 5096 69606
rect 5120 69604 5176 69606
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 4880 68570 4936 68572
rect 4960 68570 5016 68572
rect 5040 68570 5096 68572
rect 5120 68570 5176 68572
rect 4880 68518 4926 68570
rect 4926 68518 4936 68570
rect 4960 68518 4990 68570
rect 4990 68518 5002 68570
rect 5002 68518 5016 68570
rect 5040 68518 5054 68570
rect 5054 68518 5066 68570
rect 5066 68518 5096 68570
rect 5120 68518 5130 68570
rect 5130 68518 5176 68570
rect 4880 68516 4936 68518
rect 4960 68516 5016 68518
rect 5040 68516 5096 68518
rect 5120 68516 5176 68518
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 4880 67482 4936 67484
rect 4960 67482 5016 67484
rect 5040 67482 5096 67484
rect 5120 67482 5176 67484
rect 4880 67430 4926 67482
rect 4926 67430 4936 67482
rect 4960 67430 4990 67482
rect 4990 67430 5002 67482
rect 5002 67430 5016 67482
rect 5040 67430 5054 67482
rect 5054 67430 5066 67482
rect 5066 67430 5096 67482
rect 5120 67430 5130 67482
rect 5130 67430 5176 67482
rect 4880 67428 4936 67430
rect 4960 67428 5016 67430
rect 5040 67428 5096 67430
rect 5120 67428 5176 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 4880 66394 4936 66396
rect 4960 66394 5016 66396
rect 5040 66394 5096 66396
rect 5120 66394 5176 66396
rect 4880 66342 4926 66394
rect 4926 66342 4936 66394
rect 4960 66342 4990 66394
rect 4990 66342 5002 66394
rect 5002 66342 5016 66394
rect 5040 66342 5054 66394
rect 5054 66342 5066 66394
rect 5066 66342 5096 66394
rect 5120 66342 5130 66394
rect 5130 66342 5176 66394
rect 4880 66340 4936 66342
rect 4960 66340 5016 66342
rect 5040 66340 5096 66342
rect 5120 66340 5176 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 4880 65306 4936 65308
rect 4960 65306 5016 65308
rect 5040 65306 5096 65308
rect 5120 65306 5176 65308
rect 4880 65254 4926 65306
rect 4926 65254 4936 65306
rect 4960 65254 4990 65306
rect 4990 65254 5002 65306
rect 5002 65254 5016 65306
rect 5040 65254 5054 65306
rect 5054 65254 5066 65306
rect 5066 65254 5096 65306
rect 5120 65254 5130 65306
rect 5130 65254 5176 65306
rect 4880 65252 4936 65254
rect 4960 65252 5016 65254
rect 5040 65252 5096 65254
rect 5120 65252 5176 65254
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4880 64218 4936 64220
rect 4960 64218 5016 64220
rect 5040 64218 5096 64220
rect 5120 64218 5176 64220
rect 4880 64166 4926 64218
rect 4926 64166 4936 64218
rect 4960 64166 4990 64218
rect 4990 64166 5002 64218
rect 5002 64166 5016 64218
rect 5040 64166 5054 64218
rect 5054 64166 5066 64218
rect 5066 64166 5096 64218
rect 5120 64166 5130 64218
rect 5130 64166 5176 64218
rect 4880 64164 4936 64166
rect 4960 64164 5016 64166
rect 5040 64164 5096 64166
rect 5120 64164 5176 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4880 63130 4936 63132
rect 4960 63130 5016 63132
rect 5040 63130 5096 63132
rect 5120 63130 5176 63132
rect 4880 63078 4926 63130
rect 4926 63078 4936 63130
rect 4960 63078 4990 63130
rect 4990 63078 5002 63130
rect 5002 63078 5016 63130
rect 5040 63078 5054 63130
rect 5054 63078 5066 63130
rect 5066 63078 5096 63130
rect 5120 63078 5130 63130
rect 5130 63078 5176 63130
rect 4880 63076 4936 63078
rect 4960 63076 5016 63078
rect 5040 63076 5096 63078
rect 5120 63076 5176 63078
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4880 62042 4936 62044
rect 4960 62042 5016 62044
rect 5040 62042 5096 62044
rect 5120 62042 5176 62044
rect 4880 61990 4926 62042
rect 4926 61990 4936 62042
rect 4960 61990 4990 62042
rect 4990 61990 5002 62042
rect 5002 61990 5016 62042
rect 5040 61990 5054 62042
rect 5054 61990 5066 62042
rect 5066 61990 5096 62042
rect 5120 61990 5130 62042
rect 5130 61990 5176 62042
rect 4880 61988 4936 61990
rect 4960 61988 5016 61990
rect 5040 61988 5096 61990
rect 5120 61988 5176 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4880 60954 4936 60956
rect 4960 60954 5016 60956
rect 5040 60954 5096 60956
rect 5120 60954 5176 60956
rect 4880 60902 4926 60954
rect 4926 60902 4936 60954
rect 4960 60902 4990 60954
rect 4990 60902 5002 60954
rect 5002 60902 5016 60954
rect 5040 60902 5054 60954
rect 5054 60902 5066 60954
rect 5066 60902 5096 60954
rect 5120 60902 5130 60954
rect 5130 60902 5176 60954
rect 4880 60900 4936 60902
rect 4960 60900 5016 60902
rect 5040 60900 5096 60902
rect 5120 60900 5176 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4880 59866 4936 59868
rect 4960 59866 5016 59868
rect 5040 59866 5096 59868
rect 5120 59866 5176 59868
rect 4880 59814 4926 59866
rect 4926 59814 4936 59866
rect 4960 59814 4990 59866
rect 4990 59814 5002 59866
rect 5002 59814 5016 59866
rect 5040 59814 5054 59866
rect 5054 59814 5066 59866
rect 5066 59814 5096 59866
rect 5120 59814 5130 59866
rect 5130 59814 5176 59866
rect 4880 59812 4936 59814
rect 4960 59812 5016 59814
rect 5040 59812 5096 59814
rect 5120 59812 5176 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4880 58778 4936 58780
rect 4960 58778 5016 58780
rect 5040 58778 5096 58780
rect 5120 58778 5176 58780
rect 4880 58726 4926 58778
rect 4926 58726 4936 58778
rect 4960 58726 4990 58778
rect 4990 58726 5002 58778
rect 5002 58726 5016 58778
rect 5040 58726 5054 58778
rect 5054 58726 5066 58778
rect 5066 58726 5096 58778
rect 5120 58726 5130 58778
rect 5130 58726 5176 58778
rect 4880 58724 4936 58726
rect 4960 58724 5016 58726
rect 5040 58724 5096 58726
rect 5120 58724 5176 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 7562 41248 7618 41304
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 1490 13640 1546 13696
rect 1306 12960 1362 13016
rect 1490 12280 1546 12336
rect 1214 11600 1270 11656
rect 1490 10920 1546 10976
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 7286 39480 7342 39536
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 7562 38392 7618 38448
rect 7562 36644 7618 36680
rect 7562 36624 7564 36644
rect 7564 36624 7616 36644
rect 7616 36624 7618 36644
rect 7470 35536 7526 35592
rect 7562 33924 7618 33960
rect 7562 33904 7564 33924
rect 7564 33904 7616 33924
rect 7616 33904 7618 33924
rect 7470 15408 7526 15464
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1306 10240 1362 10296
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 1490 9560 1546 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 1214 8900 1270 8936
rect 1214 8880 1216 8900
rect 1216 8880 1268 8900
rect 1268 8880 1270 8900
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 1950 8200 2006 8256
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 1306 7520 1362 7576
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1306 6840 1362 6896
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 1214 6160 1270 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 40958 79908 40960 79928
rect 40960 79908 41012 79928
rect 41012 79908 41014 79928
rect 40958 79872 41014 79908
rect 43258 79872 43314 79928
rect 30470 79600 30526 79656
rect 31666 79620 31722 79656
rect 31666 79600 31668 79620
rect 31668 79600 31720 79620
rect 31720 79600 31722 79620
rect 24674 79464 24730 79520
rect 26054 79464 26110 79520
rect 26974 79464 27030 79520
rect 28170 79464 28226 79520
rect 29550 79464 29606 79520
rect 26974 79192 27030 79248
rect 28170 79056 28226 79112
rect 33966 79464 34022 79520
rect 35346 79464 35402 79520
rect 32862 79056 32918 79112
rect 34940 77818 34996 77820
rect 35020 77818 35076 77820
rect 35100 77818 35156 77820
rect 35180 77818 35236 77820
rect 34940 77766 34986 77818
rect 34986 77766 34996 77818
rect 35020 77766 35050 77818
rect 35050 77766 35062 77818
rect 35062 77766 35076 77818
rect 35100 77766 35114 77818
rect 35114 77766 35126 77818
rect 35126 77766 35156 77818
rect 35180 77766 35190 77818
rect 35190 77766 35236 77818
rect 34940 77764 34996 77766
rect 35020 77764 35076 77766
rect 35100 77764 35156 77766
rect 35180 77764 35236 77766
rect 38658 79756 38714 79792
rect 38658 79736 38660 79756
rect 38660 79736 38712 79756
rect 38712 79736 38714 79756
rect 37462 79600 37518 79656
rect 42154 79464 42210 79520
rect 65660 77818 65716 77820
rect 65740 77818 65796 77820
rect 65820 77818 65876 77820
rect 65900 77818 65956 77820
rect 65660 77766 65706 77818
rect 65706 77766 65716 77818
rect 65740 77766 65770 77818
rect 65770 77766 65782 77818
rect 65782 77766 65796 77818
rect 65820 77766 65834 77818
rect 65834 77766 65846 77818
rect 65846 77766 65876 77818
rect 65900 77766 65910 77818
rect 65910 77766 65956 77818
rect 65660 77764 65716 77766
rect 65740 77764 65796 77766
rect 65820 77764 65876 77766
rect 65900 77764 65956 77766
rect 35600 77274 35656 77276
rect 35680 77274 35736 77276
rect 35760 77274 35816 77276
rect 35840 77274 35896 77276
rect 35600 77222 35646 77274
rect 35646 77222 35656 77274
rect 35680 77222 35710 77274
rect 35710 77222 35722 77274
rect 35722 77222 35736 77274
rect 35760 77222 35774 77274
rect 35774 77222 35786 77274
rect 35786 77222 35816 77274
rect 35840 77222 35850 77274
rect 35850 77222 35896 77274
rect 35600 77220 35656 77222
rect 35680 77220 35736 77222
rect 35760 77220 35816 77222
rect 35840 77220 35896 77222
rect 34940 76730 34996 76732
rect 35020 76730 35076 76732
rect 35100 76730 35156 76732
rect 35180 76730 35236 76732
rect 34940 76678 34986 76730
rect 34986 76678 34996 76730
rect 35020 76678 35050 76730
rect 35050 76678 35062 76730
rect 35062 76678 35076 76730
rect 35100 76678 35114 76730
rect 35114 76678 35126 76730
rect 35126 76678 35156 76730
rect 35180 76678 35190 76730
rect 35190 76678 35236 76730
rect 34940 76676 34996 76678
rect 35020 76676 35076 76678
rect 35100 76676 35156 76678
rect 35180 76676 35236 76678
rect 35600 76186 35656 76188
rect 35680 76186 35736 76188
rect 35760 76186 35816 76188
rect 35840 76186 35896 76188
rect 35600 76134 35646 76186
rect 35646 76134 35656 76186
rect 35680 76134 35710 76186
rect 35710 76134 35722 76186
rect 35722 76134 35736 76186
rect 35760 76134 35774 76186
rect 35774 76134 35786 76186
rect 35786 76134 35816 76186
rect 35840 76134 35850 76186
rect 35850 76134 35896 76186
rect 35600 76132 35656 76134
rect 35680 76132 35736 76134
rect 35760 76132 35816 76134
rect 35840 76132 35896 76134
rect 34940 75642 34996 75644
rect 35020 75642 35076 75644
rect 35100 75642 35156 75644
rect 35180 75642 35236 75644
rect 34940 75590 34986 75642
rect 34986 75590 34996 75642
rect 35020 75590 35050 75642
rect 35050 75590 35062 75642
rect 35062 75590 35076 75642
rect 35100 75590 35114 75642
rect 35114 75590 35126 75642
rect 35126 75590 35156 75642
rect 35180 75590 35190 75642
rect 35190 75590 35236 75642
rect 34940 75588 34996 75590
rect 35020 75588 35076 75590
rect 35100 75588 35156 75590
rect 35180 75588 35236 75590
rect 35600 75098 35656 75100
rect 35680 75098 35736 75100
rect 35760 75098 35816 75100
rect 35840 75098 35896 75100
rect 35600 75046 35646 75098
rect 35646 75046 35656 75098
rect 35680 75046 35710 75098
rect 35710 75046 35722 75098
rect 35722 75046 35736 75098
rect 35760 75046 35774 75098
rect 35774 75046 35786 75098
rect 35786 75046 35816 75098
rect 35840 75046 35850 75098
rect 35850 75046 35896 75098
rect 35600 75044 35656 75046
rect 35680 75044 35736 75046
rect 35760 75044 35816 75046
rect 35840 75044 35896 75046
rect 34940 74554 34996 74556
rect 35020 74554 35076 74556
rect 35100 74554 35156 74556
rect 35180 74554 35236 74556
rect 34940 74502 34986 74554
rect 34986 74502 34996 74554
rect 35020 74502 35050 74554
rect 35050 74502 35062 74554
rect 35062 74502 35076 74554
rect 35100 74502 35114 74554
rect 35114 74502 35126 74554
rect 35126 74502 35156 74554
rect 35180 74502 35190 74554
rect 35190 74502 35236 74554
rect 34940 74500 34996 74502
rect 35020 74500 35076 74502
rect 35100 74500 35156 74502
rect 35180 74500 35236 74502
rect 34940 73466 34996 73468
rect 35020 73466 35076 73468
rect 35100 73466 35156 73468
rect 35180 73466 35236 73468
rect 34940 73414 34986 73466
rect 34986 73414 34996 73466
rect 35020 73414 35050 73466
rect 35050 73414 35062 73466
rect 35062 73414 35076 73466
rect 35100 73414 35114 73466
rect 35114 73414 35126 73466
rect 35126 73414 35156 73466
rect 35180 73414 35190 73466
rect 35190 73414 35236 73466
rect 34940 73412 34996 73414
rect 35020 73412 35076 73414
rect 35100 73412 35156 73414
rect 35180 73412 35236 73414
rect 35600 74010 35656 74012
rect 35680 74010 35736 74012
rect 35760 74010 35816 74012
rect 35840 74010 35896 74012
rect 35600 73958 35646 74010
rect 35646 73958 35656 74010
rect 35680 73958 35710 74010
rect 35710 73958 35722 74010
rect 35722 73958 35736 74010
rect 35760 73958 35774 74010
rect 35774 73958 35786 74010
rect 35786 73958 35816 74010
rect 35840 73958 35850 74010
rect 35850 73958 35896 74010
rect 35600 73956 35656 73958
rect 35680 73956 35736 73958
rect 35760 73956 35816 73958
rect 35840 73956 35896 73958
rect 35600 72922 35656 72924
rect 35680 72922 35736 72924
rect 35760 72922 35816 72924
rect 35840 72922 35896 72924
rect 35600 72870 35646 72922
rect 35646 72870 35656 72922
rect 35680 72870 35710 72922
rect 35710 72870 35722 72922
rect 35722 72870 35736 72922
rect 35760 72870 35774 72922
rect 35774 72870 35786 72922
rect 35786 72870 35816 72922
rect 35840 72870 35850 72922
rect 35850 72870 35896 72922
rect 35600 72868 35656 72870
rect 35680 72868 35736 72870
rect 35760 72868 35816 72870
rect 35840 72868 35896 72870
rect 34940 72378 34996 72380
rect 35020 72378 35076 72380
rect 35100 72378 35156 72380
rect 35180 72378 35236 72380
rect 34940 72326 34986 72378
rect 34986 72326 34996 72378
rect 35020 72326 35050 72378
rect 35050 72326 35062 72378
rect 35062 72326 35076 72378
rect 35100 72326 35114 72378
rect 35114 72326 35126 72378
rect 35126 72326 35156 72378
rect 35180 72326 35190 72378
rect 35190 72326 35236 72378
rect 34940 72324 34996 72326
rect 35020 72324 35076 72326
rect 35100 72324 35156 72326
rect 35180 72324 35236 72326
rect 35600 71834 35656 71836
rect 35680 71834 35736 71836
rect 35760 71834 35816 71836
rect 35840 71834 35896 71836
rect 35600 71782 35646 71834
rect 35646 71782 35656 71834
rect 35680 71782 35710 71834
rect 35710 71782 35722 71834
rect 35722 71782 35736 71834
rect 35760 71782 35774 71834
rect 35774 71782 35786 71834
rect 35786 71782 35816 71834
rect 35840 71782 35850 71834
rect 35850 71782 35896 71834
rect 35600 71780 35656 71782
rect 35680 71780 35736 71782
rect 35760 71780 35816 71782
rect 35840 71780 35896 71782
rect 34940 71290 34996 71292
rect 35020 71290 35076 71292
rect 35100 71290 35156 71292
rect 35180 71290 35236 71292
rect 34940 71238 34986 71290
rect 34986 71238 34996 71290
rect 35020 71238 35050 71290
rect 35050 71238 35062 71290
rect 35062 71238 35076 71290
rect 35100 71238 35114 71290
rect 35114 71238 35126 71290
rect 35126 71238 35156 71290
rect 35180 71238 35190 71290
rect 35190 71238 35236 71290
rect 34940 71236 34996 71238
rect 35020 71236 35076 71238
rect 35100 71236 35156 71238
rect 35180 71236 35236 71238
rect 35600 70746 35656 70748
rect 35680 70746 35736 70748
rect 35760 70746 35816 70748
rect 35840 70746 35896 70748
rect 35600 70694 35646 70746
rect 35646 70694 35656 70746
rect 35680 70694 35710 70746
rect 35710 70694 35722 70746
rect 35722 70694 35736 70746
rect 35760 70694 35774 70746
rect 35774 70694 35786 70746
rect 35786 70694 35816 70746
rect 35840 70694 35850 70746
rect 35850 70694 35896 70746
rect 35600 70692 35656 70694
rect 35680 70692 35736 70694
rect 35760 70692 35816 70694
rect 35840 70692 35896 70694
rect 34940 70202 34996 70204
rect 35020 70202 35076 70204
rect 35100 70202 35156 70204
rect 35180 70202 35236 70204
rect 34940 70150 34986 70202
rect 34986 70150 34996 70202
rect 35020 70150 35050 70202
rect 35050 70150 35062 70202
rect 35062 70150 35076 70202
rect 35100 70150 35114 70202
rect 35114 70150 35126 70202
rect 35126 70150 35156 70202
rect 35180 70150 35190 70202
rect 35190 70150 35236 70202
rect 34940 70148 34996 70150
rect 35020 70148 35076 70150
rect 35100 70148 35156 70150
rect 35180 70148 35236 70150
rect 35600 69658 35656 69660
rect 35680 69658 35736 69660
rect 35760 69658 35816 69660
rect 35840 69658 35896 69660
rect 35600 69606 35646 69658
rect 35646 69606 35656 69658
rect 35680 69606 35710 69658
rect 35710 69606 35722 69658
rect 35722 69606 35736 69658
rect 35760 69606 35774 69658
rect 35774 69606 35786 69658
rect 35786 69606 35816 69658
rect 35840 69606 35850 69658
rect 35850 69606 35896 69658
rect 35600 69604 35656 69606
rect 35680 69604 35736 69606
rect 35760 69604 35816 69606
rect 35840 69604 35896 69606
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 35600 68570 35656 68572
rect 35680 68570 35736 68572
rect 35760 68570 35816 68572
rect 35840 68570 35896 68572
rect 35600 68518 35646 68570
rect 35646 68518 35656 68570
rect 35680 68518 35710 68570
rect 35710 68518 35722 68570
rect 35722 68518 35736 68570
rect 35760 68518 35774 68570
rect 35774 68518 35786 68570
rect 35786 68518 35816 68570
rect 35840 68518 35850 68570
rect 35850 68518 35896 68570
rect 35600 68516 35656 68518
rect 35680 68516 35736 68518
rect 35760 68516 35816 68518
rect 35840 68516 35896 68518
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 35600 67482 35656 67484
rect 35680 67482 35736 67484
rect 35760 67482 35816 67484
rect 35840 67482 35896 67484
rect 35600 67430 35646 67482
rect 35646 67430 35656 67482
rect 35680 67430 35710 67482
rect 35710 67430 35722 67482
rect 35722 67430 35736 67482
rect 35760 67430 35774 67482
rect 35774 67430 35786 67482
rect 35786 67430 35816 67482
rect 35840 67430 35850 67482
rect 35850 67430 35896 67482
rect 35600 67428 35656 67430
rect 35680 67428 35736 67430
rect 35760 67428 35816 67430
rect 35840 67428 35896 67430
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 35600 66394 35656 66396
rect 35680 66394 35736 66396
rect 35760 66394 35816 66396
rect 35840 66394 35896 66396
rect 35600 66342 35646 66394
rect 35646 66342 35656 66394
rect 35680 66342 35710 66394
rect 35710 66342 35722 66394
rect 35722 66342 35736 66394
rect 35760 66342 35774 66394
rect 35774 66342 35786 66394
rect 35786 66342 35816 66394
rect 35840 66342 35850 66394
rect 35850 66342 35896 66394
rect 35600 66340 35656 66342
rect 35680 66340 35736 66342
rect 35760 66340 35816 66342
rect 35840 66340 35896 66342
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 34518 65592 34574 65648
rect 31666 65456 31722 65512
rect 66320 77274 66376 77276
rect 66400 77274 66456 77276
rect 66480 77274 66536 77276
rect 66560 77274 66616 77276
rect 66320 77222 66366 77274
rect 66366 77222 66376 77274
rect 66400 77222 66430 77274
rect 66430 77222 66442 77274
rect 66442 77222 66456 77274
rect 66480 77222 66494 77274
rect 66494 77222 66506 77274
rect 66506 77222 66536 77274
rect 66560 77222 66570 77274
rect 66570 77222 66616 77274
rect 66320 77220 66376 77222
rect 66400 77220 66456 77222
rect 66480 77220 66536 77222
rect 66560 77220 66616 77222
rect 67914 77016 67970 77072
rect 65982 76880 66038 76936
rect 65660 76730 65716 76732
rect 65740 76730 65796 76732
rect 65820 76730 65876 76732
rect 65900 76730 65956 76732
rect 65660 76678 65706 76730
rect 65706 76678 65716 76730
rect 65740 76678 65770 76730
rect 65770 76678 65782 76730
rect 65782 76678 65796 76730
rect 65820 76678 65834 76730
rect 65834 76678 65846 76730
rect 65846 76678 65876 76730
rect 65900 76678 65910 76730
rect 65910 76678 65956 76730
rect 65660 76676 65716 76678
rect 65740 76676 65796 76678
rect 65820 76676 65876 76678
rect 65900 76676 65956 76678
rect 43718 68176 43774 68232
rect 63130 76472 63186 76528
rect 61014 76356 61070 76392
rect 61014 76336 61016 76356
rect 61016 76336 61068 76356
rect 61068 76336 61070 76356
rect 66320 76186 66376 76188
rect 66400 76186 66456 76188
rect 66480 76186 66536 76188
rect 66560 76186 66616 76188
rect 66320 76134 66366 76186
rect 66366 76134 66376 76186
rect 66400 76134 66430 76186
rect 66430 76134 66442 76186
rect 66442 76134 66456 76186
rect 66480 76134 66494 76186
rect 66494 76134 66506 76186
rect 66506 76134 66536 76186
rect 66560 76134 66570 76186
rect 66570 76134 66616 76186
rect 66320 76132 66376 76134
rect 66400 76132 66456 76134
rect 66480 76132 66536 76134
rect 66560 76132 66616 76134
rect 65660 75642 65716 75644
rect 65740 75642 65796 75644
rect 65820 75642 65876 75644
rect 65900 75642 65956 75644
rect 65660 75590 65706 75642
rect 65706 75590 65716 75642
rect 65740 75590 65770 75642
rect 65770 75590 65782 75642
rect 65782 75590 65796 75642
rect 65820 75590 65834 75642
rect 65834 75590 65846 75642
rect 65846 75590 65876 75642
rect 65900 75590 65910 75642
rect 65910 75590 65956 75642
rect 65660 75588 65716 75590
rect 65740 75588 65796 75590
rect 65820 75588 65876 75590
rect 65900 75588 65956 75590
rect 66320 75098 66376 75100
rect 66400 75098 66456 75100
rect 66480 75098 66536 75100
rect 66560 75098 66616 75100
rect 66320 75046 66366 75098
rect 66366 75046 66376 75098
rect 66400 75046 66430 75098
rect 66430 75046 66442 75098
rect 66442 75046 66456 75098
rect 66480 75046 66494 75098
rect 66494 75046 66506 75098
rect 66506 75046 66536 75098
rect 66560 75046 66570 75098
rect 66570 75046 66616 75098
rect 66320 75044 66376 75046
rect 66400 75044 66456 75046
rect 66480 75044 66536 75046
rect 66560 75044 66616 75046
rect 65660 74554 65716 74556
rect 65740 74554 65796 74556
rect 65820 74554 65876 74556
rect 65900 74554 65956 74556
rect 65660 74502 65706 74554
rect 65706 74502 65716 74554
rect 65740 74502 65770 74554
rect 65770 74502 65782 74554
rect 65782 74502 65796 74554
rect 65820 74502 65834 74554
rect 65834 74502 65846 74554
rect 65846 74502 65876 74554
rect 65900 74502 65910 74554
rect 65910 74502 65956 74554
rect 65660 74500 65716 74502
rect 65740 74500 65796 74502
rect 65820 74500 65876 74502
rect 65900 74500 65956 74502
rect 66320 74010 66376 74012
rect 66400 74010 66456 74012
rect 66480 74010 66536 74012
rect 66560 74010 66616 74012
rect 66320 73958 66366 74010
rect 66366 73958 66376 74010
rect 66400 73958 66430 74010
rect 66430 73958 66442 74010
rect 66442 73958 66456 74010
rect 66480 73958 66494 74010
rect 66494 73958 66506 74010
rect 66506 73958 66536 74010
rect 66560 73958 66570 74010
rect 66570 73958 66616 74010
rect 66320 73956 66376 73958
rect 66400 73956 66456 73958
rect 66480 73956 66536 73958
rect 66560 73956 66616 73958
rect 65660 73466 65716 73468
rect 65740 73466 65796 73468
rect 65820 73466 65876 73468
rect 65900 73466 65956 73468
rect 65660 73414 65706 73466
rect 65706 73414 65716 73466
rect 65740 73414 65770 73466
rect 65770 73414 65782 73466
rect 65782 73414 65796 73466
rect 65820 73414 65834 73466
rect 65834 73414 65846 73466
rect 65846 73414 65876 73466
rect 65900 73414 65910 73466
rect 65910 73414 65956 73466
rect 65660 73412 65716 73414
rect 65740 73412 65796 73414
rect 65820 73412 65876 73414
rect 65900 73412 65956 73414
rect 66320 72922 66376 72924
rect 66400 72922 66456 72924
rect 66480 72922 66536 72924
rect 66560 72922 66616 72924
rect 66320 72870 66366 72922
rect 66366 72870 66376 72922
rect 66400 72870 66430 72922
rect 66430 72870 66442 72922
rect 66442 72870 66456 72922
rect 66480 72870 66494 72922
rect 66494 72870 66506 72922
rect 66506 72870 66536 72922
rect 66560 72870 66570 72922
rect 66570 72870 66616 72922
rect 66320 72868 66376 72870
rect 66400 72868 66456 72870
rect 66480 72868 66536 72870
rect 66560 72868 66616 72870
rect 65660 72378 65716 72380
rect 65740 72378 65796 72380
rect 65820 72378 65876 72380
rect 65900 72378 65956 72380
rect 65660 72326 65706 72378
rect 65706 72326 65716 72378
rect 65740 72326 65770 72378
rect 65770 72326 65782 72378
rect 65782 72326 65796 72378
rect 65820 72326 65834 72378
rect 65834 72326 65846 72378
rect 65846 72326 65876 72378
rect 65900 72326 65910 72378
rect 65910 72326 65956 72378
rect 65660 72324 65716 72326
rect 65740 72324 65796 72326
rect 65820 72324 65876 72326
rect 65900 72324 65956 72326
rect 66320 71834 66376 71836
rect 66400 71834 66456 71836
rect 66480 71834 66536 71836
rect 66560 71834 66616 71836
rect 66320 71782 66366 71834
rect 66366 71782 66376 71834
rect 66400 71782 66430 71834
rect 66430 71782 66442 71834
rect 66442 71782 66456 71834
rect 66480 71782 66494 71834
rect 66494 71782 66506 71834
rect 66506 71782 66536 71834
rect 66560 71782 66570 71834
rect 66570 71782 66616 71834
rect 66320 71780 66376 71782
rect 66400 71780 66456 71782
rect 66480 71780 66536 71782
rect 66560 71780 66616 71782
rect 65660 71290 65716 71292
rect 65740 71290 65796 71292
rect 65820 71290 65876 71292
rect 65900 71290 65956 71292
rect 65660 71238 65706 71290
rect 65706 71238 65716 71290
rect 65740 71238 65770 71290
rect 65770 71238 65782 71290
rect 65782 71238 65796 71290
rect 65820 71238 65834 71290
rect 65834 71238 65846 71290
rect 65846 71238 65876 71290
rect 65900 71238 65910 71290
rect 65910 71238 65956 71290
rect 65660 71236 65716 71238
rect 65740 71236 65796 71238
rect 65820 71236 65876 71238
rect 65900 71236 65956 71238
rect 66320 70746 66376 70748
rect 66400 70746 66456 70748
rect 66480 70746 66536 70748
rect 66560 70746 66616 70748
rect 66320 70694 66366 70746
rect 66366 70694 66376 70746
rect 66400 70694 66430 70746
rect 66430 70694 66442 70746
rect 66442 70694 66456 70746
rect 66480 70694 66494 70746
rect 66494 70694 66506 70746
rect 66506 70694 66536 70746
rect 66560 70694 66570 70746
rect 66570 70694 66616 70746
rect 66320 70692 66376 70694
rect 66400 70692 66456 70694
rect 66480 70692 66536 70694
rect 66560 70692 66616 70694
rect 65660 70202 65716 70204
rect 65740 70202 65796 70204
rect 65820 70202 65876 70204
rect 65900 70202 65956 70204
rect 65660 70150 65706 70202
rect 65706 70150 65716 70202
rect 65740 70150 65770 70202
rect 65770 70150 65782 70202
rect 65782 70150 65796 70202
rect 65820 70150 65834 70202
rect 65834 70150 65846 70202
rect 65846 70150 65876 70202
rect 65900 70150 65910 70202
rect 65910 70150 65956 70202
rect 65660 70148 65716 70150
rect 65740 70148 65796 70150
rect 65820 70148 65876 70150
rect 65900 70148 65956 70150
rect 66320 69658 66376 69660
rect 66400 69658 66456 69660
rect 66480 69658 66536 69660
rect 66560 69658 66616 69660
rect 66320 69606 66366 69658
rect 66366 69606 66376 69658
rect 66400 69606 66430 69658
rect 66430 69606 66442 69658
rect 66442 69606 66456 69658
rect 66480 69606 66494 69658
rect 66494 69606 66506 69658
rect 66506 69606 66536 69658
rect 66560 69606 66570 69658
rect 66570 69606 66616 69658
rect 66320 69604 66376 69606
rect 66400 69604 66456 69606
rect 66480 69604 66536 69606
rect 66560 69604 66616 69606
rect 66442 69300 66444 69320
rect 66444 69300 66496 69320
rect 66496 69300 66498 69320
rect 66442 69264 66498 69300
rect 58714 68740 58770 68776
rect 58714 68720 58716 68740
rect 58716 68720 58768 68740
rect 58768 68720 58770 68740
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 61474 68620 61476 68640
rect 61476 68620 61528 68640
rect 61528 68620 61530 68640
rect 45098 65592 45154 65648
rect 41142 64232 41198 64288
rect 61474 68584 61530 68620
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 66320 68570 66376 68572
rect 66400 68570 66456 68572
rect 66480 68570 66536 68572
rect 66560 68570 66616 68572
rect 66320 68518 66366 68570
rect 66366 68518 66376 68570
rect 66400 68518 66430 68570
rect 66430 68518 66442 68570
rect 66442 68518 66456 68570
rect 66480 68518 66494 68570
rect 66494 68518 66506 68570
rect 66506 68518 66536 68570
rect 66560 68518 66570 68570
rect 66570 68518 66616 68570
rect 66320 68516 66376 68518
rect 66400 68516 66456 68518
rect 66480 68516 66536 68518
rect 66560 68516 66616 68518
rect 66320 67482 66376 67484
rect 66400 67482 66456 67484
rect 66480 67482 66536 67484
rect 66560 67482 66616 67484
rect 66320 67430 66366 67482
rect 66366 67430 66376 67482
rect 66400 67430 66430 67482
rect 66430 67430 66442 67482
rect 66442 67430 66456 67482
rect 66480 67430 66494 67482
rect 66494 67430 66506 67482
rect 66506 67430 66536 67482
rect 66560 67430 66570 67482
rect 66570 67430 66616 67482
rect 66320 67428 66376 67430
rect 66400 67428 66456 67430
rect 66480 67428 66536 67430
rect 66560 67428 66616 67430
rect 66320 66394 66376 66396
rect 66400 66394 66456 66396
rect 66480 66394 66536 66396
rect 66560 66394 66616 66396
rect 66320 66342 66366 66394
rect 66366 66342 66376 66394
rect 66400 66342 66430 66394
rect 66430 66342 66442 66394
rect 66442 66342 66456 66394
rect 66480 66342 66494 66394
rect 66494 66342 66506 66394
rect 66506 66342 66536 66394
rect 66560 66342 66570 66394
rect 66570 66342 66616 66394
rect 66320 66340 66376 66342
rect 66400 66340 66456 66342
rect 66480 66340 66536 66342
rect 66560 66340 66616 66342
rect 72698 69808 72754 69864
rect 68650 66172 68652 66192
rect 68652 66172 68704 66192
rect 68704 66172 68706 66192
rect 68650 66136 68706 66172
rect 39946 64096 40002 64152
rect 46478 64096 46534 64152
rect 66074 64096 66130 64152
rect 84842 75928 84898 75984
rect 79322 69844 79324 69864
rect 79324 69844 79376 69864
rect 79376 69844 79378 69864
rect 79322 69808 79378 69844
rect 72422 63960 72478 64016
rect 88982 72528 89038 72584
rect 91466 77696 91522 77752
rect 91558 77424 91614 77480
rect 92202 77560 92258 77616
rect 88246 65900 88248 65920
rect 88248 65900 88300 65920
rect 88300 65900 88302 65920
rect 88246 65864 88302 65900
rect 96380 77818 96436 77820
rect 96460 77818 96516 77820
rect 96540 77818 96596 77820
rect 96620 77818 96676 77820
rect 96380 77766 96426 77818
rect 96426 77766 96436 77818
rect 96460 77766 96490 77818
rect 96490 77766 96502 77818
rect 96502 77766 96516 77818
rect 96540 77766 96554 77818
rect 96554 77766 96566 77818
rect 96566 77766 96596 77818
rect 96620 77766 96630 77818
rect 96630 77766 96676 77818
rect 96380 77764 96436 77766
rect 96460 77764 96516 77766
rect 96540 77764 96596 77766
rect 96620 77764 96676 77766
rect 96380 76730 96436 76732
rect 96460 76730 96516 76732
rect 96540 76730 96596 76732
rect 96620 76730 96676 76732
rect 96380 76678 96426 76730
rect 96426 76678 96436 76730
rect 96460 76678 96490 76730
rect 96490 76678 96502 76730
rect 96502 76678 96516 76730
rect 96540 76678 96554 76730
rect 96554 76678 96566 76730
rect 96566 76678 96596 76730
rect 96620 76678 96630 76730
rect 96630 76678 96676 76730
rect 96380 76676 96436 76678
rect 96460 76676 96516 76678
rect 96540 76676 96596 76678
rect 96620 76676 96676 76678
rect 96380 75642 96436 75644
rect 96460 75642 96516 75644
rect 96540 75642 96596 75644
rect 96620 75642 96676 75644
rect 96380 75590 96426 75642
rect 96426 75590 96436 75642
rect 96460 75590 96490 75642
rect 96490 75590 96502 75642
rect 96502 75590 96516 75642
rect 96540 75590 96554 75642
rect 96554 75590 96566 75642
rect 96566 75590 96596 75642
rect 96620 75590 96630 75642
rect 96630 75590 96676 75642
rect 96380 75588 96436 75590
rect 96460 75588 96516 75590
rect 96540 75588 96596 75590
rect 96620 75588 96676 75590
rect 97040 77274 97096 77276
rect 97120 77274 97176 77276
rect 97200 77274 97256 77276
rect 97280 77274 97336 77276
rect 97040 77222 97086 77274
rect 97086 77222 97096 77274
rect 97120 77222 97150 77274
rect 97150 77222 97162 77274
rect 97162 77222 97176 77274
rect 97200 77222 97214 77274
rect 97214 77222 97226 77274
rect 97226 77222 97256 77274
rect 97280 77222 97290 77274
rect 97290 77222 97336 77274
rect 97040 77220 97096 77222
rect 97120 77220 97176 77222
rect 97200 77220 97256 77222
rect 97280 77220 97336 77222
rect 105928 136570 105984 136572
rect 106008 136570 106064 136572
rect 106088 136570 106144 136572
rect 106168 136570 106224 136572
rect 105928 136518 105974 136570
rect 105974 136518 105984 136570
rect 106008 136518 106038 136570
rect 106038 136518 106050 136570
rect 106050 136518 106064 136570
rect 106088 136518 106102 136570
rect 106102 136518 106114 136570
rect 106114 136518 106144 136570
rect 106168 136518 106178 136570
rect 106178 136518 106224 136570
rect 105928 136516 105984 136518
rect 106008 136516 106064 136518
rect 106088 136516 106144 136518
rect 106168 136516 106224 136518
rect 97040 76186 97096 76188
rect 97120 76186 97176 76188
rect 97200 76186 97256 76188
rect 97280 76186 97336 76188
rect 97040 76134 97086 76186
rect 97086 76134 97096 76186
rect 97120 76134 97150 76186
rect 97150 76134 97162 76186
rect 97162 76134 97176 76186
rect 97200 76134 97214 76186
rect 97214 76134 97226 76186
rect 97226 76134 97256 76186
rect 97280 76134 97290 76186
rect 97290 76134 97336 76186
rect 97040 76132 97096 76134
rect 97120 76132 97176 76134
rect 97200 76132 97256 76134
rect 97280 76132 97336 76134
rect 96380 74554 96436 74556
rect 96460 74554 96516 74556
rect 96540 74554 96596 74556
rect 96620 74554 96676 74556
rect 96380 74502 96426 74554
rect 96426 74502 96436 74554
rect 96460 74502 96490 74554
rect 96490 74502 96502 74554
rect 96502 74502 96516 74554
rect 96540 74502 96554 74554
rect 96554 74502 96566 74554
rect 96566 74502 96596 74554
rect 96620 74502 96630 74554
rect 96630 74502 96676 74554
rect 96380 74500 96436 74502
rect 96460 74500 96516 74502
rect 96540 74500 96596 74502
rect 96620 74500 96676 74502
rect 97040 75098 97096 75100
rect 97120 75098 97176 75100
rect 97200 75098 97256 75100
rect 97280 75098 97336 75100
rect 97040 75046 97086 75098
rect 97086 75046 97096 75098
rect 97120 75046 97150 75098
rect 97150 75046 97162 75098
rect 97162 75046 97176 75098
rect 97200 75046 97214 75098
rect 97214 75046 97226 75098
rect 97226 75046 97256 75098
rect 97280 75046 97290 75098
rect 97290 75046 97336 75098
rect 97040 75044 97096 75046
rect 97120 75044 97176 75046
rect 97200 75044 97256 75046
rect 97280 75044 97336 75046
rect 96380 73466 96436 73468
rect 96460 73466 96516 73468
rect 96540 73466 96596 73468
rect 96620 73466 96676 73468
rect 96380 73414 96426 73466
rect 96426 73414 96436 73466
rect 96460 73414 96490 73466
rect 96490 73414 96502 73466
rect 96502 73414 96516 73466
rect 96540 73414 96554 73466
rect 96554 73414 96566 73466
rect 96566 73414 96596 73466
rect 96620 73414 96630 73466
rect 96630 73414 96676 73466
rect 96380 73412 96436 73414
rect 96460 73412 96516 73414
rect 96540 73412 96596 73414
rect 96620 73412 96676 73414
rect 97040 74010 97096 74012
rect 97120 74010 97176 74012
rect 97200 74010 97256 74012
rect 97280 74010 97336 74012
rect 97040 73958 97086 74010
rect 97086 73958 97096 74010
rect 97120 73958 97150 74010
rect 97150 73958 97162 74010
rect 97162 73958 97176 74010
rect 97200 73958 97214 74010
rect 97214 73958 97226 74010
rect 97226 73958 97256 74010
rect 97280 73958 97290 74010
rect 97290 73958 97336 74010
rect 97040 73956 97096 73958
rect 97120 73956 97176 73958
rect 97200 73956 97256 73958
rect 97280 73956 97336 73958
rect 97040 72922 97096 72924
rect 97120 72922 97176 72924
rect 97200 72922 97256 72924
rect 97280 72922 97336 72924
rect 97040 72870 97086 72922
rect 97086 72870 97096 72922
rect 97120 72870 97150 72922
rect 97150 72870 97162 72922
rect 97162 72870 97176 72922
rect 97200 72870 97214 72922
rect 97214 72870 97226 72922
rect 97226 72870 97256 72922
rect 97280 72870 97290 72922
rect 97290 72870 97336 72922
rect 97040 72868 97096 72870
rect 97120 72868 97176 72870
rect 97200 72868 97256 72870
rect 97280 72868 97336 72870
rect 96380 72378 96436 72380
rect 96460 72378 96516 72380
rect 96540 72378 96596 72380
rect 96620 72378 96676 72380
rect 96380 72326 96426 72378
rect 96426 72326 96436 72378
rect 96460 72326 96490 72378
rect 96490 72326 96502 72378
rect 96502 72326 96516 72378
rect 96540 72326 96554 72378
rect 96554 72326 96566 72378
rect 96566 72326 96596 72378
rect 96620 72326 96630 72378
rect 96630 72326 96676 72378
rect 96380 72324 96436 72326
rect 96460 72324 96516 72326
rect 96540 72324 96596 72326
rect 96620 72324 96676 72326
rect 96380 71290 96436 71292
rect 96460 71290 96516 71292
rect 96540 71290 96596 71292
rect 96620 71290 96676 71292
rect 96380 71238 96426 71290
rect 96426 71238 96436 71290
rect 96460 71238 96490 71290
rect 96490 71238 96502 71290
rect 96502 71238 96516 71290
rect 96540 71238 96554 71290
rect 96554 71238 96566 71290
rect 96566 71238 96596 71290
rect 96620 71238 96630 71290
rect 96630 71238 96676 71290
rect 96380 71236 96436 71238
rect 96460 71236 96516 71238
rect 96540 71236 96596 71238
rect 96620 71236 96676 71238
rect 97040 71834 97096 71836
rect 97120 71834 97176 71836
rect 97200 71834 97256 71836
rect 97280 71834 97336 71836
rect 97040 71782 97086 71834
rect 97086 71782 97096 71834
rect 97120 71782 97150 71834
rect 97150 71782 97162 71834
rect 97162 71782 97176 71834
rect 97200 71782 97214 71834
rect 97214 71782 97226 71834
rect 97226 71782 97256 71834
rect 97280 71782 97290 71834
rect 97290 71782 97336 71834
rect 97040 71780 97096 71782
rect 97120 71780 97176 71782
rect 97200 71780 97256 71782
rect 97280 71780 97336 71782
rect 98826 74160 98882 74216
rect 98550 73364 98606 73400
rect 98550 73344 98552 73364
rect 98552 73344 98604 73364
rect 98604 73344 98606 73364
rect 99102 73208 99158 73264
rect 102506 95032 102562 95088
rect 102414 93332 102470 93388
rect 102230 76472 102286 76528
rect 99470 74432 99526 74488
rect 99470 73344 99526 73400
rect 97040 70746 97096 70748
rect 97120 70746 97176 70748
rect 97200 70746 97256 70748
rect 97280 70746 97336 70748
rect 97040 70694 97086 70746
rect 97086 70694 97096 70746
rect 97120 70694 97150 70746
rect 97150 70694 97162 70746
rect 97162 70694 97176 70746
rect 97200 70694 97214 70746
rect 97214 70694 97226 70746
rect 97226 70694 97256 70746
rect 97280 70694 97290 70746
rect 97290 70694 97336 70746
rect 97040 70692 97096 70694
rect 97120 70692 97176 70694
rect 97200 70692 97256 70694
rect 97280 70692 97336 70694
rect 96380 70202 96436 70204
rect 96460 70202 96516 70204
rect 96540 70202 96596 70204
rect 96620 70202 96676 70204
rect 96380 70150 96426 70202
rect 96426 70150 96436 70202
rect 96460 70150 96490 70202
rect 96490 70150 96502 70202
rect 96502 70150 96516 70202
rect 96540 70150 96554 70202
rect 96554 70150 96566 70202
rect 96566 70150 96596 70202
rect 96620 70150 96630 70202
rect 96630 70150 96676 70202
rect 96380 70148 96436 70150
rect 96460 70148 96516 70150
rect 96540 70148 96596 70150
rect 96620 70148 96676 70150
rect 97722 71068 97724 71088
rect 97724 71068 97776 71088
rect 97776 71068 97778 71088
rect 97722 71032 97778 71068
rect 99654 73208 99710 73264
rect 97538 69944 97594 70000
rect 98182 71032 98238 71088
rect 103610 77016 103666 77072
rect 103886 129804 103942 129840
rect 103886 129784 103888 129804
rect 103888 129784 103940 129804
rect 103940 129784 103942 129804
rect 103886 92248 103942 92304
rect 103794 76880 103850 76936
rect 103702 76336 103758 76392
rect 103518 75928 103574 75984
rect 106664 136026 106720 136028
rect 106744 136026 106800 136028
rect 106824 136026 106880 136028
rect 106904 136026 106960 136028
rect 106664 135974 106710 136026
rect 106710 135974 106720 136026
rect 106744 135974 106774 136026
rect 106774 135974 106786 136026
rect 106786 135974 106800 136026
rect 106824 135974 106838 136026
rect 106838 135974 106850 136026
rect 106850 135974 106880 136026
rect 106904 135974 106914 136026
rect 106914 135974 106960 136026
rect 106664 135972 106720 135974
rect 106744 135972 106800 135974
rect 106824 135972 106880 135974
rect 106904 135972 106960 135974
rect 105928 135482 105984 135484
rect 106008 135482 106064 135484
rect 106088 135482 106144 135484
rect 106168 135482 106224 135484
rect 105928 135430 105974 135482
rect 105974 135430 105984 135482
rect 106008 135430 106038 135482
rect 106038 135430 106050 135482
rect 106050 135430 106064 135482
rect 106088 135430 106102 135482
rect 106102 135430 106114 135482
rect 106114 135430 106144 135482
rect 106168 135430 106178 135482
rect 106178 135430 106224 135482
rect 105928 135428 105984 135430
rect 106008 135428 106064 135430
rect 106088 135428 106144 135430
rect 106168 135428 106224 135430
rect 106664 134938 106720 134940
rect 106744 134938 106800 134940
rect 106824 134938 106880 134940
rect 106904 134938 106960 134940
rect 106664 134886 106710 134938
rect 106710 134886 106720 134938
rect 106744 134886 106774 134938
rect 106774 134886 106786 134938
rect 106786 134886 106800 134938
rect 106824 134886 106838 134938
rect 106838 134886 106850 134938
rect 106850 134886 106880 134938
rect 106904 134886 106914 134938
rect 106914 134886 106960 134938
rect 106664 134884 106720 134886
rect 106744 134884 106800 134886
rect 106824 134884 106880 134886
rect 106904 134884 106960 134886
rect 105928 134394 105984 134396
rect 106008 134394 106064 134396
rect 106088 134394 106144 134396
rect 106168 134394 106224 134396
rect 105928 134342 105974 134394
rect 105974 134342 105984 134394
rect 106008 134342 106038 134394
rect 106038 134342 106050 134394
rect 106050 134342 106064 134394
rect 106088 134342 106102 134394
rect 106102 134342 106114 134394
rect 106114 134342 106144 134394
rect 106168 134342 106178 134394
rect 106178 134342 106224 134394
rect 105928 134340 105984 134342
rect 106008 134340 106064 134342
rect 106088 134340 106144 134342
rect 106168 134340 106224 134342
rect 106664 133850 106720 133852
rect 106744 133850 106800 133852
rect 106824 133850 106880 133852
rect 106904 133850 106960 133852
rect 106664 133798 106710 133850
rect 106710 133798 106720 133850
rect 106744 133798 106774 133850
rect 106774 133798 106786 133850
rect 106786 133798 106800 133850
rect 106824 133798 106838 133850
rect 106838 133798 106850 133850
rect 106850 133798 106880 133850
rect 106904 133798 106914 133850
rect 106914 133798 106960 133850
rect 106664 133796 106720 133798
rect 106744 133796 106800 133798
rect 106824 133796 106880 133798
rect 106904 133796 106960 133798
rect 105928 133306 105984 133308
rect 106008 133306 106064 133308
rect 106088 133306 106144 133308
rect 106168 133306 106224 133308
rect 105928 133254 105974 133306
rect 105974 133254 105984 133306
rect 106008 133254 106038 133306
rect 106038 133254 106050 133306
rect 106050 133254 106064 133306
rect 106088 133254 106102 133306
rect 106102 133254 106114 133306
rect 106114 133254 106144 133306
rect 106168 133254 106178 133306
rect 106178 133254 106224 133306
rect 105928 133252 105984 133254
rect 106008 133252 106064 133254
rect 106088 133252 106144 133254
rect 106168 133252 106224 133254
rect 106664 132762 106720 132764
rect 106744 132762 106800 132764
rect 106824 132762 106880 132764
rect 106904 132762 106960 132764
rect 106664 132710 106710 132762
rect 106710 132710 106720 132762
rect 106744 132710 106774 132762
rect 106774 132710 106786 132762
rect 106786 132710 106800 132762
rect 106824 132710 106838 132762
rect 106838 132710 106850 132762
rect 106850 132710 106880 132762
rect 106904 132710 106914 132762
rect 106914 132710 106960 132762
rect 106664 132708 106720 132710
rect 106744 132708 106800 132710
rect 106824 132708 106880 132710
rect 106904 132708 106960 132710
rect 105928 132218 105984 132220
rect 106008 132218 106064 132220
rect 106088 132218 106144 132220
rect 106168 132218 106224 132220
rect 105928 132166 105974 132218
rect 105974 132166 105984 132218
rect 106008 132166 106038 132218
rect 106038 132166 106050 132218
rect 106050 132166 106064 132218
rect 106088 132166 106102 132218
rect 106102 132166 106114 132218
rect 106114 132166 106144 132218
rect 106168 132166 106178 132218
rect 106178 132166 106224 132218
rect 105928 132164 105984 132166
rect 106008 132164 106064 132166
rect 106088 132164 106144 132166
rect 106168 132164 106224 132166
rect 106664 131674 106720 131676
rect 106744 131674 106800 131676
rect 106824 131674 106880 131676
rect 106904 131674 106960 131676
rect 106664 131622 106710 131674
rect 106710 131622 106720 131674
rect 106744 131622 106774 131674
rect 106774 131622 106786 131674
rect 106786 131622 106800 131674
rect 106824 131622 106838 131674
rect 106838 131622 106850 131674
rect 106850 131622 106880 131674
rect 106904 131622 106914 131674
rect 106914 131622 106960 131674
rect 106664 131620 106720 131622
rect 106744 131620 106800 131622
rect 106824 131620 106880 131622
rect 106904 131620 106960 131622
rect 105928 131130 105984 131132
rect 106008 131130 106064 131132
rect 106088 131130 106144 131132
rect 106168 131130 106224 131132
rect 105928 131078 105974 131130
rect 105974 131078 105984 131130
rect 106008 131078 106038 131130
rect 106038 131078 106050 131130
rect 106050 131078 106064 131130
rect 106088 131078 106102 131130
rect 106102 131078 106114 131130
rect 106114 131078 106144 131130
rect 106168 131078 106178 131130
rect 106178 131078 106224 131130
rect 105928 131076 105984 131078
rect 106008 131076 106064 131078
rect 106088 131076 106144 131078
rect 106168 131076 106224 131078
rect 106664 130586 106720 130588
rect 106744 130586 106800 130588
rect 106824 130586 106880 130588
rect 106904 130586 106960 130588
rect 106664 130534 106710 130586
rect 106710 130534 106720 130586
rect 106744 130534 106774 130586
rect 106774 130534 106786 130586
rect 106786 130534 106800 130586
rect 106824 130534 106838 130586
rect 106838 130534 106850 130586
rect 106850 130534 106880 130586
rect 106904 130534 106914 130586
rect 106914 130534 106960 130586
rect 106664 130532 106720 130534
rect 106744 130532 106800 130534
rect 106824 130532 106880 130534
rect 106904 130532 106960 130534
rect 105928 130042 105984 130044
rect 106008 130042 106064 130044
rect 106088 130042 106144 130044
rect 106168 130042 106224 130044
rect 105928 129990 105974 130042
rect 105974 129990 105984 130042
rect 106008 129990 106038 130042
rect 106038 129990 106050 130042
rect 106050 129990 106064 130042
rect 106088 129990 106102 130042
rect 106102 129990 106114 130042
rect 106114 129990 106144 130042
rect 106168 129990 106178 130042
rect 106178 129990 106224 130042
rect 105928 129988 105984 129990
rect 106008 129988 106064 129990
rect 106088 129988 106144 129990
rect 106168 129988 106224 129990
rect 106664 129498 106720 129500
rect 106744 129498 106800 129500
rect 106824 129498 106880 129500
rect 106904 129498 106960 129500
rect 106664 129446 106710 129498
rect 106710 129446 106720 129498
rect 106744 129446 106774 129498
rect 106774 129446 106786 129498
rect 106786 129446 106800 129498
rect 106824 129446 106838 129498
rect 106838 129446 106850 129498
rect 106850 129446 106880 129498
rect 106904 129446 106914 129498
rect 106914 129446 106960 129498
rect 106664 129444 106720 129446
rect 106744 129444 106800 129446
rect 106824 129444 106880 129446
rect 106904 129444 106960 129446
rect 105928 128954 105984 128956
rect 106008 128954 106064 128956
rect 106088 128954 106144 128956
rect 106168 128954 106224 128956
rect 105928 128902 105974 128954
rect 105974 128902 105984 128954
rect 106008 128902 106038 128954
rect 106038 128902 106050 128954
rect 106050 128902 106064 128954
rect 106088 128902 106102 128954
rect 106102 128902 106114 128954
rect 106114 128902 106144 128954
rect 106168 128902 106178 128954
rect 106178 128902 106224 128954
rect 105928 128900 105984 128902
rect 106008 128900 106064 128902
rect 106088 128900 106144 128902
rect 106168 128900 106224 128902
rect 106664 128410 106720 128412
rect 106744 128410 106800 128412
rect 106824 128410 106880 128412
rect 106904 128410 106960 128412
rect 106664 128358 106710 128410
rect 106710 128358 106720 128410
rect 106744 128358 106774 128410
rect 106774 128358 106786 128410
rect 106786 128358 106800 128410
rect 106824 128358 106838 128410
rect 106838 128358 106850 128410
rect 106850 128358 106880 128410
rect 106904 128358 106914 128410
rect 106914 128358 106960 128410
rect 106664 128356 106720 128358
rect 106744 128356 106800 128358
rect 106824 128356 106880 128358
rect 106904 128356 106960 128358
rect 105928 127866 105984 127868
rect 106008 127866 106064 127868
rect 106088 127866 106144 127868
rect 106168 127866 106224 127868
rect 105928 127814 105974 127866
rect 105974 127814 105984 127866
rect 106008 127814 106038 127866
rect 106038 127814 106050 127866
rect 106050 127814 106064 127866
rect 106088 127814 106102 127866
rect 106102 127814 106114 127866
rect 106114 127814 106144 127866
rect 106168 127814 106178 127866
rect 106178 127814 106224 127866
rect 105928 127812 105984 127814
rect 106008 127812 106064 127814
rect 106088 127812 106144 127814
rect 106168 127812 106224 127814
rect 106664 127322 106720 127324
rect 106744 127322 106800 127324
rect 106824 127322 106880 127324
rect 106904 127322 106960 127324
rect 106664 127270 106710 127322
rect 106710 127270 106720 127322
rect 106744 127270 106774 127322
rect 106774 127270 106786 127322
rect 106786 127270 106800 127322
rect 106824 127270 106838 127322
rect 106838 127270 106850 127322
rect 106850 127270 106880 127322
rect 106904 127270 106914 127322
rect 106914 127270 106960 127322
rect 106664 127268 106720 127270
rect 106744 127268 106800 127270
rect 106824 127268 106880 127270
rect 106904 127268 106960 127270
rect 105928 126778 105984 126780
rect 106008 126778 106064 126780
rect 106088 126778 106144 126780
rect 106168 126778 106224 126780
rect 105928 126726 105974 126778
rect 105974 126726 105984 126778
rect 106008 126726 106038 126778
rect 106038 126726 106050 126778
rect 106050 126726 106064 126778
rect 106088 126726 106102 126778
rect 106102 126726 106114 126778
rect 106114 126726 106144 126778
rect 106168 126726 106178 126778
rect 106178 126726 106224 126778
rect 105928 126724 105984 126726
rect 106008 126724 106064 126726
rect 106088 126724 106144 126726
rect 106168 126724 106224 126726
rect 106664 126234 106720 126236
rect 106744 126234 106800 126236
rect 106824 126234 106880 126236
rect 106904 126234 106960 126236
rect 106664 126182 106710 126234
rect 106710 126182 106720 126234
rect 106744 126182 106774 126234
rect 106774 126182 106786 126234
rect 106786 126182 106800 126234
rect 106824 126182 106838 126234
rect 106838 126182 106850 126234
rect 106850 126182 106880 126234
rect 106904 126182 106914 126234
rect 106914 126182 106960 126234
rect 106664 126180 106720 126182
rect 106744 126180 106800 126182
rect 106824 126180 106880 126182
rect 106904 126180 106960 126182
rect 105928 125690 105984 125692
rect 106008 125690 106064 125692
rect 106088 125690 106144 125692
rect 106168 125690 106224 125692
rect 105928 125638 105974 125690
rect 105974 125638 105984 125690
rect 106008 125638 106038 125690
rect 106038 125638 106050 125690
rect 106050 125638 106064 125690
rect 106088 125638 106102 125690
rect 106102 125638 106114 125690
rect 106114 125638 106144 125690
rect 106168 125638 106178 125690
rect 106178 125638 106224 125690
rect 105928 125636 105984 125638
rect 106008 125636 106064 125638
rect 106088 125636 106144 125638
rect 106168 125636 106224 125638
rect 106664 125146 106720 125148
rect 106744 125146 106800 125148
rect 106824 125146 106880 125148
rect 106904 125146 106960 125148
rect 106664 125094 106710 125146
rect 106710 125094 106720 125146
rect 106744 125094 106774 125146
rect 106774 125094 106786 125146
rect 106786 125094 106800 125146
rect 106824 125094 106838 125146
rect 106838 125094 106850 125146
rect 106850 125094 106880 125146
rect 106904 125094 106914 125146
rect 106914 125094 106960 125146
rect 106664 125092 106720 125094
rect 106744 125092 106800 125094
rect 106824 125092 106880 125094
rect 106904 125092 106960 125094
rect 105928 124602 105984 124604
rect 106008 124602 106064 124604
rect 106088 124602 106144 124604
rect 106168 124602 106224 124604
rect 105928 124550 105974 124602
rect 105974 124550 105984 124602
rect 106008 124550 106038 124602
rect 106038 124550 106050 124602
rect 106050 124550 106064 124602
rect 106088 124550 106102 124602
rect 106102 124550 106114 124602
rect 106114 124550 106144 124602
rect 106168 124550 106178 124602
rect 106178 124550 106224 124602
rect 105928 124548 105984 124550
rect 106008 124548 106064 124550
rect 106088 124548 106144 124550
rect 106168 124548 106224 124550
rect 106664 124058 106720 124060
rect 106744 124058 106800 124060
rect 106824 124058 106880 124060
rect 106904 124058 106960 124060
rect 106664 124006 106710 124058
rect 106710 124006 106720 124058
rect 106744 124006 106774 124058
rect 106774 124006 106786 124058
rect 106786 124006 106800 124058
rect 106824 124006 106838 124058
rect 106838 124006 106850 124058
rect 106850 124006 106880 124058
rect 106904 124006 106914 124058
rect 106914 124006 106960 124058
rect 106664 124004 106720 124006
rect 106744 124004 106800 124006
rect 106824 124004 106880 124006
rect 106904 124004 106960 124006
rect 105928 123514 105984 123516
rect 106008 123514 106064 123516
rect 106088 123514 106144 123516
rect 106168 123514 106224 123516
rect 105928 123462 105974 123514
rect 105974 123462 105984 123514
rect 106008 123462 106038 123514
rect 106038 123462 106050 123514
rect 106050 123462 106064 123514
rect 106088 123462 106102 123514
rect 106102 123462 106114 123514
rect 106114 123462 106144 123514
rect 106168 123462 106178 123514
rect 106178 123462 106224 123514
rect 105928 123460 105984 123462
rect 106008 123460 106064 123462
rect 106088 123460 106144 123462
rect 106168 123460 106224 123462
rect 106664 122970 106720 122972
rect 106744 122970 106800 122972
rect 106824 122970 106880 122972
rect 106904 122970 106960 122972
rect 106664 122918 106710 122970
rect 106710 122918 106720 122970
rect 106744 122918 106774 122970
rect 106774 122918 106786 122970
rect 106786 122918 106800 122970
rect 106824 122918 106838 122970
rect 106838 122918 106850 122970
rect 106850 122918 106880 122970
rect 106904 122918 106914 122970
rect 106914 122918 106960 122970
rect 106664 122916 106720 122918
rect 106744 122916 106800 122918
rect 106824 122916 106880 122918
rect 106904 122916 106960 122918
rect 105928 122426 105984 122428
rect 106008 122426 106064 122428
rect 106088 122426 106144 122428
rect 106168 122426 106224 122428
rect 105928 122374 105974 122426
rect 105974 122374 105984 122426
rect 106008 122374 106038 122426
rect 106038 122374 106050 122426
rect 106050 122374 106064 122426
rect 106088 122374 106102 122426
rect 106102 122374 106114 122426
rect 106114 122374 106144 122426
rect 106168 122374 106178 122426
rect 106178 122374 106224 122426
rect 105928 122372 105984 122374
rect 106008 122372 106064 122374
rect 106088 122372 106144 122374
rect 106168 122372 106224 122374
rect 106664 121882 106720 121884
rect 106744 121882 106800 121884
rect 106824 121882 106880 121884
rect 106904 121882 106960 121884
rect 106664 121830 106710 121882
rect 106710 121830 106720 121882
rect 106744 121830 106774 121882
rect 106774 121830 106786 121882
rect 106786 121830 106800 121882
rect 106824 121830 106838 121882
rect 106838 121830 106850 121882
rect 106850 121830 106880 121882
rect 106904 121830 106914 121882
rect 106914 121830 106960 121882
rect 106664 121828 106720 121830
rect 106744 121828 106800 121830
rect 106824 121828 106880 121830
rect 106904 121828 106960 121830
rect 105928 121338 105984 121340
rect 106008 121338 106064 121340
rect 106088 121338 106144 121340
rect 106168 121338 106224 121340
rect 105928 121286 105974 121338
rect 105974 121286 105984 121338
rect 106008 121286 106038 121338
rect 106038 121286 106050 121338
rect 106050 121286 106064 121338
rect 106088 121286 106102 121338
rect 106102 121286 106114 121338
rect 106114 121286 106144 121338
rect 106168 121286 106178 121338
rect 106178 121286 106224 121338
rect 105928 121284 105984 121286
rect 106008 121284 106064 121286
rect 106088 121284 106144 121286
rect 106168 121284 106224 121286
rect 106664 120794 106720 120796
rect 106744 120794 106800 120796
rect 106824 120794 106880 120796
rect 106904 120794 106960 120796
rect 106664 120742 106710 120794
rect 106710 120742 106720 120794
rect 106744 120742 106774 120794
rect 106774 120742 106786 120794
rect 106786 120742 106800 120794
rect 106824 120742 106838 120794
rect 106838 120742 106850 120794
rect 106850 120742 106880 120794
rect 106904 120742 106914 120794
rect 106914 120742 106960 120794
rect 106664 120740 106720 120742
rect 106744 120740 106800 120742
rect 106824 120740 106880 120742
rect 106904 120740 106960 120742
rect 105928 120250 105984 120252
rect 106008 120250 106064 120252
rect 106088 120250 106144 120252
rect 106168 120250 106224 120252
rect 105928 120198 105974 120250
rect 105974 120198 105984 120250
rect 106008 120198 106038 120250
rect 106038 120198 106050 120250
rect 106050 120198 106064 120250
rect 106088 120198 106102 120250
rect 106102 120198 106114 120250
rect 106114 120198 106144 120250
rect 106168 120198 106178 120250
rect 106178 120198 106224 120250
rect 105928 120196 105984 120198
rect 106008 120196 106064 120198
rect 106088 120196 106144 120198
rect 106168 120196 106224 120198
rect 106664 119706 106720 119708
rect 106744 119706 106800 119708
rect 106824 119706 106880 119708
rect 106904 119706 106960 119708
rect 106664 119654 106710 119706
rect 106710 119654 106720 119706
rect 106744 119654 106774 119706
rect 106774 119654 106786 119706
rect 106786 119654 106800 119706
rect 106824 119654 106838 119706
rect 106838 119654 106850 119706
rect 106850 119654 106880 119706
rect 106904 119654 106914 119706
rect 106914 119654 106960 119706
rect 106664 119652 106720 119654
rect 106744 119652 106800 119654
rect 106824 119652 106880 119654
rect 106904 119652 106960 119654
rect 105928 119162 105984 119164
rect 106008 119162 106064 119164
rect 106088 119162 106144 119164
rect 106168 119162 106224 119164
rect 105928 119110 105974 119162
rect 105974 119110 105984 119162
rect 106008 119110 106038 119162
rect 106038 119110 106050 119162
rect 106050 119110 106064 119162
rect 106088 119110 106102 119162
rect 106102 119110 106114 119162
rect 106114 119110 106144 119162
rect 106168 119110 106178 119162
rect 106178 119110 106224 119162
rect 105928 119108 105984 119110
rect 106008 119108 106064 119110
rect 106088 119108 106144 119110
rect 106168 119108 106224 119110
rect 106664 118618 106720 118620
rect 106744 118618 106800 118620
rect 106824 118618 106880 118620
rect 106904 118618 106960 118620
rect 106664 118566 106710 118618
rect 106710 118566 106720 118618
rect 106744 118566 106774 118618
rect 106774 118566 106786 118618
rect 106786 118566 106800 118618
rect 106824 118566 106838 118618
rect 106838 118566 106850 118618
rect 106850 118566 106880 118618
rect 106904 118566 106914 118618
rect 106914 118566 106960 118618
rect 106664 118564 106720 118566
rect 106744 118564 106800 118566
rect 106824 118564 106880 118566
rect 106904 118564 106960 118566
rect 105928 118074 105984 118076
rect 106008 118074 106064 118076
rect 106088 118074 106144 118076
rect 106168 118074 106224 118076
rect 105928 118022 105974 118074
rect 105974 118022 105984 118074
rect 106008 118022 106038 118074
rect 106038 118022 106050 118074
rect 106050 118022 106064 118074
rect 106088 118022 106102 118074
rect 106102 118022 106114 118074
rect 106114 118022 106144 118074
rect 106168 118022 106178 118074
rect 106178 118022 106224 118074
rect 105928 118020 105984 118022
rect 106008 118020 106064 118022
rect 106088 118020 106144 118022
rect 106168 118020 106224 118022
rect 106664 117530 106720 117532
rect 106744 117530 106800 117532
rect 106824 117530 106880 117532
rect 106904 117530 106960 117532
rect 106664 117478 106710 117530
rect 106710 117478 106720 117530
rect 106744 117478 106774 117530
rect 106774 117478 106786 117530
rect 106786 117478 106800 117530
rect 106824 117478 106838 117530
rect 106838 117478 106850 117530
rect 106850 117478 106880 117530
rect 106904 117478 106914 117530
rect 106914 117478 106960 117530
rect 106664 117476 106720 117478
rect 106744 117476 106800 117478
rect 106824 117476 106880 117478
rect 106904 117476 106960 117478
rect 105928 116986 105984 116988
rect 106008 116986 106064 116988
rect 106088 116986 106144 116988
rect 106168 116986 106224 116988
rect 105928 116934 105974 116986
rect 105974 116934 105984 116986
rect 106008 116934 106038 116986
rect 106038 116934 106050 116986
rect 106050 116934 106064 116986
rect 106088 116934 106102 116986
rect 106102 116934 106114 116986
rect 106114 116934 106144 116986
rect 106168 116934 106178 116986
rect 106178 116934 106224 116986
rect 105928 116932 105984 116934
rect 106008 116932 106064 116934
rect 106088 116932 106144 116934
rect 106168 116932 106224 116934
rect 106664 116442 106720 116444
rect 106744 116442 106800 116444
rect 106824 116442 106880 116444
rect 106904 116442 106960 116444
rect 106664 116390 106710 116442
rect 106710 116390 106720 116442
rect 106744 116390 106774 116442
rect 106774 116390 106786 116442
rect 106786 116390 106800 116442
rect 106824 116390 106838 116442
rect 106838 116390 106850 116442
rect 106850 116390 106880 116442
rect 106904 116390 106914 116442
rect 106914 116390 106960 116442
rect 106664 116388 106720 116390
rect 106744 116388 106800 116390
rect 106824 116388 106880 116390
rect 106904 116388 106960 116390
rect 105928 115898 105984 115900
rect 106008 115898 106064 115900
rect 106088 115898 106144 115900
rect 106168 115898 106224 115900
rect 105928 115846 105974 115898
rect 105974 115846 105984 115898
rect 106008 115846 106038 115898
rect 106038 115846 106050 115898
rect 106050 115846 106064 115898
rect 106088 115846 106102 115898
rect 106102 115846 106114 115898
rect 106114 115846 106144 115898
rect 106168 115846 106178 115898
rect 106178 115846 106224 115898
rect 105928 115844 105984 115846
rect 106008 115844 106064 115846
rect 106088 115844 106144 115846
rect 106168 115844 106224 115846
rect 106664 115354 106720 115356
rect 106744 115354 106800 115356
rect 106824 115354 106880 115356
rect 106904 115354 106960 115356
rect 106664 115302 106710 115354
rect 106710 115302 106720 115354
rect 106744 115302 106774 115354
rect 106774 115302 106786 115354
rect 106786 115302 106800 115354
rect 106824 115302 106838 115354
rect 106838 115302 106850 115354
rect 106850 115302 106880 115354
rect 106904 115302 106914 115354
rect 106914 115302 106960 115354
rect 106664 115300 106720 115302
rect 106744 115300 106800 115302
rect 106824 115300 106880 115302
rect 106904 115300 106960 115302
rect 105928 114810 105984 114812
rect 106008 114810 106064 114812
rect 106088 114810 106144 114812
rect 106168 114810 106224 114812
rect 105928 114758 105974 114810
rect 105974 114758 105984 114810
rect 106008 114758 106038 114810
rect 106038 114758 106050 114810
rect 106050 114758 106064 114810
rect 106088 114758 106102 114810
rect 106102 114758 106114 114810
rect 106114 114758 106144 114810
rect 106168 114758 106178 114810
rect 106178 114758 106224 114810
rect 105928 114756 105984 114758
rect 106008 114756 106064 114758
rect 106088 114756 106144 114758
rect 106168 114756 106224 114758
rect 106664 114266 106720 114268
rect 106744 114266 106800 114268
rect 106824 114266 106880 114268
rect 106904 114266 106960 114268
rect 106664 114214 106710 114266
rect 106710 114214 106720 114266
rect 106744 114214 106774 114266
rect 106774 114214 106786 114266
rect 106786 114214 106800 114266
rect 106824 114214 106838 114266
rect 106838 114214 106850 114266
rect 106850 114214 106880 114266
rect 106904 114214 106914 114266
rect 106914 114214 106960 114266
rect 106664 114212 106720 114214
rect 106744 114212 106800 114214
rect 106824 114212 106880 114214
rect 106904 114212 106960 114214
rect 105928 113722 105984 113724
rect 106008 113722 106064 113724
rect 106088 113722 106144 113724
rect 106168 113722 106224 113724
rect 105928 113670 105974 113722
rect 105974 113670 105984 113722
rect 106008 113670 106038 113722
rect 106038 113670 106050 113722
rect 106050 113670 106064 113722
rect 106088 113670 106102 113722
rect 106102 113670 106114 113722
rect 106114 113670 106144 113722
rect 106168 113670 106178 113722
rect 106178 113670 106224 113722
rect 105928 113668 105984 113670
rect 106008 113668 106064 113670
rect 106088 113668 106144 113670
rect 106168 113668 106224 113670
rect 106664 113178 106720 113180
rect 106744 113178 106800 113180
rect 106824 113178 106880 113180
rect 106904 113178 106960 113180
rect 106664 113126 106710 113178
rect 106710 113126 106720 113178
rect 106744 113126 106774 113178
rect 106774 113126 106786 113178
rect 106786 113126 106800 113178
rect 106824 113126 106838 113178
rect 106838 113126 106850 113178
rect 106850 113126 106880 113178
rect 106904 113126 106914 113178
rect 106914 113126 106960 113178
rect 106664 113124 106720 113126
rect 106744 113124 106800 113126
rect 106824 113124 106880 113126
rect 106904 113124 106960 113126
rect 105928 112634 105984 112636
rect 106008 112634 106064 112636
rect 106088 112634 106144 112636
rect 106168 112634 106224 112636
rect 105928 112582 105974 112634
rect 105974 112582 105984 112634
rect 106008 112582 106038 112634
rect 106038 112582 106050 112634
rect 106050 112582 106064 112634
rect 106088 112582 106102 112634
rect 106102 112582 106114 112634
rect 106114 112582 106144 112634
rect 106168 112582 106178 112634
rect 106178 112582 106224 112634
rect 105928 112580 105984 112582
rect 106008 112580 106064 112582
rect 106088 112580 106144 112582
rect 106168 112580 106224 112582
rect 106664 112090 106720 112092
rect 106744 112090 106800 112092
rect 106824 112090 106880 112092
rect 106904 112090 106960 112092
rect 106664 112038 106710 112090
rect 106710 112038 106720 112090
rect 106744 112038 106774 112090
rect 106774 112038 106786 112090
rect 106786 112038 106800 112090
rect 106824 112038 106838 112090
rect 106838 112038 106850 112090
rect 106850 112038 106880 112090
rect 106904 112038 106914 112090
rect 106914 112038 106960 112090
rect 106664 112036 106720 112038
rect 106744 112036 106800 112038
rect 106824 112036 106880 112038
rect 106904 112036 106960 112038
rect 105928 111546 105984 111548
rect 106008 111546 106064 111548
rect 106088 111546 106144 111548
rect 106168 111546 106224 111548
rect 105928 111494 105974 111546
rect 105974 111494 105984 111546
rect 106008 111494 106038 111546
rect 106038 111494 106050 111546
rect 106050 111494 106064 111546
rect 106088 111494 106102 111546
rect 106102 111494 106114 111546
rect 106114 111494 106144 111546
rect 106168 111494 106178 111546
rect 106178 111494 106224 111546
rect 105928 111492 105984 111494
rect 106008 111492 106064 111494
rect 106088 111492 106144 111494
rect 106168 111492 106224 111494
rect 106664 111002 106720 111004
rect 106744 111002 106800 111004
rect 106824 111002 106880 111004
rect 106904 111002 106960 111004
rect 106664 110950 106710 111002
rect 106710 110950 106720 111002
rect 106744 110950 106774 111002
rect 106774 110950 106786 111002
rect 106786 110950 106800 111002
rect 106824 110950 106838 111002
rect 106838 110950 106850 111002
rect 106850 110950 106880 111002
rect 106904 110950 106914 111002
rect 106914 110950 106960 111002
rect 106664 110948 106720 110950
rect 106744 110948 106800 110950
rect 106824 110948 106880 110950
rect 106904 110948 106960 110950
rect 105928 110458 105984 110460
rect 106008 110458 106064 110460
rect 106088 110458 106144 110460
rect 106168 110458 106224 110460
rect 105928 110406 105974 110458
rect 105974 110406 105984 110458
rect 106008 110406 106038 110458
rect 106038 110406 106050 110458
rect 106050 110406 106064 110458
rect 106088 110406 106102 110458
rect 106102 110406 106114 110458
rect 106114 110406 106144 110458
rect 106168 110406 106178 110458
rect 106178 110406 106224 110458
rect 105928 110404 105984 110406
rect 106008 110404 106064 110406
rect 106088 110404 106144 110406
rect 106168 110404 106224 110406
rect 106664 109914 106720 109916
rect 106744 109914 106800 109916
rect 106824 109914 106880 109916
rect 106904 109914 106960 109916
rect 106664 109862 106710 109914
rect 106710 109862 106720 109914
rect 106744 109862 106774 109914
rect 106774 109862 106786 109914
rect 106786 109862 106800 109914
rect 106824 109862 106838 109914
rect 106838 109862 106850 109914
rect 106850 109862 106880 109914
rect 106904 109862 106914 109914
rect 106914 109862 106960 109914
rect 106664 109860 106720 109862
rect 106744 109860 106800 109862
rect 106824 109860 106880 109862
rect 106904 109860 106960 109862
rect 105928 109370 105984 109372
rect 106008 109370 106064 109372
rect 106088 109370 106144 109372
rect 106168 109370 106224 109372
rect 105928 109318 105974 109370
rect 105974 109318 105984 109370
rect 106008 109318 106038 109370
rect 106038 109318 106050 109370
rect 106050 109318 106064 109370
rect 106088 109318 106102 109370
rect 106102 109318 106114 109370
rect 106114 109318 106144 109370
rect 106168 109318 106178 109370
rect 106178 109318 106224 109370
rect 105928 109316 105984 109318
rect 106008 109316 106064 109318
rect 106088 109316 106144 109318
rect 106168 109316 106224 109318
rect 106664 108826 106720 108828
rect 106744 108826 106800 108828
rect 106824 108826 106880 108828
rect 106904 108826 106960 108828
rect 106664 108774 106710 108826
rect 106710 108774 106720 108826
rect 106744 108774 106774 108826
rect 106774 108774 106786 108826
rect 106786 108774 106800 108826
rect 106824 108774 106838 108826
rect 106838 108774 106850 108826
rect 106850 108774 106880 108826
rect 106904 108774 106914 108826
rect 106914 108774 106960 108826
rect 106664 108772 106720 108774
rect 106744 108772 106800 108774
rect 106824 108772 106880 108774
rect 106904 108772 106960 108774
rect 105928 108282 105984 108284
rect 106008 108282 106064 108284
rect 106088 108282 106144 108284
rect 106168 108282 106224 108284
rect 105928 108230 105974 108282
rect 105974 108230 105984 108282
rect 106008 108230 106038 108282
rect 106038 108230 106050 108282
rect 106050 108230 106064 108282
rect 106088 108230 106102 108282
rect 106102 108230 106114 108282
rect 106114 108230 106144 108282
rect 106168 108230 106178 108282
rect 106178 108230 106224 108282
rect 105928 108228 105984 108230
rect 106008 108228 106064 108230
rect 106088 108228 106144 108230
rect 106168 108228 106224 108230
rect 106664 107738 106720 107740
rect 106744 107738 106800 107740
rect 106824 107738 106880 107740
rect 106904 107738 106960 107740
rect 106664 107686 106710 107738
rect 106710 107686 106720 107738
rect 106744 107686 106774 107738
rect 106774 107686 106786 107738
rect 106786 107686 106800 107738
rect 106824 107686 106838 107738
rect 106838 107686 106850 107738
rect 106850 107686 106880 107738
rect 106904 107686 106914 107738
rect 106914 107686 106960 107738
rect 106664 107684 106720 107686
rect 106744 107684 106800 107686
rect 106824 107684 106880 107686
rect 106904 107684 106960 107686
rect 105928 107194 105984 107196
rect 106008 107194 106064 107196
rect 106088 107194 106144 107196
rect 106168 107194 106224 107196
rect 105928 107142 105974 107194
rect 105974 107142 105984 107194
rect 106008 107142 106038 107194
rect 106038 107142 106050 107194
rect 106050 107142 106064 107194
rect 106088 107142 106102 107194
rect 106102 107142 106114 107194
rect 106114 107142 106144 107194
rect 106168 107142 106178 107194
rect 106178 107142 106224 107194
rect 105928 107140 105984 107142
rect 106008 107140 106064 107142
rect 106088 107140 106144 107142
rect 106168 107140 106224 107142
rect 106664 106650 106720 106652
rect 106744 106650 106800 106652
rect 106824 106650 106880 106652
rect 106904 106650 106960 106652
rect 106664 106598 106710 106650
rect 106710 106598 106720 106650
rect 106744 106598 106774 106650
rect 106774 106598 106786 106650
rect 106786 106598 106800 106650
rect 106824 106598 106838 106650
rect 106838 106598 106850 106650
rect 106850 106598 106880 106650
rect 106904 106598 106914 106650
rect 106914 106598 106960 106650
rect 106664 106596 106720 106598
rect 106744 106596 106800 106598
rect 106824 106596 106880 106598
rect 106904 106596 106960 106598
rect 105928 106106 105984 106108
rect 106008 106106 106064 106108
rect 106088 106106 106144 106108
rect 106168 106106 106224 106108
rect 105928 106054 105974 106106
rect 105974 106054 105984 106106
rect 106008 106054 106038 106106
rect 106038 106054 106050 106106
rect 106050 106054 106064 106106
rect 106088 106054 106102 106106
rect 106102 106054 106114 106106
rect 106114 106054 106144 106106
rect 106168 106054 106178 106106
rect 106178 106054 106224 106106
rect 105928 106052 105984 106054
rect 106008 106052 106064 106054
rect 106088 106052 106144 106054
rect 106168 106052 106224 106054
rect 106664 105562 106720 105564
rect 106744 105562 106800 105564
rect 106824 105562 106880 105564
rect 106904 105562 106960 105564
rect 106664 105510 106710 105562
rect 106710 105510 106720 105562
rect 106744 105510 106774 105562
rect 106774 105510 106786 105562
rect 106786 105510 106800 105562
rect 106824 105510 106838 105562
rect 106838 105510 106850 105562
rect 106850 105510 106880 105562
rect 106904 105510 106914 105562
rect 106914 105510 106960 105562
rect 106664 105508 106720 105510
rect 106744 105508 106800 105510
rect 106824 105508 106880 105510
rect 106904 105508 106960 105510
rect 105928 105018 105984 105020
rect 106008 105018 106064 105020
rect 106088 105018 106144 105020
rect 106168 105018 106224 105020
rect 105928 104966 105974 105018
rect 105974 104966 105984 105018
rect 106008 104966 106038 105018
rect 106038 104966 106050 105018
rect 106050 104966 106064 105018
rect 106088 104966 106102 105018
rect 106102 104966 106114 105018
rect 106114 104966 106144 105018
rect 106168 104966 106178 105018
rect 106178 104966 106224 105018
rect 105928 104964 105984 104966
rect 106008 104964 106064 104966
rect 106088 104964 106144 104966
rect 106168 104964 106224 104966
rect 106664 104474 106720 104476
rect 106744 104474 106800 104476
rect 106824 104474 106880 104476
rect 106904 104474 106960 104476
rect 106664 104422 106710 104474
rect 106710 104422 106720 104474
rect 106744 104422 106774 104474
rect 106774 104422 106786 104474
rect 106786 104422 106800 104474
rect 106824 104422 106838 104474
rect 106838 104422 106850 104474
rect 106850 104422 106880 104474
rect 106904 104422 106914 104474
rect 106914 104422 106960 104474
rect 106664 104420 106720 104422
rect 106744 104420 106800 104422
rect 106824 104420 106880 104422
rect 106904 104420 106960 104422
rect 105928 103930 105984 103932
rect 106008 103930 106064 103932
rect 106088 103930 106144 103932
rect 106168 103930 106224 103932
rect 105928 103878 105974 103930
rect 105974 103878 105984 103930
rect 106008 103878 106038 103930
rect 106038 103878 106050 103930
rect 106050 103878 106064 103930
rect 106088 103878 106102 103930
rect 106102 103878 106114 103930
rect 106114 103878 106144 103930
rect 106168 103878 106178 103930
rect 106178 103878 106224 103930
rect 105928 103876 105984 103878
rect 106008 103876 106064 103878
rect 106088 103876 106144 103878
rect 106168 103876 106224 103878
rect 106664 103386 106720 103388
rect 106744 103386 106800 103388
rect 106824 103386 106880 103388
rect 106904 103386 106960 103388
rect 106664 103334 106710 103386
rect 106710 103334 106720 103386
rect 106744 103334 106774 103386
rect 106774 103334 106786 103386
rect 106786 103334 106800 103386
rect 106824 103334 106838 103386
rect 106838 103334 106850 103386
rect 106850 103334 106880 103386
rect 106904 103334 106914 103386
rect 106914 103334 106960 103386
rect 106664 103332 106720 103334
rect 106744 103332 106800 103334
rect 106824 103332 106880 103334
rect 106904 103332 106960 103334
rect 105928 102842 105984 102844
rect 106008 102842 106064 102844
rect 106088 102842 106144 102844
rect 106168 102842 106224 102844
rect 105928 102790 105974 102842
rect 105974 102790 105984 102842
rect 106008 102790 106038 102842
rect 106038 102790 106050 102842
rect 106050 102790 106064 102842
rect 106088 102790 106102 102842
rect 106102 102790 106114 102842
rect 106114 102790 106144 102842
rect 106168 102790 106178 102842
rect 106178 102790 106224 102842
rect 105928 102788 105984 102790
rect 106008 102788 106064 102790
rect 106088 102788 106144 102790
rect 106168 102788 106224 102790
rect 106664 102298 106720 102300
rect 106744 102298 106800 102300
rect 106824 102298 106880 102300
rect 106904 102298 106960 102300
rect 106664 102246 106710 102298
rect 106710 102246 106720 102298
rect 106744 102246 106774 102298
rect 106774 102246 106786 102298
rect 106786 102246 106800 102298
rect 106824 102246 106838 102298
rect 106838 102246 106850 102298
rect 106850 102246 106880 102298
rect 106904 102246 106914 102298
rect 106914 102246 106960 102298
rect 106664 102244 106720 102246
rect 106744 102244 106800 102246
rect 106824 102244 106880 102246
rect 106904 102244 106960 102246
rect 105928 101754 105984 101756
rect 106008 101754 106064 101756
rect 106088 101754 106144 101756
rect 106168 101754 106224 101756
rect 105928 101702 105974 101754
rect 105974 101702 105984 101754
rect 106008 101702 106038 101754
rect 106038 101702 106050 101754
rect 106050 101702 106064 101754
rect 106088 101702 106102 101754
rect 106102 101702 106114 101754
rect 106114 101702 106144 101754
rect 106168 101702 106178 101754
rect 106178 101702 106224 101754
rect 105928 101700 105984 101702
rect 106008 101700 106064 101702
rect 106088 101700 106144 101702
rect 106168 101700 106224 101702
rect 106664 101210 106720 101212
rect 106744 101210 106800 101212
rect 106824 101210 106880 101212
rect 106904 101210 106960 101212
rect 106664 101158 106710 101210
rect 106710 101158 106720 101210
rect 106744 101158 106774 101210
rect 106774 101158 106786 101210
rect 106786 101158 106800 101210
rect 106824 101158 106838 101210
rect 106838 101158 106850 101210
rect 106850 101158 106880 101210
rect 106904 101158 106914 101210
rect 106914 101158 106960 101210
rect 106664 101156 106720 101158
rect 106744 101156 106800 101158
rect 106824 101156 106880 101158
rect 106904 101156 106960 101158
rect 105928 100666 105984 100668
rect 106008 100666 106064 100668
rect 106088 100666 106144 100668
rect 106168 100666 106224 100668
rect 105928 100614 105974 100666
rect 105974 100614 105984 100666
rect 106008 100614 106038 100666
rect 106038 100614 106050 100666
rect 106050 100614 106064 100666
rect 106088 100614 106102 100666
rect 106102 100614 106114 100666
rect 106114 100614 106144 100666
rect 106168 100614 106178 100666
rect 106178 100614 106224 100666
rect 105928 100612 105984 100614
rect 106008 100612 106064 100614
rect 106088 100612 106144 100614
rect 106168 100612 106224 100614
rect 106664 100122 106720 100124
rect 106744 100122 106800 100124
rect 106824 100122 106880 100124
rect 106904 100122 106960 100124
rect 106664 100070 106710 100122
rect 106710 100070 106720 100122
rect 106744 100070 106774 100122
rect 106774 100070 106786 100122
rect 106786 100070 106800 100122
rect 106824 100070 106838 100122
rect 106838 100070 106850 100122
rect 106850 100070 106880 100122
rect 106904 100070 106914 100122
rect 106914 100070 106960 100122
rect 106664 100068 106720 100070
rect 106744 100068 106800 100070
rect 106824 100068 106880 100070
rect 106904 100068 106960 100070
rect 105928 99578 105984 99580
rect 106008 99578 106064 99580
rect 106088 99578 106144 99580
rect 106168 99578 106224 99580
rect 105928 99526 105974 99578
rect 105974 99526 105984 99578
rect 106008 99526 106038 99578
rect 106038 99526 106050 99578
rect 106050 99526 106064 99578
rect 106088 99526 106102 99578
rect 106102 99526 106114 99578
rect 106114 99526 106144 99578
rect 106168 99526 106178 99578
rect 106178 99526 106224 99578
rect 105928 99524 105984 99526
rect 106008 99524 106064 99526
rect 106088 99524 106144 99526
rect 106168 99524 106224 99526
rect 106664 99034 106720 99036
rect 106744 99034 106800 99036
rect 106824 99034 106880 99036
rect 106904 99034 106960 99036
rect 106664 98982 106710 99034
rect 106710 98982 106720 99034
rect 106744 98982 106774 99034
rect 106774 98982 106786 99034
rect 106786 98982 106800 99034
rect 106824 98982 106838 99034
rect 106838 98982 106850 99034
rect 106850 98982 106880 99034
rect 106904 98982 106914 99034
rect 106914 98982 106960 99034
rect 106664 98980 106720 98982
rect 106744 98980 106800 98982
rect 106824 98980 106880 98982
rect 106904 98980 106960 98982
rect 105928 98490 105984 98492
rect 106008 98490 106064 98492
rect 106088 98490 106144 98492
rect 106168 98490 106224 98492
rect 105928 98438 105974 98490
rect 105974 98438 105984 98490
rect 106008 98438 106038 98490
rect 106038 98438 106050 98490
rect 106050 98438 106064 98490
rect 106088 98438 106102 98490
rect 106102 98438 106114 98490
rect 106114 98438 106144 98490
rect 106168 98438 106178 98490
rect 106178 98438 106224 98490
rect 105928 98436 105984 98438
rect 106008 98436 106064 98438
rect 106088 98436 106144 98438
rect 106168 98436 106224 98438
rect 106664 97946 106720 97948
rect 106744 97946 106800 97948
rect 106824 97946 106880 97948
rect 106904 97946 106960 97948
rect 106664 97894 106710 97946
rect 106710 97894 106720 97946
rect 106744 97894 106774 97946
rect 106774 97894 106786 97946
rect 106786 97894 106800 97946
rect 106824 97894 106838 97946
rect 106838 97894 106850 97946
rect 106850 97894 106880 97946
rect 106904 97894 106914 97946
rect 106914 97894 106960 97946
rect 106664 97892 106720 97894
rect 106744 97892 106800 97894
rect 106824 97892 106880 97894
rect 106904 97892 106960 97894
rect 105928 97402 105984 97404
rect 106008 97402 106064 97404
rect 106088 97402 106144 97404
rect 106168 97402 106224 97404
rect 105928 97350 105974 97402
rect 105974 97350 105984 97402
rect 106008 97350 106038 97402
rect 106038 97350 106050 97402
rect 106050 97350 106064 97402
rect 106088 97350 106102 97402
rect 106102 97350 106114 97402
rect 106114 97350 106144 97402
rect 106168 97350 106178 97402
rect 106178 97350 106224 97402
rect 105928 97348 105984 97350
rect 106008 97348 106064 97350
rect 106088 97348 106144 97350
rect 106168 97348 106224 97350
rect 106664 96858 106720 96860
rect 106744 96858 106800 96860
rect 106824 96858 106880 96860
rect 106904 96858 106960 96860
rect 106664 96806 106710 96858
rect 106710 96806 106720 96858
rect 106744 96806 106774 96858
rect 106774 96806 106786 96858
rect 106786 96806 106800 96858
rect 106824 96806 106838 96858
rect 106838 96806 106850 96858
rect 106850 96806 106880 96858
rect 106904 96806 106914 96858
rect 106914 96806 106960 96858
rect 106664 96804 106720 96806
rect 106744 96804 106800 96806
rect 106824 96804 106880 96806
rect 106904 96804 106960 96806
rect 105928 96314 105984 96316
rect 106008 96314 106064 96316
rect 106088 96314 106144 96316
rect 106168 96314 106224 96316
rect 105928 96262 105974 96314
rect 105974 96262 105984 96314
rect 106008 96262 106038 96314
rect 106038 96262 106050 96314
rect 106050 96262 106064 96314
rect 106088 96262 106102 96314
rect 106102 96262 106114 96314
rect 106114 96262 106144 96314
rect 106168 96262 106178 96314
rect 106178 96262 106224 96314
rect 105928 96260 105984 96262
rect 106008 96260 106064 96262
rect 106088 96260 106144 96262
rect 106168 96260 106224 96262
rect 106664 95770 106720 95772
rect 106744 95770 106800 95772
rect 106824 95770 106880 95772
rect 106904 95770 106960 95772
rect 106664 95718 106710 95770
rect 106710 95718 106720 95770
rect 106744 95718 106774 95770
rect 106774 95718 106786 95770
rect 106786 95718 106800 95770
rect 106824 95718 106838 95770
rect 106838 95718 106850 95770
rect 106850 95718 106880 95770
rect 106904 95718 106914 95770
rect 106914 95718 106960 95770
rect 106664 95716 106720 95718
rect 106744 95716 106800 95718
rect 106824 95716 106880 95718
rect 106904 95716 106960 95718
rect 105928 95226 105984 95228
rect 106008 95226 106064 95228
rect 106088 95226 106144 95228
rect 106168 95226 106224 95228
rect 105928 95174 105974 95226
rect 105974 95174 105984 95226
rect 106008 95174 106038 95226
rect 106038 95174 106050 95226
rect 106050 95174 106064 95226
rect 106088 95174 106102 95226
rect 106102 95174 106114 95226
rect 106114 95174 106144 95226
rect 106168 95174 106178 95226
rect 106178 95174 106224 95226
rect 105928 95172 105984 95174
rect 106008 95172 106064 95174
rect 106088 95172 106144 95174
rect 106168 95172 106224 95174
rect 106664 94682 106720 94684
rect 106744 94682 106800 94684
rect 106824 94682 106880 94684
rect 106904 94682 106960 94684
rect 106664 94630 106710 94682
rect 106710 94630 106720 94682
rect 106744 94630 106774 94682
rect 106774 94630 106786 94682
rect 106786 94630 106800 94682
rect 106824 94630 106838 94682
rect 106838 94630 106850 94682
rect 106850 94630 106880 94682
rect 106904 94630 106914 94682
rect 106914 94630 106960 94682
rect 106664 94628 106720 94630
rect 106744 94628 106800 94630
rect 106824 94628 106880 94630
rect 106904 94628 106960 94630
rect 105928 94138 105984 94140
rect 106008 94138 106064 94140
rect 106088 94138 106144 94140
rect 106168 94138 106224 94140
rect 105928 94086 105974 94138
rect 105974 94086 105984 94138
rect 106008 94086 106038 94138
rect 106038 94086 106050 94138
rect 106050 94086 106064 94138
rect 106088 94086 106102 94138
rect 106102 94086 106114 94138
rect 106114 94086 106144 94138
rect 106168 94086 106178 94138
rect 106178 94086 106224 94138
rect 105928 94084 105984 94086
rect 106008 94084 106064 94086
rect 106088 94084 106144 94086
rect 106168 94084 106224 94086
rect 106664 93594 106720 93596
rect 106744 93594 106800 93596
rect 106824 93594 106880 93596
rect 106904 93594 106960 93596
rect 106664 93542 106710 93594
rect 106710 93542 106720 93594
rect 106744 93542 106774 93594
rect 106774 93542 106786 93594
rect 106786 93542 106800 93594
rect 106824 93542 106838 93594
rect 106838 93542 106850 93594
rect 106850 93542 106880 93594
rect 106904 93542 106914 93594
rect 106914 93542 106960 93594
rect 106664 93540 106720 93542
rect 106744 93540 106800 93542
rect 106824 93540 106880 93542
rect 106904 93540 106960 93542
rect 105928 93050 105984 93052
rect 106008 93050 106064 93052
rect 106088 93050 106144 93052
rect 106168 93050 106224 93052
rect 105928 92998 105974 93050
rect 105974 92998 105984 93050
rect 106008 92998 106038 93050
rect 106038 92998 106050 93050
rect 106050 92998 106064 93050
rect 106088 92998 106102 93050
rect 106102 92998 106114 93050
rect 106114 92998 106144 93050
rect 106168 92998 106178 93050
rect 106178 92998 106224 93050
rect 105928 92996 105984 92998
rect 106008 92996 106064 92998
rect 106088 92996 106144 92998
rect 106168 92996 106224 92998
rect 106664 92506 106720 92508
rect 106744 92506 106800 92508
rect 106824 92506 106880 92508
rect 106904 92506 106960 92508
rect 106664 92454 106710 92506
rect 106710 92454 106720 92506
rect 106744 92454 106774 92506
rect 106774 92454 106786 92506
rect 106786 92454 106800 92506
rect 106824 92454 106838 92506
rect 106838 92454 106850 92506
rect 106850 92454 106880 92506
rect 106904 92454 106914 92506
rect 106914 92454 106960 92506
rect 106664 92452 106720 92454
rect 106744 92452 106800 92454
rect 106824 92452 106880 92454
rect 106904 92452 106960 92454
rect 105928 91962 105984 91964
rect 106008 91962 106064 91964
rect 106088 91962 106144 91964
rect 106168 91962 106224 91964
rect 105928 91910 105974 91962
rect 105974 91910 105984 91962
rect 106008 91910 106038 91962
rect 106038 91910 106050 91962
rect 106050 91910 106064 91962
rect 106088 91910 106102 91962
rect 106102 91910 106114 91962
rect 106114 91910 106144 91962
rect 106168 91910 106178 91962
rect 106178 91910 106224 91962
rect 105928 91908 105984 91910
rect 106008 91908 106064 91910
rect 106088 91908 106144 91910
rect 106168 91908 106224 91910
rect 106664 91418 106720 91420
rect 106744 91418 106800 91420
rect 106824 91418 106880 91420
rect 106904 91418 106960 91420
rect 106664 91366 106710 91418
rect 106710 91366 106720 91418
rect 106744 91366 106774 91418
rect 106774 91366 106786 91418
rect 106786 91366 106800 91418
rect 106824 91366 106838 91418
rect 106838 91366 106850 91418
rect 106850 91366 106880 91418
rect 106904 91366 106914 91418
rect 106914 91366 106960 91418
rect 106664 91364 106720 91366
rect 106744 91364 106800 91366
rect 106824 91364 106880 91366
rect 106904 91364 106960 91366
rect 105928 90874 105984 90876
rect 106008 90874 106064 90876
rect 106088 90874 106144 90876
rect 106168 90874 106224 90876
rect 105928 90822 105974 90874
rect 105974 90822 105984 90874
rect 106008 90822 106038 90874
rect 106038 90822 106050 90874
rect 106050 90822 106064 90874
rect 106088 90822 106102 90874
rect 106102 90822 106114 90874
rect 106114 90822 106144 90874
rect 106168 90822 106178 90874
rect 106178 90822 106224 90874
rect 105928 90820 105984 90822
rect 106008 90820 106064 90822
rect 106088 90820 106144 90822
rect 106168 90820 106224 90822
rect 106664 90330 106720 90332
rect 106744 90330 106800 90332
rect 106824 90330 106880 90332
rect 106904 90330 106960 90332
rect 106664 90278 106710 90330
rect 106710 90278 106720 90330
rect 106744 90278 106774 90330
rect 106774 90278 106786 90330
rect 106786 90278 106800 90330
rect 106824 90278 106838 90330
rect 106838 90278 106850 90330
rect 106850 90278 106880 90330
rect 106904 90278 106914 90330
rect 106914 90278 106960 90330
rect 106664 90276 106720 90278
rect 106744 90276 106800 90278
rect 106824 90276 106880 90278
rect 106904 90276 106960 90278
rect 105928 89786 105984 89788
rect 106008 89786 106064 89788
rect 106088 89786 106144 89788
rect 106168 89786 106224 89788
rect 105928 89734 105974 89786
rect 105974 89734 105984 89786
rect 106008 89734 106038 89786
rect 106038 89734 106050 89786
rect 106050 89734 106064 89786
rect 106088 89734 106102 89786
rect 106102 89734 106114 89786
rect 106114 89734 106144 89786
rect 106168 89734 106178 89786
rect 106178 89734 106224 89786
rect 105928 89732 105984 89734
rect 106008 89732 106064 89734
rect 106088 89732 106144 89734
rect 106168 89732 106224 89734
rect 106664 89242 106720 89244
rect 106744 89242 106800 89244
rect 106824 89242 106880 89244
rect 106904 89242 106960 89244
rect 106664 89190 106710 89242
rect 106710 89190 106720 89242
rect 106744 89190 106774 89242
rect 106774 89190 106786 89242
rect 106786 89190 106800 89242
rect 106824 89190 106838 89242
rect 106838 89190 106850 89242
rect 106850 89190 106880 89242
rect 106904 89190 106914 89242
rect 106914 89190 106960 89242
rect 106664 89188 106720 89190
rect 106744 89188 106800 89190
rect 106824 89188 106880 89190
rect 106904 89188 106960 89190
rect 105928 88698 105984 88700
rect 106008 88698 106064 88700
rect 106088 88698 106144 88700
rect 106168 88698 106224 88700
rect 105928 88646 105974 88698
rect 105974 88646 105984 88698
rect 106008 88646 106038 88698
rect 106038 88646 106050 88698
rect 106050 88646 106064 88698
rect 106088 88646 106102 88698
rect 106102 88646 106114 88698
rect 106114 88646 106144 88698
rect 106168 88646 106178 88698
rect 106178 88646 106224 88698
rect 105928 88644 105984 88646
rect 106008 88644 106064 88646
rect 106088 88644 106144 88646
rect 106168 88644 106224 88646
rect 106664 88154 106720 88156
rect 106744 88154 106800 88156
rect 106824 88154 106880 88156
rect 106904 88154 106960 88156
rect 106664 88102 106710 88154
rect 106710 88102 106720 88154
rect 106744 88102 106774 88154
rect 106774 88102 106786 88154
rect 106786 88102 106800 88154
rect 106824 88102 106838 88154
rect 106838 88102 106850 88154
rect 106850 88102 106880 88154
rect 106904 88102 106914 88154
rect 106914 88102 106960 88154
rect 106664 88100 106720 88102
rect 106744 88100 106800 88102
rect 106824 88100 106880 88102
rect 106904 88100 106960 88102
rect 105928 87610 105984 87612
rect 106008 87610 106064 87612
rect 106088 87610 106144 87612
rect 106168 87610 106224 87612
rect 105928 87558 105974 87610
rect 105974 87558 105984 87610
rect 106008 87558 106038 87610
rect 106038 87558 106050 87610
rect 106050 87558 106064 87610
rect 106088 87558 106102 87610
rect 106102 87558 106114 87610
rect 106114 87558 106144 87610
rect 106168 87558 106178 87610
rect 106178 87558 106224 87610
rect 105928 87556 105984 87558
rect 106008 87556 106064 87558
rect 106088 87556 106144 87558
rect 106168 87556 106224 87558
rect 106664 87066 106720 87068
rect 106744 87066 106800 87068
rect 106824 87066 106880 87068
rect 106904 87066 106960 87068
rect 106664 87014 106710 87066
rect 106710 87014 106720 87066
rect 106744 87014 106774 87066
rect 106774 87014 106786 87066
rect 106786 87014 106800 87066
rect 106824 87014 106838 87066
rect 106838 87014 106850 87066
rect 106850 87014 106880 87066
rect 106904 87014 106914 87066
rect 106914 87014 106960 87066
rect 106664 87012 106720 87014
rect 106744 87012 106800 87014
rect 106824 87012 106880 87014
rect 106904 87012 106960 87014
rect 105928 86522 105984 86524
rect 106008 86522 106064 86524
rect 106088 86522 106144 86524
rect 106168 86522 106224 86524
rect 105928 86470 105974 86522
rect 105974 86470 105984 86522
rect 106008 86470 106038 86522
rect 106038 86470 106050 86522
rect 106050 86470 106064 86522
rect 106088 86470 106102 86522
rect 106102 86470 106114 86522
rect 106114 86470 106144 86522
rect 106168 86470 106178 86522
rect 106178 86470 106224 86522
rect 105928 86468 105984 86470
rect 106008 86468 106064 86470
rect 106088 86468 106144 86470
rect 106168 86468 106224 86470
rect 106664 85978 106720 85980
rect 106744 85978 106800 85980
rect 106824 85978 106880 85980
rect 106904 85978 106960 85980
rect 106664 85926 106710 85978
rect 106710 85926 106720 85978
rect 106744 85926 106774 85978
rect 106774 85926 106786 85978
rect 106786 85926 106800 85978
rect 106824 85926 106838 85978
rect 106838 85926 106850 85978
rect 106850 85926 106880 85978
rect 106904 85926 106914 85978
rect 106914 85926 106960 85978
rect 106664 85924 106720 85926
rect 106744 85924 106800 85926
rect 106824 85924 106880 85926
rect 106904 85924 106960 85926
rect 105928 85434 105984 85436
rect 106008 85434 106064 85436
rect 106088 85434 106144 85436
rect 106168 85434 106224 85436
rect 105928 85382 105974 85434
rect 105974 85382 105984 85434
rect 106008 85382 106038 85434
rect 106038 85382 106050 85434
rect 106050 85382 106064 85434
rect 106088 85382 106102 85434
rect 106102 85382 106114 85434
rect 106114 85382 106144 85434
rect 106168 85382 106178 85434
rect 106178 85382 106224 85434
rect 105928 85380 105984 85382
rect 106008 85380 106064 85382
rect 106088 85380 106144 85382
rect 106168 85380 106224 85382
rect 106664 84890 106720 84892
rect 106744 84890 106800 84892
rect 106824 84890 106880 84892
rect 106904 84890 106960 84892
rect 106664 84838 106710 84890
rect 106710 84838 106720 84890
rect 106744 84838 106774 84890
rect 106774 84838 106786 84890
rect 106786 84838 106800 84890
rect 106824 84838 106838 84890
rect 106838 84838 106850 84890
rect 106850 84838 106880 84890
rect 106904 84838 106914 84890
rect 106914 84838 106960 84890
rect 106664 84836 106720 84838
rect 106744 84836 106800 84838
rect 106824 84836 106880 84838
rect 106904 84836 106960 84838
rect 105928 84346 105984 84348
rect 106008 84346 106064 84348
rect 106088 84346 106144 84348
rect 106168 84346 106224 84348
rect 105928 84294 105974 84346
rect 105974 84294 105984 84346
rect 106008 84294 106038 84346
rect 106038 84294 106050 84346
rect 106050 84294 106064 84346
rect 106088 84294 106102 84346
rect 106102 84294 106114 84346
rect 106114 84294 106144 84346
rect 106168 84294 106178 84346
rect 106178 84294 106224 84346
rect 105928 84292 105984 84294
rect 106008 84292 106064 84294
rect 106088 84292 106144 84294
rect 106168 84292 106224 84294
rect 106664 83802 106720 83804
rect 106744 83802 106800 83804
rect 106824 83802 106880 83804
rect 106904 83802 106960 83804
rect 106664 83750 106710 83802
rect 106710 83750 106720 83802
rect 106744 83750 106774 83802
rect 106774 83750 106786 83802
rect 106786 83750 106800 83802
rect 106824 83750 106838 83802
rect 106838 83750 106850 83802
rect 106850 83750 106880 83802
rect 106904 83750 106914 83802
rect 106914 83750 106960 83802
rect 106664 83748 106720 83750
rect 106744 83748 106800 83750
rect 106824 83748 106880 83750
rect 106904 83748 106960 83750
rect 105928 83258 105984 83260
rect 106008 83258 106064 83260
rect 106088 83258 106144 83260
rect 106168 83258 106224 83260
rect 105928 83206 105974 83258
rect 105974 83206 105984 83258
rect 106008 83206 106038 83258
rect 106038 83206 106050 83258
rect 106050 83206 106064 83258
rect 106088 83206 106102 83258
rect 106102 83206 106114 83258
rect 106114 83206 106144 83258
rect 106168 83206 106178 83258
rect 106178 83206 106224 83258
rect 105928 83204 105984 83206
rect 106008 83204 106064 83206
rect 106088 83204 106144 83206
rect 106168 83204 106224 83206
rect 106664 82714 106720 82716
rect 106744 82714 106800 82716
rect 106824 82714 106880 82716
rect 106904 82714 106960 82716
rect 106664 82662 106710 82714
rect 106710 82662 106720 82714
rect 106744 82662 106774 82714
rect 106774 82662 106786 82714
rect 106786 82662 106800 82714
rect 106824 82662 106838 82714
rect 106838 82662 106850 82714
rect 106850 82662 106880 82714
rect 106904 82662 106914 82714
rect 106914 82662 106960 82714
rect 106664 82660 106720 82662
rect 106744 82660 106800 82662
rect 106824 82660 106880 82662
rect 106904 82660 106960 82662
rect 105928 82170 105984 82172
rect 106008 82170 106064 82172
rect 106088 82170 106144 82172
rect 106168 82170 106224 82172
rect 105928 82118 105974 82170
rect 105974 82118 105984 82170
rect 106008 82118 106038 82170
rect 106038 82118 106050 82170
rect 106050 82118 106064 82170
rect 106088 82118 106102 82170
rect 106102 82118 106114 82170
rect 106114 82118 106144 82170
rect 106168 82118 106178 82170
rect 106178 82118 106224 82170
rect 105928 82116 105984 82118
rect 106008 82116 106064 82118
rect 106088 82116 106144 82118
rect 106168 82116 106224 82118
rect 106664 81626 106720 81628
rect 106744 81626 106800 81628
rect 106824 81626 106880 81628
rect 106904 81626 106960 81628
rect 106664 81574 106710 81626
rect 106710 81574 106720 81626
rect 106744 81574 106774 81626
rect 106774 81574 106786 81626
rect 106786 81574 106800 81626
rect 106824 81574 106838 81626
rect 106838 81574 106850 81626
rect 106850 81574 106880 81626
rect 106904 81574 106914 81626
rect 106914 81574 106960 81626
rect 106664 81572 106720 81574
rect 106744 81572 106800 81574
rect 106824 81572 106880 81574
rect 106904 81572 106960 81574
rect 105928 81082 105984 81084
rect 106008 81082 106064 81084
rect 106088 81082 106144 81084
rect 106168 81082 106224 81084
rect 105928 81030 105974 81082
rect 105974 81030 105984 81082
rect 106008 81030 106038 81082
rect 106038 81030 106050 81082
rect 106050 81030 106064 81082
rect 106088 81030 106102 81082
rect 106102 81030 106114 81082
rect 106114 81030 106144 81082
rect 106168 81030 106178 81082
rect 106178 81030 106224 81082
rect 105928 81028 105984 81030
rect 106008 81028 106064 81030
rect 106088 81028 106144 81030
rect 106168 81028 106224 81030
rect 106664 80538 106720 80540
rect 106744 80538 106800 80540
rect 106824 80538 106880 80540
rect 106904 80538 106960 80540
rect 106664 80486 106710 80538
rect 106710 80486 106720 80538
rect 106744 80486 106774 80538
rect 106774 80486 106786 80538
rect 106786 80486 106800 80538
rect 106824 80486 106838 80538
rect 106838 80486 106850 80538
rect 106850 80486 106880 80538
rect 106904 80486 106914 80538
rect 106914 80486 106960 80538
rect 106664 80484 106720 80486
rect 106744 80484 106800 80486
rect 106824 80484 106880 80486
rect 106904 80484 106960 80486
rect 105928 79994 105984 79996
rect 106008 79994 106064 79996
rect 106088 79994 106144 79996
rect 106168 79994 106224 79996
rect 105928 79942 105974 79994
rect 105974 79942 105984 79994
rect 106008 79942 106038 79994
rect 106038 79942 106050 79994
rect 106050 79942 106064 79994
rect 106088 79942 106102 79994
rect 106102 79942 106114 79994
rect 106114 79942 106144 79994
rect 106168 79942 106178 79994
rect 106178 79942 106224 79994
rect 105928 79940 105984 79942
rect 106008 79940 106064 79942
rect 106088 79940 106144 79942
rect 106168 79940 106224 79942
rect 106664 79450 106720 79452
rect 106744 79450 106800 79452
rect 106824 79450 106880 79452
rect 106904 79450 106960 79452
rect 106664 79398 106710 79450
rect 106710 79398 106720 79450
rect 106744 79398 106774 79450
rect 106774 79398 106786 79450
rect 106786 79398 106800 79450
rect 106824 79398 106838 79450
rect 106838 79398 106850 79450
rect 106850 79398 106880 79450
rect 106904 79398 106914 79450
rect 106914 79398 106960 79450
rect 106664 79396 106720 79398
rect 106744 79396 106800 79398
rect 106824 79396 106880 79398
rect 106904 79396 106960 79398
rect 105928 78906 105984 78908
rect 106008 78906 106064 78908
rect 106088 78906 106144 78908
rect 106168 78906 106224 78908
rect 105928 78854 105974 78906
rect 105974 78854 105984 78906
rect 106008 78854 106038 78906
rect 106038 78854 106050 78906
rect 106050 78854 106064 78906
rect 106088 78854 106102 78906
rect 106102 78854 106114 78906
rect 106114 78854 106144 78906
rect 106168 78854 106178 78906
rect 106178 78854 106224 78906
rect 105928 78852 105984 78854
rect 106008 78852 106064 78854
rect 106088 78852 106144 78854
rect 106168 78852 106224 78854
rect 106664 78362 106720 78364
rect 106744 78362 106800 78364
rect 106824 78362 106880 78364
rect 106904 78362 106960 78364
rect 106664 78310 106710 78362
rect 106710 78310 106720 78362
rect 106744 78310 106774 78362
rect 106774 78310 106786 78362
rect 106786 78310 106800 78362
rect 106824 78310 106838 78362
rect 106838 78310 106850 78362
rect 106850 78310 106880 78362
rect 106904 78310 106914 78362
rect 106914 78310 106960 78362
rect 106664 78308 106720 78310
rect 106744 78308 106800 78310
rect 106824 78308 106880 78310
rect 106904 78308 106960 78310
rect 105928 77818 105984 77820
rect 106008 77818 106064 77820
rect 106088 77818 106144 77820
rect 106168 77818 106224 77820
rect 105928 77766 105974 77818
rect 105974 77766 105984 77818
rect 106008 77766 106038 77818
rect 106038 77766 106050 77818
rect 106050 77766 106064 77818
rect 106088 77766 106102 77818
rect 106102 77766 106114 77818
rect 106114 77766 106144 77818
rect 106168 77766 106178 77818
rect 106178 77766 106224 77818
rect 105928 77764 105984 77766
rect 106008 77764 106064 77766
rect 106088 77764 106144 77766
rect 106168 77764 106224 77766
rect 106664 77274 106720 77276
rect 106744 77274 106800 77276
rect 106824 77274 106880 77276
rect 106904 77274 106960 77276
rect 106664 77222 106710 77274
rect 106710 77222 106720 77274
rect 106744 77222 106774 77274
rect 106774 77222 106786 77274
rect 106786 77222 106800 77274
rect 106824 77222 106838 77274
rect 106838 77222 106850 77274
rect 106850 77222 106880 77274
rect 106904 77222 106914 77274
rect 106914 77222 106960 77274
rect 106664 77220 106720 77222
rect 106744 77220 106800 77222
rect 106824 77220 106880 77222
rect 106904 77220 106960 77222
rect 100390 74432 100446 74488
rect 100206 74196 100208 74216
rect 100208 74196 100260 74216
rect 100260 74196 100262 74216
rect 100206 74160 100262 74196
rect 96380 69114 96436 69116
rect 96460 69114 96516 69116
rect 96540 69114 96596 69116
rect 96620 69114 96676 69116
rect 96380 69062 96426 69114
rect 96426 69062 96436 69114
rect 96460 69062 96490 69114
rect 96490 69062 96502 69114
rect 96502 69062 96516 69114
rect 96540 69062 96554 69114
rect 96554 69062 96566 69114
rect 96566 69062 96596 69114
rect 96620 69062 96630 69114
rect 96630 69062 96676 69114
rect 96380 69060 96436 69062
rect 96460 69060 96516 69062
rect 96540 69060 96596 69062
rect 96620 69060 96676 69062
rect 96380 68026 96436 68028
rect 96460 68026 96516 68028
rect 96540 68026 96596 68028
rect 96620 68026 96676 68028
rect 96380 67974 96426 68026
rect 96426 67974 96436 68026
rect 96460 67974 96490 68026
rect 96490 67974 96502 68026
rect 96502 67974 96516 68026
rect 96540 67974 96554 68026
rect 96554 67974 96566 68026
rect 96566 67974 96596 68026
rect 96620 67974 96630 68026
rect 96630 67974 96676 68026
rect 96380 67972 96436 67974
rect 96460 67972 96516 67974
rect 96540 67972 96596 67974
rect 96620 67972 96676 67974
rect 96380 66938 96436 66940
rect 96460 66938 96516 66940
rect 96540 66938 96596 66940
rect 96620 66938 96676 66940
rect 96380 66886 96426 66938
rect 96426 66886 96436 66938
rect 96460 66886 96490 66938
rect 96490 66886 96502 66938
rect 96502 66886 96516 66938
rect 96540 66886 96554 66938
rect 96554 66886 96566 66938
rect 96566 66886 96596 66938
rect 96620 66886 96630 66938
rect 96630 66886 96676 66938
rect 96380 66884 96436 66886
rect 96460 66884 96516 66886
rect 96540 66884 96596 66886
rect 96620 66884 96676 66886
rect 97040 69658 97096 69660
rect 97120 69658 97176 69660
rect 97200 69658 97256 69660
rect 97280 69658 97336 69660
rect 97040 69606 97086 69658
rect 97086 69606 97096 69658
rect 97120 69606 97150 69658
rect 97150 69606 97162 69658
rect 97162 69606 97176 69658
rect 97200 69606 97214 69658
rect 97214 69606 97226 69658
rect 97226 69606 97256 69658
rect 97280 69606 97290 69658
rect 97290 69606 97336 69658
rect 97040 69604 97096 69606
rect 97120 69604 97176 69606
rect 97200 69604 97256 69606
rect 97280 69604 97336 69606
rect 97040 68570 97096 68572
rect 97120 68570 97176 68572
rect 97200 68570 97256 68572
rect 97280 68570 97336 68572
rect 97040 68518 97086 68570
rect 97086 68518 97096 68570
rect 97120 68518 97150 68570
rect 97150 68518 97162 68570
rect 97162 68518 97176 68570
rect 97200 68518 97214 68570
rect 97214 68518 97226 68570
rect 97226 68518 97256 68570
rect 97280 68518 97290 68570
rect 97290 68518 97336 68570
rect 97040 68516 97096 68518
rect 97120 68516 97176 68518
rect 97200 68516 97256 68518
rect 97280 68516 97336 68518
rect 97538 67632 97594 67688
rect 97040 67482 97096 67484
rect 97120 67482 97176 67484
rect 97200 67482 97256 67484
rect 97280 67482 97336 67484
rect 97040 67430 97086 67482
rect 97086 67430 97096 67482
rect 97120 67430 97150 67482
rect 97150 67430 97162 67482
rect 97162 67430 97176 67482
rect 97200 67430 97214 67482
rect 97214 67430 97226 67482
rect 97226 67430 97256 67482
rect 97280 67430 97290 67482
rect 97290 67430 97336 67482
rect 97040 67428 97096 67430
rect 97120 67428 97176 67430
rect 97200 67428 97256 67430
rect 97280 67428 97336 67430
rect 97040 66394 97096 66396
rect 97120 66394 97176 66396
rect 97200 66394 97256 66396
rect 97280 66394 97336 66396
rect 97040 66342 97086 66394
rect 97086 66342 97096 66394
rect 97120 66342 97150 66394
rect 97150 66342 97162 66394
rect 97162 66342 97176 66394
rect 97200 66342 97214 66394
rect 97214 66342 97226 66394
rect 97226 66342 97256 66394
rect 97280 66342 97290 66394
rect 97290 66342 97336 66394
rect 97040 66340 97096 66342
rect 97120 66340 97176 66342
rect 97200 66340 97256 66342
rect 97280 66340 97336 66342
rect 98826 70896 98882 70952
rect 100574 74196 100576 74216
rect 100576 74196 100628 74216
rect 100628 74196 100630 74216
rect 100574 74160 100630 74196
rect 100022 69944 100078 70000
rect 101034 70932 101036 70952
rect 101036 70932 101088 70952
rect 101088 70932 101090 70952
rect 101034 70896 101090 70932
rect 100298 68892 100300 68912
rect 100300 68892 100352 68912
rect 100352 68892 100354 68912
rect 100298 68856 100354 68892
rect 102506 73752 102562 73808
rect 108486 80316 108488 80336
rect 108488 80316 108540 80336
rect 108540 80316 108542 80336
rect 108486 80280 108542 80316
rect 108394 79600 108450 79656
rect 108394 78956 108396 78976
rect 108396 78956 108448 78976
rect 108448 78956 108450 78976
rect 108394 78920 108450 78956
rect 108394 78240 108450 78296
rect 108394 77560 108450 77616
rect 108394 76900 108450 76936
rect 108394 76880 108396 76900
rect 108396 76880 108448 76900
rect 108448 76880 108450 76900
rect 108394 76236 108396 76256
rect 108396 76236 108448 76256
rect 108448 76236 108450 76256
rect 108394 76200 108450 76236
rect 108394 75520 108450 75576
rect 108394 74840 108450 74896
rect 104714 73772 104770 73808
rect 104714 73752 104716 73772
rect 104716 73752 104768 73772
rect 104768 73752 104770 73772
rect 108394 74160 108450 74216
rect 108486 73480 108542 73536
rect 103518 70896 103574 70952
rect 100850 68332 100906 68368
rect 100850 68312 100852 68332
rect 100852 68312 100904 68332
rect 100904 68312 100906 68332
rect 100850 67632 100906 67688
rect 102138 67768 102194 67824
rect 102966 67804 102968 67824
rect 102968 67804 103020 67824
rect 103020 67804 103022 67824
rect 102966 67768 103022 67804
rect 96380 65850 96436 65852
rect 96460 65850 96516 65852
rect 96540 65850 96596 65852
rect 96620 65850 96676 65852
rect 96380 65798 96426 65850
rect 96426 65798 96436 65850
rect 96460 65798 96490 65850
rect 96490 65798 96502 65850
rect 96502 65798 96516 65850
rect 96540 65798 96554 65850
rect 96554 65798 96566 65850
rect 96566 65798 96596 65850
rect 96620 65798 96630 65850
rect 96630 65798 96676 65850
rect 96380 65796 96436 65798
rect 96460 65796 96516 65798
rect 96540 65796 96596 65798
rect 96620 65796 96676 65798
rect 95882 64096 95938 64152
rect 77850 63824 77906 63880
rect 104898 68332 104954 68368
rect 108486 72800 108542 72856
rect 108486 72120 108542 72176
rect 108486 71440 108542 71496
rect 108486 70760 108542 70816
rect 104898 68312 104900 68332
rect 104900 68312 104952 68332
rect 104952 68312 104954 68332
rect 108486 70080 108542 70136
rect 108486 69400 108542 69456
rect 108486 67360 108542 67416
rect 102598 25100 102600 25120
rect 102600 25100 102652 25120
rect 102652 25100 102654 25120
rect 102230 25032 102286 25088
rect 102598 25064 102654 25100
rect 102782 23468 102784 23488
rect 102784 23468 102836 23488
rect 102836 23468 102838 23488
rect 102782 23432 102838 23468
rect 102138 22204 102194 22260
rect 23478 9696 23534 9752
rect 25778 9696 25834 9752
rect 28170 9696 28226 9752
rect 29550 9696 29606 9752
rect 30470 9696 30526 9752
rect 16026 9596 16028 9616
rect 16028 9596 16080 9616
rect 16080 9596 16082 9616
rect 16026 9560 16082 9596
rect 1398 5480 1454 5536
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1306 4800 1362 4856
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 24674 9560 24730 9616
rect 26698 8880 26754 8936
rect 90638 9560 90694 9616
rect 90822 9560 90878 9616
rect 90546 8336 90602 8392
rect 31666 8200 31722 8256
rect 32954 8200 33010 8256
rect 34242 8200 34298 8256
rect 35438 8200 35494 8256
rect 36358 8200 36414 8256
rect 37462 8200 37518 8256
rect 38750 8200 38806 8256
rect 41326 8200 41382 8256
rect 42154 8200 42210 8256
rect 43442 8200 43498 8256
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 39946 4528 40002 4584
rect 66320 7642 66376 7644
rect 66400 7642 66456 7644
rect 66480 7642 66536 7644
rect 66560 7642 66616 7644
rect 66320 7590 66366 7642
rect 66366 7590 66376 7642
rect 66400 7590 66430 7642
rect 66430 7590 66442 7642
rect 66442 7590 66456 7642
rect 66480 7590 66494 7642
rect 66494 7590 66506 7642
rect 66506 7590 66536 7642
rect 66560 7590 66570 7642
rect 66570 7590 66616 7642
rect 66320 7588 66376 7590
rect 66400 7588 66456 7590
rect 66480 7588 66536 7590
rect 66560 7588 66616 7590
rect 106664 66394 106720 66396
rect 106744 66394 106800 66396
rect 106824 66394 106880 66396
rect 106904 66394 106960 66396
rect 106664 66342 106710 66394
rect 106710 66342 106720 66394
rect 106744 66342 106774 66394
rect 106774 66342 106786 66394
rect 106786 66342 106800 66394
rect 106824 66342 106838 66394
rect 106838 66342 106850 66394
rect 106850 66342 106880 66394
rect 106904 66342 106914 66394
rect 106914 66342 106960 66394
rect 106664 66340 106720 66342
rect 106744 66340 106800 66342
rect 106824 66340 106880 66342
rect 106904 66340 106960 66342
rect 105928 65850 105984 65852
rect 106008 65850 106064 65852
rect 106088 65850 106144 65852
rect 106168 65850 106224 65852
rect 105928 65798 105974 65850
rect 105974 65798 105984 65850
rect 106008 65798 106038 65850
rect 106038 65798 106050 65850
rect 106050 65798 106064 65850
rect 106088 65798 106102 65850
rect 106102 65798 106114 65850
rect 106114 65798 106144 65850
rect 106168 65798 106178 65850
rect 106178 65798 106224 65850
rect 105928 65796 105984 65798
rect 106008 65796 106064 65798
rect 106088 65796 106144 65798
rect 106168 65796 106224 65798
rect 106664 65306 106720 65308
rect 106744 65306 106800 65308
rect 106824 65306 106880 65308
rect 106904 65306 106960 65308
rect 106664 65254 106710 65306
rect 106710 65254 106720 65306
rect 106744 65254 106774 65306
rect 106774 65254 106786 65306
rect 106786 65254 106800 65306
rect 106824 65254 106838 65306
rect 106838 65254 106850 65306
rect 106850 65254 106880 65306
rect 106904 65254 106914 65306
rect 106914 65254 106960 65306
rect 106664 65252 106720 65254
rect 106744 65252 106800 65254
rect 106824 65252 106880 65254
rect 106904 65252 106960 65254
rect 105928 64762 105984 64764
rect 106008 64762 106064 64764
rect 106088 64762 106144 64764
rect 106168 64762 106224 64764
rect 105928 64710 105974 64762
rect 105974 64710 105984 64762
rect 106008 64710 106038 64762
rect 106038 64710 106050 64762
rect 106050 64710 106064 64762
rect 106088 64710 106102 64762
rect 106102 64710 106114 64762
rect 106114 64710 106144 64762
rect 106168 64710 106178 64762
rect 106178 64710 106224 64762
rect 105928 64708 105984 64710
rect 106008 64708 106064 64710
rect 106088 64708 106144 64710
rect 106168 64708 106224 64710
rect 106664 64218 106720 64220
rect 106744 64218 106800 64220
rect 106824 64218 106880 64220
rect 106904 64218 106960 64220
rect 106664 64166 106710 64218
rect 106710 64166 106720 64218
rect 106744 64166 106774 64218
rect 106774 64166 106786 64218
rect 106786 64166 106800 64218
rect 106824 64166 106838 64218
rect 106838 64166 106850 64218
rect 106850 64166 106880 64218
rect 106904 64166 106914 64218
rect 106914 64166 106960 64218
rect 106664 64164 106720 64166
rect 106744 64164 106800 64166
rect 106824 64164 106880 64166
rect 106904 64164 106960 64166
rect 105928 63674 105984 63676
rect 106008 63674 106064 63676
rect 106088 63674 106144 63676
rect 106168 63674 106224 63676
rect 105928 63622 105974 63674
rect 105974 63622 105984 63674
rect 106008 63622 106038 63674
rect 106038 63622 106050 63674
rect 106050 63622 106064 63674
rect 106088 63622 106102 63674
rect 106102 63622 106114 63674
rect 106114 63622 106144 63674
rect 106168 63622 106178 63674
rect 106178 63622 106224 63674
rect 105928 63620 105984 63622
rect 106008 63620 106064 63622
rect 106088 63620 106144 63622
rect 106168 63620 106224 63622
rect 106664 63130 106720 63132
rect 106744 63130 106800 63132
rect 106824 63130 106880 63132
rect 106904 63130 106960 63132
rect 106664 63078 106710 63130
rect 106710 63078 106720 63130
rect 106744 63078 106774 63130
rect 106774 63078 106786 63130
rect 106786 63078 106800 63130
rect 106824 63078 106838 63130
rect 106838 63078 106850 63130
rect 106850 63078 106880 63130
rect 106904 63078 106914 63130
rect 106914 63078 106960 63130
rect 106664 63076 106720 63078
rect 106744 63076 106800 63078
rect 106824 63076 106880 63078
rect 106904 63076 106960 63078
rect 105928 62586 105984 62588
rect 106008 62586 106064 62588
rect 106088 62586 106144 62588
rect 106168 62586 106224 62588
rect 105928 62534 105974 62586
rect 105974 62534 105984 62586
rect 106008 62534 106038 62586
rect 106038 62534 106050 62586
rect 106050 62534 106064 62586
rect 106088 62534 106102 62586
rect 106102 62534 106114 62586
rect 106114 62534 106144 62586
rect 106168 62534 106178 62586
rect 106178 62534 106224 62586
rect 105928 62532 105984 62534
rect 106008 62532 106064 62534
rect 106088 62532 106144 62534
rect 106168 62532 106224 62534
rect 106664 62042 106720 62044
rect 106744 62042 106800 62044
rect 106824 62042 106880 62044
rect 106904 62042 106960 62044
rect 106664 61990 106710 62042
rect 106710 61990 106720 62042
rect 106744 61990 106774 62042
rect 106774 61990 106786 62042
rect 106786 61990 106800 62042
rect 106824 61990 106838 62042
rect 106838 61990 106850 62042
rect 106850 61990 106880 62042
rect 106904 61990 106914 62042
rect 106914 61990 106960 62042
rect 106664 61988 106720 61990
rect 106744 61988 106800 61990
rect 106824 61988 106880 61990
rect 106904 61988 106960 61990
rect 105928 61498 105984 61500
rect 106008 61498 106064 61500
rect 106088 61498 106144 61500
rect 106168 61498 106224 61500
rect 105928 61446 105974 61498
rect 105974 61446 105984 61498
rect 106008 61446 106038 61498
rect 106038 61446 106050 61498
rect 106050 61446 106064 61498
rect 106088 61446 106102 61498
rect 106102 61446 106114 61498
rect 106114 61446 106144 61498
rect 106168 61446 106178 61498
rect 106178 61446 106224 61498
rect 105928 61444 105984 61446
rect 106008 61444 106064 61446
rect 106088 61444 106144 61446
rect 106168 61444 106224 61446
rect 106664 60954 106720 60956
rect 106744 60954 106800 60956
rect 106824 60954 106880 60956
rect 106904 60954 106960 60956
rect 106664 60902 106710 60954
rect 106710 60902 106720 60954
rect 106744 60902 106774 60954
rect 106774 60902 106786 60954
rect 106786 60902 106800 60954
rect 106824 60902 106838 60954
rect 106838 60902 106850 60954
rect 106850 60902 106880 60954
rect 106904 60902 106914 60954
rect 106914 60902 106960 60954
rect 106664 60900 106720 60902
rect 106744 60900 106800 60902
rect 106824 60900 106880 60902
rect 106904 60900 106960 60902
rect 105928 60410 105984 60412
rect 106008 60410 106064 60412
rect 106088 60410 106144 60412
rect 106168 60410 106224 60412
rect 105928 60358 105974 60410
rect 105974 60358 105984 60410
rect 106008 60358 106038 60410
rect 106038 60358 106050 60410
rect 106050 60358 106064 60410
rect 106088 60358 106102 60410
rect 106102 60358 106114 60410
rect 106114 60358 106144 60410
rect 106168 60358 106178 60410
rect 106178 60358 106224 60410
rect 105928 60356 105984 60358
rect 106008 60356 106064 60358
rect 106088 60356 106144 60358
rect 106168 60356 106224 60358
rect 106664 59866 106720 59868
rect 106744 59866 106800 59868
rect 106824 59866 106880 59868
rect 106904 59866 106960 59868
rect 106664 59814 106710 59866
rect 106710 59814 106720 59866
rect 106744 59814 106774 59866
rect 106774 59814 106786 59866
rect 106786 59814 106800 59866
rect 106824 59814 106838 59866
rect 106838 59814 106850 59866
rect 106850 59814 106880 59866
rect 106904 59814 106914 59866
rect 106914 59814 106960 59866
rect 106664 59812 106720 59814
rect 106744 59812 106800 59814
rect 106824 59812 106880 59814
rect 106904 59812 106960 59814
rect 104346 59744 104402 59800
rect 105928 59322 105984 59324
rect 106008 59322 106064 59324
rect 106088 59322 106144 59324
rect 106168 59322 106224 59324
rect 105928 59270 105974 59322
rect 105974 59270 105984 59322
rect 106008 59270 106038 59322
rect 106038 59270 106050 59322
rect 106050 59270 106064 59322
rect 106088 59270 106102 59322
rect 106102 59270 106114 59322
rect 106114 59270 106144 59322
rect 106168 59270 106178 59322
rect 106178 59270 106224 59322
rect 105928 59268 105984 59270
rect 106008 59268 106064 59270
rect 106088 59268 106144 59270
rect 106168 59268 106224 59270
rect 106664 58778 106720 58780
rect 106744 58778 106800 58780
rect 106824 58778 106880 58780
rect 106904 58778 106960 58780
rect 106664 58726 106710 58778
rect 106710 58726 106720 58778
rect 106744 58726 106774 58778
rect 106774 58726 106786 58778
rect 106786 58726 106800 58778
rect 106824 58726 106838 58778
rect 106838 58726 106850 58778
rect 106850 58726 106880 58778
rect 106904 58726 106914 58778
rect 106914 58726 106960 58778
rect 106664 58724 106720 58726
rect 106744 58724 106800 58726
rect 106824 58724 106880 58726
rect 106904 58724 106960 58726
rect 105928 58234 105984 58236
rect 106008 58234 106064 58236
rect 106088 58234 106144 58236
rect 106168 58234 106224 58236
rect 105928 58182 105974 58234
rect 105974 58182 105984 58234
rect 106008 58182 106038 58234
rect 106038 58182 106050 58234
rect 106050 58182 106064 58234
rect 106088 58182 106102 58234
rect 106102 58182 106114 58234
rect 106114 58182 106144 58234
rect 106168 58182 106178 58234
rect 106178 58182 106224 58234
rect 105928 58180 105984 58182
rect 106008 58180 106064 58182
rect 106088 58180 106144 58182
rect 106168 58180 106224 58182
rect 106664 57690 106720 57692
rect 106744 57690 106800 57692
rect 106824 57690 106880 57692
rect 106904 57690 106960 57692
rect 106664 57638 106710 57690
rect 106710 57638 106720 57690
rect 106744 57638 106774 57690
rect 106774 57638 106786 57690
rect 106786 57638 106800 57690
rect 106824 57638 106838 57690
rect 106838 57638 106850 57690
rect 106850 57638 106880 57690
rect 106904 57638 106914 57690
rect 106914 57638 106960 57690
rect 106664 57636 106720 57638
rect 106744 57636 106800 57638
rect 106824 57636 106880 57638
rect 106904 57636 106960 57638
rect 105928 57146 105984 57148
rect 106008 57146 106064 57148
rect 106088 57146 106144 57148
rect 106168 57146 106224 57148
rect 105928 57094 105974 57146
rect 105974 57094 105984 57146
rect 106008 57094 106038 57146
rect 106038 57094 106050 57146
rect 106050 57094 106064 57146
rect 106088 57094 106102 57146
rect 106102 57094 106114 57146
rect 106114 57094 106144 57146
rect 106168 57094 106178 57146
rect 106178 57094 106224 57146
rect 105928 57092 105984 57094
rect 106008 57092 106064 57094
rect 106088 57092 106144 57094
rect 106168 57092 106224 57094
rect 106664 56602 106720 56604
rect 106744 56602 106800 56604
rect 106824 56602 106880 56604
rect 106904 56602 106960 56604
rect 106664 56550 106710 56602
rect 106710 56550 106720 56602
rect 106744 56550 106774 56602
rect 106774 56550 106786 56602
rect 106786 56550 106800 56602
rect 106824 56550 106838 56602
rect 106838 56550 106850 56602
rect 106850 56550 106880 56602
rect 106904 56550 106914 56602
rect 106914 56550 106960 56602
rect 106664 56548 106720 56550
rect 106744 56548 106800 56550
rect 106824 56548 106880 56550
rect 106904 56548 106960 56550
rect 105928 56058 105984 56060
rect 106008 56058 106064 56060
rect 106088 56058 106144 56060
rect 106168 56058 106224 56060
rect 105928 56006 105974 56058
rect 105974 56006 105984 56058
rect 106008 56006 106038 56058
rect 106038 56006 106050 56058
rect 106050 56006 106064 56058
rect 106088 56006 106102 56058
rect 106102 56006 106114 56058
rect 106114 56006 106144 56058
rect 106168 56006 106178 56058
rect 106178 56006 106224 56058
rect 105928 56004 105984 56006
rect 106008 56004 106064 56006
rect 106088 56004 106144 56006
rect 106168 56004 106224 56006
rect 106664 55514 106720 55516
rect 106744 55514 106800 55516
rect 106824 55514 106880 55516
rect 106904 55514 106960 55516
rect 106664 55462 106710 55514
rect 106710 55462 106720 55514
rect 106744 55462 106774 55514
rect 106774 55462 106786 55514
rect 106786 55462 106800 55514
rect 106824 55462 106838 55514
rect 106838 55462 106850 55514
rect 106850 55462 106880 55514
rect 106904 55462 106914 55514
rect 106914 55462 106960 55514
rect 106664 55460 106720 55462
rect 106744 55460 106800 55462
rect 106824 55460 106880 55462
rect 106904 55460 106960 55462
rect 105928 54970 105984 54972
rect 106008 54970 106064 54972
rect 106088 54970 106144 54972
rect 106168 54970 106224 54972
rect 105928 54918 105974 54970
rect 105974 54918 105984 54970
rect 106008 54918 106038 54970
rect 106038 54918 106050 54970
rect 106050 54918 106064 54970
rect 106088 54918 106102 54970
rect 106102 54918 106114 54970
rect 106114 54918 106144 54970
rect 106168 54918 106178 54970
rect 106178 54918 106224 54970
rect 105928 54916 105984 54918
rect 106008 54916 106064 54918
rect 106088 54916 106144 54918
rect 106168 54916 106224 54918
rect 106664 54426 106720 54428
rect 106744 54426 106800 54428
rect 106824 54426 106880 54428
rect 106904 54426 106960 54428
rect 106664 54374 106710 54426
rect 106710 54374 106720 54426
rect 106744 54374 106774 54426
rect 106774 54374 106786 54426
rect 106786 54374 106800 54426
rect 106824 54374 106838 54426
rect 106838 54374 106850 54426
rect 106850 54374 106880 54426
rect 106904 54374 106914 54426
rect 106914 54374 106960 54426
rect 106664 54372 106720 54374
rect 106744 54372 106800 54374
rect 106824 54372 106880 54374
rect 106904 54372 106960 54374
rect 105928 53882 105984 53884
rect 106008 53882 106064 53884
rect 106088 53882 106144 53884
rect 106168 53882 106224 53884
rect 105928 53830 105974 53882
rect 105974 53830 105984 53882
rect 106008 53830 106038 53882
rect 106038 53830 106050 53882
rect 106050 53830 106064 53882
rect 106088 53830 106102 53882
rect 106102 53830 106114 53882
rect 106114 53830 106144 53882
rect 106168 53830 106178 53882
rect 106178 53830 106224 53882
rect 105928 53828 105984 53830
rect 106008 53828 106064 53830
rect 106088 53828 106144 53830
rect 106168 53828 106224 53830
rect 106664 53338 106720 53340
rect 106744 53338 106800 53340
rect 106824 53338 106880 53340
rect 106904 53338 106960 53340
rect 106664 53286 106710 53338
rect 106710 53286 106720 53338
rect 106744 53286 106774 53338
rect 106774 53286 106786 53338
rect 106786 53286 106800 53338
rect 106824 53286 106838 53338
rect 106838 53286 106850 53338
rect 106850 53286 106880 53338
rect 106904 53286 106914 53338
rect 106914 53286 106960 53338
rect 106664 53284 106720 53286
rect 106744 53284 106800 53286
rect 106824 53284 106880 53286
rect 106904 53284 106960 53286
rect 105928 52794 105984 52796
rect 106008 52794 106064 52796
rect 106088 52794 106144 52796
rect 106168 52794 106224 52796
rect 105928 52742 105974 52794
rect 105974 52742 105984 52794
rect 106008 52742 106038 52794
rect 106038 52742 106050 52794
rect 106050 52742 106064 52794
rect 106088 52742 106102 52794
rect 106102 52742 106114 52794
rect 106114 52742 106144 52794
rect 106168 52742 106178 52794
rect 106178 52742 106224 52794
rect 105928 52740 105984 52742
rect 106008 52740 106064 52742
rect 106088 52740 106144 52742
rect 106168 52740 106224 52742
rect 106664 52250 106720 52252
rect 106744 52250 106800 52252
rect 106824 52250 106880 52252
rect 106904 52250 106960 52252
rect 106664 52198 106710 52250
rect 106710 52198 106720 52250
rect 106744 52198 106774 52250
rect 106774 52198 106786 52250
rect 106786 52198 106800 52250
rect 106824 52198 106838 52250
rect 106838 52198 106850 52250
rect 106850 52198 106880 52250
rect 106904 52198 106914 52250
rect 106914 52198 106960 52250
rect 106664 52196 106720 52198
rect 106744 52196 106800 52198
rect 106824 52196 106880 52198
rect 106904 52196 106960 52198
rect 105928 51706 105984 51708
rect 106008 51706 106064 51708
rect 106088 51706 106144 51708
rect 106168 51706 106224 51708
rect 105928 51654 105974 51706
rect 105974 51654 105984 51706
rect 106008 51654 106038 51706
rect 106038 51654 106050 51706
rect 106050 51654 106064 51706
rect 106088 51654 106102 51706
rect 106102 51654 106114 51706
rect 106114 51654 106144 51706
rect 106168 51654 106178 51706
rect 106178 51654 106224 51706
rect 105928 51652 105984 51654
rect 106008 51652 106064 51654
rect 106088 51652 106144 51654
rect 106168 51652 106224 51654
rect 106664 51162 106720 51164
rect 106744 51162 106800 51164
rect 106824 51162 106880 51164
rect 106904 51162 106960 51164
rect 106664 51110 106710 51162
rect 106710 51110 106720 51162
rect 106744 51110 106774 51162
rect 106774 51110 106786 51162
rect 106786 51110 106800 51162
rect 106824 51110 106838 51162
rect 106838 51110 106850 51162
rect 106850 51110 106880 51162
rect 106904 51110 106914 51162
rect 106914 51110 106960 51162
rect 106664 51108 106720 51110
rect 106744 51108 106800 51110
rect 106824 51108 106880 51110
rect 106904 51108 106960 51110
rect 105928 50618 105984 50620
rect 106008 50618 106064 50620
rect 106088 50618 106144 50620
rect 106168 50618 106224 50620
rect 105928 50566 105974 50618
rect 105974 50566 105984 50618
rect 106008 50566 106038 50618
rect 106038 50566 106050 50618
rect 106050 50566 106064 50618
rect 106088 50566 106102 50618
rect 106102 50566 106114 50618
rect 106114 50566 106144 50618
rect 106168 50566 106178 50618
rect 106178 50566 106224 50618
rect 105928 50564 105984 50566
rect 106008 50564 106064 50566
rect 106088 50564 106144 50566
rect 106168 50564 106224 50566
rect 106664 50074 106720 50076
rect 106744 50074 106800 50076
rect 106824 50074 106880 50076
rect 106904 50074 106960 50076
rect 106664 50022 106710 50074
rect 106710 50022 106720 50074
rect 106744 50022 106774 50074
rect 106774 50022 106786 50074
rect 106786 50022 106800 50074
rect 106824 50022 106838 50074
rect 106838 50022 106850 50074
rect 106850 50022 106880 50074
rect 106904 50022 106914 50074
rect 106914 50022 106960 50074
rect 106664 50020 106720 50022
rect 106744 50020 106800 50022
rect 106824 50020 106880 50022
rect 106904 50020 106960 50022
rect 105928 49530 105984 49532
rect 106008 49530 106064 49532
rect 106088 49530 106144 49532
rect 106168 49530 106224 49532
rect 105928 49478 105974 49530
rect 105974 49478 105984 49530
rect 106008 49478 106038 49530
rect 106038 49478 106050 49530
rect 106050 49478 106064 49530
rect 106088 49478 106102 49530
rect 106102 49478 106114 49530
rect 106114 49478 106144 49530
rect 106168 49478 106178 49530
rect 106178 49478 106224 49530
rect 105928 49476 105984 49478
rect 106008 49476 106064 49478
rect 106088 49476 106144 49478
rect 106168 49476 106224 49478
rect 106664 48986 106720 48988
rect 106744 48986 106800 48988
rect 106824 48986 106880 48988
rect 106904 48986 106960 48988
rect 106664 48934 106710 48986
rect 106710 48934 106720 48986
rect 106744 48934 106774 48986
rect 106774 48934 106786 48986
rect 106786 48934 106800 48986
rect 106824 48934 106838 48986
rect 106838 48934 106850 48986
rect 106850 48934 106880 48986
rect 106904 48934 106914 48986
rect 106914 48934 106960 48986
rect 106664 48932 106720 48934
rect 106744 48932 106800 48934
rect 106824 48932 106880 48934
rect 106904 48932 106960 48934
rect 105928 48442 105984 48444
rect 106008 48442 106064 48444
rect 106088 48442 106144 48444
rect 106168 48442 106224 48444
rect 105928 48390 105974 48442
rect 105974 48390 105984 48442
rect 106008 48390 106038 48442
rect 106038 48390 106050 48442
rect 106050 48390 106064 48442
rect 106088 48390 106102 48442
rect 106102 48390 106114 48442
rect 106114 48390 106144 48442
rect 106168 48390 106178 48442
rect 106178 48390 106224 48442
rect 105928 48388 105984 48390
rect 106008 48388 106064 48390
rect 106088 48388 106144 48390
rect 106168 48388 106224 48390
rect 106664 47898 106720 47900
rect 106744 47898 106800 47900
rect 106824 47898 106880 47900
rect 106904 47898 106960 47900
rect 106664 47846 106710 47898
rect 106710 47846 106720 47898
rect 106744 47846 106774 47898
rect 106774 47846 106786 47898
rect 106786 47846 106800 47898
rect 106824 47846 106838 47898
rect 106838 47846 106850 47898
rect 106850 47846 106880 47898
rect 106904 47846 106914 47898
rect 106914 47846 106960 47898
rect 106664 47844 106720 47846
rect 106744 47844 106800 47846
rect 106824 47844 106880 47846
rect 106904 47844 106960 47846
rect 105928 47354 105984 47356
rect 106008 47354 106064 47356
rect 106088 47354 106144 47356
rect 106168 47354 106224 47356
rect 105928 47302 105974 47354
rect 105974 47302 105984 47354
rect 106008 47302 106038 47354
rect 106038 47302 106050 47354
rect 106050 47302 106064 47354
rect 106088 47302 106102 47354
rect 106102 47302 106114 47354
rect 106114 47302 106144 47354
rect 106168 47302 106178 47354
rect 106178 47302 106224 47354
rect 105928 47300 105984 47302
rect 106008 47300 106064 47302
rect 106088 47300 106144 47302
rect 106168 47300 106224 47302
rect 106664 46810 106720 46812
rect 106744 46810 106800 46812
rect 106824 46810 106880 46812
rect 106904 46810 106960 46812
rect 106664 46758 106710 46810
rect 106710 46758 106720 46810
rect 106744 46758 106774 46810
rect 106774 46758 106786 46810
rect 106786 46758 106800 46810
rect 106824 46758 106838 46810
rect 106838 46758 106850 46810
rect 106850 46758 106880 46810
rect 106904 46758 106914 46810
rect 106914 46758 106960 46810
rect 106664 46756 106720 46758
rect 106744 46756 106800 46758
rect 106824 46756 106880 46758
rect 106904 46756 106960 46758
rect 105928 46266 105984 46268
rect 106008 46266 106064 46268
rect 106088 46266 106144 46268
rect 106168 46266 106224 46268
rect 105928 46214 105974 46266
rect 105974 46214 105984 46266
rect 106008 46214 106038 46266
rect 106038 46214 106050 46266
rect 106050 46214 106064 46266
rect 106088 46214 106102 46266
rect 106102 46214 106114 46266
rect 106114 46214 106144 46266
rect 106168 46214 106178 46266
rect 106178 46214 106224 46266
rect 105928 46212 105984 46214
rect 106008 46212 106064 46214
rect 106088 46212 106144 46214
rect 106168 46212 106224 46214
rect 106664 45722 106720 45724
rect 106744 45722 106800 45724
rect 106824 45722 106880 45724
rect 106904 45722 106960 45724
rect 106664 45670 106710 45722
rect 106710 45670 106720 45722
rect 106744 45670 106774 45722
rect 106774 45670 106786 45722
rect 106786 45670 106800 45722
rect 106824 45670 106838 45722
rect 106838 45670 106850 45722
rect 106850 45670 106880 45722
rect 106904 45670 106914 45722
rect 106914 45670 106960 45722
rect 106664 45668 106720 45670
rect 106744 45668 106800 45670
rect 106824 45668 106880 45670
rect 106904 45668 106960 45670
rect 105928 45178 105984 45180
rect 106008 45178 106064 45180
rect 106088 45178 106144 45180
rect 106168 45178 106224 45180
rect 105928 45126 105974 45178
rect 105974 45126 105984 45178
rect 106008 45126 106038 45178
rect 106038 45126 106050 45178
rect 106050 45126 106064 45178
rect 106088 45126 106102 45178
rect 106102 45126 106114 45178
rect 106114 45126 106144 45178
rect 106168 45126 106178 45178
rect 106178 45126 106224 45178
rect 105928 45124 105984 45126
rect 106008 45124 106064 45126
rect 106088 45124 106144 45126
rect 106168 45124 106224 45126
rect 106664 44634 106720 44636
rect 106744 44634 106800 44636
rect 106824 44634 106880 44636
rect 106904 44634 106960 44636
rect 106664 44582 106710 44634
rect 106710 44582 106720 44634
rect 106744 44582 106774 44634
rect 106774 44582 106786 44634
rect 106786 44582 106800 44634
rect 106824 44582 106838 44634
rect 106838 44582 106850 44634
rect 106850 44582 106880 44634
rect 106904 44582 106914 44634
rect 106914 44582 106960 44634
rect 106664 44580 106720 44582
rect 106744 44580 106800 44582
rect 106824 44580 106880 44582
rect 106904 44580 106960 44582
rect 105928 44090 105984 44092
rect 106008 44090 106064 44092
rect 106088 44090 106144 44092
rect 106168 44090 106224 44092
rect 105928 44038 105974 44090
rect 105974 44038 105984 44090
rect 106008 44038 106038 44090
rect 106038 44038 106050 44090
rect 106050 44038 106064 44090
rect 106088 44038 106102 44090
rect 106102 44038 106114 44090
rect 106114 44038 106144 44090
rect 106168 44038 106178 44090
rect 106178 44038 106224 44090
rect 105928 44036 105984 44038
rect 106008 44036 106064 44038
rect 106088 44036 106144 44038
rect 106168 44036 106224 44038
rect 106664 43546 106720 43548
rect 106744 43546 106800 43548
rect 106824 43546 106880 43548
rect 106904 43546 106960 43548
rect 106664 43494 106710 43546
rect 106710 43494 106720 43546
rect 106744 43494 106774 43546
rect 106774 43494 106786 43546
rect 106786 43494 106800 43546
rect 106824 43494 106838 43546
rect 106838 43494 106850 43546
rect 106850 43494 106880 43546
rect 106904 43494 106914 43546
rect 106914 43494 106960 43546
rect 106664 43492 106720 43494
rect 106744 43492 106800 43494
rect 106824 43492 106880 43494
rect 106904 43492 106960 43494
rect 105928 43002 105984 43004
rect 106008 43002 106064 43004
rect 106088 43002 106144 43004
rect 106168 43002 106224 43004
rect 105928 42950 105974 43002
rect 105974 42950 105984 43002
rect 106008 42950 106038 43002
rect 106038 42950 106050 43002
rect 106050 42950 106064 43002
rect 106088 42950 106102 43002
rect 106102 42950 106114 43002
rect 106114 42950 106144 43002
rect 106168 42950 106178 43002
rect 106178 42950 106224 43002
rect 105928 42948 105984 42950
rect 106008 42948 106064 42950
rect 106088 42948 106144 42950
rect 106168 42948 106224 42950
rect 106664 42458 106720 42460
rect 106744 42458 106800 42460
rect 106824 42458 106880 42460
rect 106904 42458 106960 42460
rect 106664 42406 106710 42458
rect 106710 42406 106720 42458
rect 106744 42406 106774 42458
rect 106774 42406 106786 42458
rect 106786 42406 106800 42458
rect 106824 42406 106838 42458
rect 106838 42406 106850 42458
rect 106850 42406 106880 42458
rect 106904 42406 106914 42458
rect 106914 42406 106960 42458
rect 106664 42404 106720 42406
rect 106744 42404 106800 42406
rect 106824 42404 106880 42406
rect 106904 42404 106960 42406
rect 105928 41914 105984 41916
rect 106008 41914 106064 41916
rect 106088 41914 106144 41916
rect 106168 41914 106224 41916
rect 105928 41862 105974 41914
rect 105974 41862 105984 41914
rect 106008 41862 106038 41914
rect 106038 41862 106050 41914
rect 106050 41862 106064 41914
rect 106088 41862 106102 41914
rect 106102 41862 106114 41914
rect 106114 41862 106144 41914
rect 106168 41862 106178 41914
rect 106178 41862 106224 41914
rect 105928 41860 105984 41862
rect 106008 41860 106064 41862
rect 106088 41860 106144 41862
rect 106168 41860 106224 41862
rect 106664 41370 106720 41372
rect 106744 41370 106800 41372
rect 106824 41370 106880 41372
rect 106904 41370 106960 41372
rect 106664 41318 106710 41370
rect 106710 41318 106720 41370
rect 106744 41318 106774 41370
rect 106774 41318 106786 41370
rect 106786 41318 106800 41370
rect 106824 41318 106838 41370
rect 106838 41318 106850 41370
rect 106850 41318 106880 41370
rect 106904 41318 106914 41370
rect 106914 41318 106960 41370
rect 106664 41316 106720 41318
rect 106744 41316 106800 41318
rect 106824 41316 106880 41318
rect 106904 41316 106960 41318
rect 105928 40826 105984 40828
rect 106008 40826 106064 40828
rect 106088 40826 106144 40828
rect 106168 40826 106224 40828
rect 105928 40774 105974 40826
rect 105974 40774 105984 40826
rect 106008 40774 106038 40826
rect 106038 40774 106050 40826
rect 106050 40774 106064 40826
rect 106088 40774 106102 40826
rect 106102 40774 106114 40826
rect 106114 40774 106144 40826
rect 106168 40774 106178 40826
rect 106178 40774 106224 40826
rect 105928 40772 105984 40774
rect 106008 40772 106064 40774
rect 106088 40772 106144 40774
rect 106168 40772 106224 40774
rect 106664 40282 106720 40284
rect 106744 40282 106800 40284
rect 106824 40282 106880 40284
rect 106904 40282 106960 40284
rect 106664 40230 106710 40282
rect 106710 40230 106720 40282
rect 106744 40230 106774 40282
rect 106774 40230 106786 40282
rect 106786 40230 106800 40282
rect 106824 40230 106838 40282
rect 106838 40230 106850 40282
rect 106850 40230 106880 40282
rect 106904 40230 106914 40282
rect 106914 40230 106960 40282
rect 106664 40228 106720 40230
rect 106744 40228 106800 40230
rect 106824 40228 106880 40230
rect 106904 40228 106960 40230
rect 105928 39738 105984 39740
rect 106008 39738 106064 39740
rect 106088 39738 106144 39740
rect 106168 39738 106224 39740
rect 105928 39686 105974 39738
rect 105974 39686 105984 39738
rect 106008 39686 106038 39738
rect 106038 39686 106050 39738
rect 106050 39686 106064 39738
rect 106088 39686 106102 39738
rect 106102 39686 106114 39738
rect 106114 39686 106144 39738
rect 106168 39686 106178 39738
rect 106178 39686 106224 39738
rect 105928 39684 105984 39686
rect 106008 39684 106064 39686
rect 106088 39684 106144 39686
rect 106168 39684 106224 39686
rect 106664 39194 106720 39196
rect 106744 39194 106800 39196
rect 106824 39194 106880 39196
rect 106904 39194 106960 39196
rect 106664 39142 106710 39194
rect 106710 39142 106720 39194
rect 106744 39142 106774 39194
rect 106774 39142 106786 39194
rect 106786 39142 106800 39194
rect 106824 39142 106838 39194
rect 106838 39142 106850 39194
rect 106850 39142 106880 39194
rect 106904 39142 106914 39194
rect 106914 39142 106960 39194
rect 106664 39140 106720 39142
rect 106744 39140 106800 39142
rect 106824 39140 106880 39142
rect 106904 39140 106960 39142
rect 105928 38650 105984 38652
rect 106008 38650 106064 38652
rect 106088 38650 106144 38652
rect 106168 38650 106224 38652
rect 105928 38598 105974 38650
rect 105974 38598 105984 38650
rect 106008 38598 106038 38650
rect 106038 38598 106050 38650
rect 106050 38598 106064 38650
rect 106088 38598 106102 38650
rect 106102 38598 106114 38650
rect 106114 38598 106144 38650
rect 106168 38598 106178 38650
rect 106178 38598 106224 38650
rect 105928 38596 105984 38598
rect 106008 38596 106064 38598
rect 106088 38596 106144 38598
rect 106168 38596 106224 38598
rect 106664 38106 106720 38108
rect 106744 38106 106800 38108
rect 106824 38106 106880 38108
rect 106904 38106 106960 38108
rect 106664 38054 106710 38106
rect 106710 38054 106720 38106
rect 106744 38054 106774 38106
rect 106774 38054 106786 38106
rect 106786 38054 106800 38106
rect 106824 38054 106838 38106
rect 106838 38054 106850 38106
rect 106850 38054 106880 38106
rect 106904 38054 106914 38106
rect 106914 38054 106960 38106
rect 106664 38052 106720 38054
rect 106744 38052 106800 38054
rect 106824 38052 106880 38054
rect 106904 38052 106960 38054
rect 105928 37562 105984 37564
rect 106008 37562 106064 37564
rect 106088 37562 106144 37564
rect 106168 37562 106224 37564
rect 105928 37510 105974 37562
rect 105974 37510 105984 37562
rect 106008 37510 106038 37562
rect 106038 37510 106050 37562
rect 106050 37510 106064 37562
rect 106088 37510 106102 37562
rect 106102 37510 106114 37562
rect 106114 37510 106144 37562
rect 106168 37510 106178 37562
rect 106178 37510 106224 37562
rect 105928 37508 105984 37510
rect 106008 37508 106064 37510
rect 106088 37508 106144 37510
rect 106168 37508 106224 37510
rect 106664 37018 106720 37020
rect 106744 37018 106800 37020
rect 106824 37018 106880 37020
rect 106904 37018 106960 37020
rect 106664 36966 106710 37018
rect 106710 36966 106720 37018
rect 106744 36966 106774 37018
rect 106774 36966 106786 37018
rect 106786 36966 106800 37018
rect 106824 36966 106838 37018
rect 106838 36966 106850 37018
rect 106850 36966 106880 37018
rect 106904 36966 106914 37018
rect 106914 36966 106960 37018
rect 106664 36964 106720 36966
rect 106744 36964 106800 36966
rect 106824 36964 106880 36966
rect 106904 36964 106960 36966
rect 105928 36474 105984 36476
rect 106008 36474 106064 36476
rect 106088 36474 106144 36476
rect 106168 36474 106224 36476
rect 105928 36422 105974 36474
rect 105974 36422 105984 36474
rect 106008 36422 106038 36474
rect 106038 36422 106050 36474
rect 106050 36422 106064 36474
rect 106088 36422 106102 36474
rect 106102 36422 106114 36474
rect 106114 36422 106144 36474
rect 106168 36422 106178 36474
rect 106178 36422 106224 36474
rect 105928 36420 105984 36422
rect 106008 36420 106064 36422
rect 106088 36420 106144 36422
rect 106168 36420 106224 36422
rect 106664 35930 106720 35932
rect 106744 35930 106800 35932
rect 106824 35930 106880 35932
rect 106904 35930 106960 35932
rect 106664 35878 106710 35930
rect 106710 35878 106720 35930
rect 106744 35878 106774 35930
rect 106774 35878 106786 35930
rect 106786 35878 106800 35930
rect 106824 35878 106838 35930
rect 106838 35878 106850 35930
rect 106850 35878 106880 35930
rect 106904 35878 106914 35930
rect 106914 35878 106960 35930
rect 106664 35876 106720 35878
rect 106744 35876 106800 35878
rect 106824 35876 106880 35878
rect 106904 35876 106960 35878
rect 105928 35386 105984 35388
rect 106008 35386 106064 35388
rect 106088 35386 106144 35388
rect 106168 35386 106224 35388
rect 105928 35334 105974 35386
rect 105974 35334 105984 35386
rect 106008 35334 106038 35386
rect 106038 35334 106050 35386
rect 106050 35334 106064 35386
rect 106088 35334 106102 35386
rect 106102 35334 106114 35386
rect 106114 35334 106144 35386
rect 106168 35334 106178 35386
rect 106178 35334 106224 35386
rect 105928 35332 105984 35334
rect 106008 35332 106064 35334
rect 106088 35332 106144 35334
rect 106168 35332 106224 35334
rect 106664 34842 106720 34844
rect 106744 34842 106800 34844
rect 106824 34842 106880 34844
rect 106904 34842 106960 34844
rect 106664 34790 106710 34842
rect 106710 34790 106720 34842
rect 106744 34790 106774 34842
rect 106774 34790 106786 34842
rect 106786 34790 106800 34842
rect 106824 34790 106838 34842
rect 106838 34790 106850 34842
rect 106850 34790 106880 34842
rect 106904 34790 106914 34842
rect 106914 34790 106960 34842
rect 106664 34788 106720 34790
rect 106744 34788 106800 34790
rect 106824 34788 106880 34790
rect 106904 34788 106960 34790
rect 105928 34298 105984 34300
rect 106008 34298 106064 34300
rect 106088 34298 106144 34300
rect 106168 34298 106224 34300
rect 105928 34246 105974 34298
rect 105974 34246 105984 34298
rect 106008 34246 106038 34298
rect 106038 34246 106050 34298
rect 106050 34246 106064 34298
rect 106088 34246 106102 34298
rect 106102 34246 106114 34298
rect 106114 34246 106144 34298
rect 106168 34246 106178 34298
rect 106178 34246 106224 34298
rect 105928 34244 105984 34246
rect 106008 34244 106064 34246
rect 106088 34244 106144 34246
rect 106168 34244 106224 34246
rect 106664 33754 106720 33756
rect 106744 33754 106800 33756
rect 106824 33754 106880 33756
rect 106904 33754 106960 33756
rect 106664 33702 106710 33754
rect 106710 33702 106720 33754
rect 106744 33702 106774 33754
rect 106774 33702 106786 33754
rect 106786 33702 106800 33754
rect 106824 33702 106838 33754
rect 106838 33702 106850 33754
rect 106850 33702 106880 33754
rect 106904 33702 106914 33754
rect 106914 33702 106960 33754
rect 106664 33700 106720 33702
rect 106744 33700 106800 33702
rect 106824 33700 106880 33702
rect 106904 33700 106960 33702
rect 105928 33210 105984 33212
rect 106008 33210 106064 33212
rect 106088 33210 106144 33212
rect 106168 33210 106224 33212
rect 105928 33158 105974 33210
rect 105974 33158 105984 33210
rect 106008 33158 106038 33210
rect 106038 33158 106050 33210
rect 106050 33158 106064 33210
rect 106088 33158 106102 33210
rect 106102 33158 106114 33210
rect 106114 33158 106144 33210
rect 106168 33158 106178 33210
rect 106178 33158 106224 33210
rect 105928 33156 105984 33158
rect 106008 33156 106064 33158
rect 106088 33156 106144 33158
rect 106168 33156 106224 33158
rect 106664 32666 106720 32668
rect 106744 32666 106800 32668
rect 106824 32666 106880 32668
rect 106904 32666 106960 32668
rect 106664 32614 106710 32666
rect 106710 32614 106720 32666
rect 106744 32614 106774 32666
rect 106774 32614 106786 32666
rect 106786 32614 106800 32666
rect 106824 32614 106838 32666
rect 106838 32614 106850 32666
rect 106850 32614 106880 32666
rect 106904 32614 106914 32666
rect 106914 32614 106960 32666
rect 106664 32612 106720 32614
rect 106744 32612 106800 32614
rect 106824 32612 106880 32614
rect 106904 32612 106960 32614
rect 105928 32122 105984 32124
rect 106008 32122 106064 32124
rect 106088 32122 106144 32124
rect 106168 32122 106224 32124
rect 105928 32070 105974 32122
rect 105974 32070 105984 32122
rect 106008 32070 106038 32122
rect 106038 32070 106050 32122
rect 106050 32070 106064 32122
rect 106088 32070 106102 32122
rect 106102 32070 106114 32122
rect 106114 32070 106144 32122
rect 106168 32070 106178 32122
rect 106178 32070 106224 32122
rect 105928 32068 105984 32070
rect 106008 32068 106064 32070
rect 106088 32068 106144 32070
rect 106168 32068 106224 32070
rect 106664 31578 106720 31580
rect 106744 31578 106800 31580
rect 106824 31578 106880 31580
rect 106904 31578 106960 31580
rect 106664 31526 106710 31578
rect 106710 31526 106720 31578
rect 106744 31526 106774 31578
rect 106774 31526 106786 31578
rect 106786 31526 106800 31578
rect 106824 31526 106838 31578
rect 106838 31526 106850 31578
rect 106850 31526 106880 31578
rect 106904 31526 106914 31578
rect 106914 31526 106960 31578
rect 106664 31524 106720 31526
rect 106744 31524 106800 31526
rect 106824 31524 106880 31526
rect 106904 31524 106960 31526
rect 105928 31034 105984 31036
rect 106008 31034 106064 31036
rect 106088 31034 106144 31036
rect 106168 31034 106224 31036
rect 105928 30982 105974 31034
rect 105974 30982 105984 31034
rect 106008 30982 106038 31034
rect 106038 30982 106050 31034
rect 106050 30982 106064 31034
rect 106088 30982 106102 31034
rect 106102 30982 106114 31034
rect 106114 30982 106144 31034
rect 106168 30982 106178 31034
rect 106178 30982 106224 31034
rect 105928 30980 105984 30982
rect 106008 30980 106064 30982
rect 106088 30980 106144 30982
rect 106168 30980 106224 30982
rect 106664 30490 106720 30492
rect 106744 30490 106800 30492
rect 106824 30490 106880 30492
rect 106904 30490 106960 30492
rect 106664 30438 106710 30490
rect 106710 30438 106720 30490
rect 106744 30438 106774 30490
rect 106774 30438 106786 30490
rect 106786 30438 106800 30490
rect 106824 30438 106838 30490
rect 106838 30438 106850 30490
rect 106850 30438 106880 30490
rect 106904 30438 106914 30490
rect 106914 30438 106960 30490
rect 106664 30436 106720 30438
rect 106744 30436 106800 30438
rect 106824 30436 106880 30438
rect 106904 30436 106960 30438
rect 105928 29946 105984 29948
rect 106008 29946 106064 29948
rect 106088 29946 106144 29948
rect 106168 29946 106224 29948
rect 105928 29894 105974 29946
rect 105974 29894 105984 29946
rect 106008 29894 106038 29946
rect 106038 29894 106050 29946
rect 106050 29894 106064 29946
rect 106088 29894 106102 29946
rect 106102 29894 106114 29946
rect 106114 29894 106144 29946
rect 106168 29894 106178 29946
rect 106178 29894 106224 29946
rect 105928 29892 105984 29894
rect 106008 29892 106064 29894
rect 106088 29892 106144 29894
rect 106168 29892 106224 29894
rect 106664 29402 106720 29404
rect 106744 29402 106800 29404
rect 106824 29402 106880 29404
rect 106904 29402 106960 29404
rect 106664 29350 106710 29402
rect 106710 29350 106720 29402
rect 106744 29350 106774 29402
rect 106774 29350 106786 29402
rect 106786 29350 106800 29402
rect 106824 29350 106838 29402
rect 106838 29350 106850 29402
rect 106850 29350 106880 29402
rect 106904 29350 106914 29402
rect 106914 29350 106960 29402
rect 106664 29348 106720 29350
rect 106744 29348 106800 29350
rect 106824 29348 106880 29350
rect 106904 29348 106960 29350
rect 105928 28858 105984 28860
rect 106008 28858 106064 28860
rect 106088 28858 106144 28860
rect 106168 28858 106224 28860
rect 105928 28806 105974 28858
rect 105974 28806 105984 28858
rect 106008 28806 106038 28858
rect 106038 28806 106050 28858
rect 106050 28806 106064 28858
rect 106088 28806 106102 28858
rect 106102 28806 106114 28858
rect 106114 28806 106144 28858
rect 106168 28806 106178 28858
rect 106178 28806 106224 28858
rect 105928 28804 105984 28806
rect 106008 28804 106064 28806
rect 106088 28804 106144 28806
rect 106168 28804 106224 28806
rect 106664 28314 106720 28316
rect 106744 28314 106800 28316
rect 106824 28314 106880 28316
rect 106904 28314 106960 28316
rect 106664 28262 106710 28314
rect 106710 28262 106720 28314
rect 106744 28262 106774 28314
rect 106774 28262 106786 28314
rect 106786 28262 106800 28314
rect 106824 28262 106838 28314
rect 106838 28262 106850 28314
rect 106850 28262 106880 28314
rect 106904 28262 106914 28314
rect 106914 28262 106960 28314
rect 106664 28260 106720 28262
rect 106744 28260 106800 28262
rect 106824 28260 106880 28262
rect 106904 28260 106960 28262
rect 105928 27770 105984 27772
rect 106008 27770 106064 27772
rect 106088 27770 106144 27772
rect 106168 27770 106224 27772
rect 105928 27718 105974 27770
rect 105974 27718 105984 27770
rect 106008 27718 106038 27770
rect 106038 27718 106050 27770
rect 106050 27718 106064 27770
rect 106088 27718 106102 27770
rect 106102 27718 106114 27770
rect 106114 27718 106144 27770
rect 106168 27718 106178 27770
rect 106178 27718 106224 27770
rect 105928 27716 105984 27718
rect 106008 27716 106064 27718
rect 106088 27716 106144 27718
rect 106168 27716 106224 27718
rect 106664 27226 106720 27228
rect 106744 27226 106800 27228
rect 106824 27226 106880 27228
rect 106904 27226 106960 27228
rect 106664 27174 106710 27226
rect 106710 27174 106720 27226
rect 106744 27174 106774 27226
rect 106774 27174 106786 27226
rect 106786 27174 106800 27226
rect 106824 27174 106838 27226
rect 106838 27174 106850 27226
rect 106850 27174 106880 27226
rect 106904 27174 106914 27226
rect 106914 27174 106960 27226
rect 106664 27172 106720 27174
rect 106744 27172 106800 27174
rect 106824 27172 106880 27174
rect 106904 27172 106960 27174
rect 105928 26682 105984 26684
rect 106008 26682 106064 26684
rect 106088 26682 106144 26684
rect 106168 26682 106224 26684
rect 105928 26630 105974 26682
rect 105974 26630 105984 26682
rect 106008 26630 106038 26682
rect 106038 26630 106050 26682
rect 106050 26630 106064 26682
rect 106088 26630 106102 26682
rect 106102 26630 106114 26682
rect 106114 26630 106144 26682
rect 106168 26630 106178 26682
rect 106178 26630 106224 26682
rect 105928 26628 105984 26630
rect 106008 26628 106064 26630
rect 106088 26628 106144 26630
rect 106168 26628 106224 26630
rect 106664 26138 106720 26140
rect 106744 26138 106800 26140
rect 106824 26138 106880 26140
rect 106904 26138 106960 26140
rect 106664 26086 106710 26138
rect 106710 26086 106720 26138
rect 106744 26086 106774 26138
rect 106774 26086 106786 26138
rect 106786 26086 106800 26138
rect 106824 26086 106838 26138
rect 106838 26086 106850 26138
rect 106850 26086 106880 26138
rect 106904 26086 106914 26138
rect 106914 26086 106960 26138
rect 106664 26084 106720 26086
rect 106744 26084 106800 26086
rect 106824 26084 106880 26086
rect 106904 26084 106960 26086
rect 105928 25594 105984 25596
rect 106008 25594 106064 25596
rect 106088 25594 106144 25596
rect 106168 25594 106224 25596
rect 105928 25542 105974 25594
rect 105974 25542 105984 25594
rect 106008 25542 106038 25594
rect 106038 25542 106050 25594
rect 106050 25542 106064 25594
rect 106088 25542 106102 25594
rect 106102 25542 106114 25594
rect 106114 25542 106144 25594
rect 106168 25542 106178 25594
rect 106178 25542 106224 25594
rect 105928 25540 105984 25542
rect 106008 25540 106064 25542
rect 106088 25540 106144 25542
rect 106168 25540 106224 25542
rect 106664 25050 106720 25052
rect 106744 25050 106800 25052
rect 106824 25050 106880 25052
rect 106904 25050 106960 25052
rect 106664 24998 106710 25050
rect 106710 24998 106720 25050
rect 106744 24998 106774 25050
rect 106774 24998 106786 25050
rect 106786 24998 106800 25050
rect 106824 24998 106838 25050
rect 106838 24998 106850 25050
rect 106850 24998 106880 25050
rect 106904 24998 106914 25050
rect 106914 24998 106960 25050
rect 106664 24996 106720 24998
rect 106744 24996 106800 24998
rect 106824 24996 106880 24998
rect 106904 24996 106960 24998
rect 105928 24506 105984 24508
rect 106008 24506 106064 24508
rect 106088 24506 106144 24508
rect 106168 24506 106224 24508
rect 105928 24454 105974 24506
rect 105974 24454 105984 24506
rect 106008 24454 106038 24506
rect 106038 24454 106050 24506
rect 106050 24454 106064 24506
rect 106088 24454 106102 24506
rect 106102 24454 106114 24506
rect 106114 24454 106144 24506
rect 106168 24454 106178 24506
rect 106178 24454 106224 24506
rect 105928 24452 105984 24454
rect 106008 24452 106064 24454
rect 106088 24452 106144 24454
rect 106168 24452 106224 24454
rect 106664 23962 106720 23964
rect 106744 23962 106800 23964
rect 106824 23962 106880 23964
rect 106904 23962 106960 23964
rect 106664 23910 106710 23962
rect 106710 23910 106720 23962
rect 106744 23910 106774 23962
rect 106774 23910 106786 23962
rect 106786 23910 106800 23962
rect 106824 23910 106838 23962
rect 106838 23910 106850 23962
rect 106850 23910 106880 23962
rect 106904 23910 106914 23962
rect 106914 23910 106960 23962
rect 106664 23908 106720 23910
rect 106744 23908 106800 23910
rect 106824 23908 106880 23910
rect 106904 23908 106960 23910
rect 105928 23418 105984 23420
rect 106008 23418 106064 23420
rect 106088 23418 106144 23420
rect 106168 23418 106224 23420
rect 105928 23366 105974 23418
rect 105974 23366 105984 23418
rect 106008 23366 106038 23418
rect 106038 23366 106050 23418
rect 106050 23366 106064 23418
rect 106088 23366 106102 23418
rect 106102 23366 106114 23418
rect 106114 23366 106144 23418
rect 106168 23366 106178 23418
rect 106178 23366 106224 23418
rect 105928 23364 105984 23366
rect 106008 23364 106064 23366
rect 106088 23364 106144 23366
rect 106168 23364 106224 23366
rect 106664 22874 106720 22876
rect 106744 22874 106800 22876
rect 106824 22874 106880 22876
rect 106904 22874 106960 22876
rect 106664 22822 106710 22874
rect 106710 22822 106720 22874
rect 106744 22822 106774 22874
rect 106774 22822 106786 22874
rect 106786 22822 106800 22874
rect 106824 22822 106838 22874
rect 106838 22822 106850 22874
rect 106850 22822 106880 22874
rect 106904 22822 106914 22874
rect 106914 22822 106960 22874
rect 106664 22820 106720 22822
rect 106744 22820 106800 22822
rect 106824 22820 106880 22822
rect 106904 22820 106960 22822
rect 105928 22330 105984 22332
rect 106008 22330 106064 22332
rect 106088 22330 106144 22332
rect 106168 22330 106224 22332
rect 105928 22278 105974 22330
rect 105974 22278 105984 22330
rect 106008 22278 106038 22330
rect 106038 22278 106050 22330
rect 106050 22278 106064 22330
rect 106088 22278 106102 22330
rect 106102 22278 106114 22330
rect 106114 22278 106144 22330
rect 106168 22278 106178 22330
rect 106178 22278 106224 22330
rect 105928 22276 105984 22278
rect 106008 22276 106064 22278
rect 106088 22276 106144 22278
rect 106168 22276 106224 22278
rect 106664 21786 106720 21788
rect 106744 21786 106800 21788
rect 106824 21786 106880 21788
rect 106904 21786 106960 21788
rect 106664 21734 106710 21786
rect 106710 21734 106720 21786
rect 106744 21734 106774 21786
rect 106774 21734 106786 21786
rect 106786 21734 106800 21786
rect 106824 21734 106838 21786
rect 106838 21734 106850 21786
rect 106850 21734 106880 21786
rect 106904 21734 106914 21786
rect 106914 21734 106960 21786
rect 106664 21732 106720 21734
rect 106744 21732 106800 21734
rect 106824 21732 106880 21734
rect 106904 21732 106960 21734
rect 105928 21242 105984 21244
rect 106008 21242 106064 21244
rect 106088 21242 106144 21244
rect 106168 21242 106224 21244
rect 105928 21190 105974 21242
rect 105974 21190 105984 21242
rect 106008 21190 106038 21242
rect 106038 21190 106050 21242
rect 106050 21190 106064 21242
rect 106088 21190 106102 21242
rect 106102 21190 106114 21242
rect 106114 21190 106144 21242
rect 106168 21190 106178 21242
rect 106178 21190 106224 21242
rect 105928 21188 105984 21190
rect 106008 21188 106064 21190
rect 106088 21188 106144 21190
rect 106168 21188 106224 21190
rect 106664 20698 106720 20700
rect 106744 20698 106800 20700
rect 106824 20698 106880 20700
rect 106904 20698 106960 20700
rect 106664 20646 106710 20698
rect 106710 20646 106720 20698
rect 106744 20646 106774 20698
rect 106774 20646 106786 20698
rect 106786 20646 106800 20698
rect 106824 20646 106838 20698
rect 106838 20646 106850 20698
rect 106850 20646 106880 20698
rect 106904 20646 106914 20698
rect 106914 20646 106960 20698
rect 106664 20644 106720 20646
rect 106744 20644 106800 20646
rect 106824 20644 106880 20646
rect 106904 20644 106960 20646
rect 105928 20154 105984 20156
rect 106008 20154 106064 20156
rect 106088 20154 106144 20156
rect 106168 20154 106224 20156
rect 105928 20102 105974 20154
rect 105974 20102 105984 20154
rect 106008 20102 106038 20154
rect 106038 20102 106050 20154
rect 106050 20102 106064 20154
rect 106088 20102 106102 20154
rect 106102 20102 106114 20154
rect 106114 20102 106144 20154
rect 106168 20102 106178 20154
rect 106178 20102 106224 20154
rect 105928 20100 105984 20102
rect 106008 20100 106064 20102
rect 106088 20100 106144 20102
rect 106168 20100 106224 20102
rect 106664 19610 106720 19612
rect 106744 19610 106800 19612
rect 106824 19610 106880 19612
rect 106904 19610 106960 19612
rect 106664 19558 106710 19610
rect 106710 19558 106720 19610
rect 106744 19558 106774 19610
rect 106774 19558 106786 19610
rect 106786 19558 106800 19610
rect 106824 19558 106838 19610
rect 106838 19558 106850 19610
rect 106850 19558 106880 19610
rect 106904 19558 106914 19610
rect 106914 19558 106960 19610
rect 106664 19556 106720 19558
rect 106744 19556 106800 19558
rect 106824 19556 106880 19558
rect 106904 19556 106960 19558
rect 105928 19066 105984 19068
rect 106008 19066 106064 19068
rect 106088 19066 106144 19068
rect 106168 19066 106224 19068
rect 105928 19014 105974 19066
rect 105974 19014 105984 19066
rect 106008 19014 106038 19066
rect 106038 19014 106050 19066
rect 106050 19014 106064 19066
rect 106088 19014 106102 19066
rect 106102 19014 106114 19066
rect 106114 19014 106144 19066
rect 106168 19014 106178 19066
rect 106178 19014 106224 19066
rect 105928 19012 105984 19014
rect 106008 19012 106064 19014
rect 106088 19012 106144 19014
rect 106168 19012 106224 19014
rect 106664 18522 106720 18524
rect 106744 18522 106800 18524
rect 106824 18522 106880 18524
rect 106904 18522 106960 18524
rect 106664 18470 106710 18522
rect 106710 18470 106720 18522
rect 106744 18470 106774 18522
rect 106774 18470 106786 18522
rect 106786 18470 106800 18522
rect 106824 18470 106838 18522
rect 106838 18470 106850 18522
rect 106850 18470 106880 18522
rect 106904 18470 106914 18522
rect 106914 18470 106960 18522
rect 106664 18468 106720 18470
rect 106744 18468 106800 18470
rect 106824 18468 106880 18470
rect 106904 18468 106960 18470
rect 105928 17978 105984 17980
rect 106008 17978 106064 17980
rect 106088 17978 106144 17980
rect 106168 17978 106224 17980
rect 105928 17926 105974 17978
rect 105974 17926 105984 17978
rect 106008 17926 106038 17978
rect 106038 17926 106050 17978
rect 106050 17926 106064 17978
rect 106088 17926 106102 17978
rect 106102 17926 106114 17978
rect 106114 17926 106144 17978
rect 106168 17926 106178 17978
rect 106178 17926 106224 17978
rect 105928 17924 105984 17926
rect 106008 17924 106064 17926
rect 106088 17924 106144 17926
rect 106168 17924 106224 17926
rect 106664 17434 106720 17436
rect 106744 17434 106800 17436
rect 106824 17434 106880 17436
rect 106904 17434 106960 17436
rect 106664 17382 106710 17434
rect 106710 17382 106720 17434
rect 106744 17382 106774 17434
rect 106774 17382 106786 17434
rect 106786 17382 106800 17434
rect 106824 17382 106838 17434
rect 106838 17382 106850 17434
rect 106850 17382 106880 17434
rect 106904 17382 106914 17434
rect 106914 17382 106960 17434
rect 106664 17380 106720 17382
rect 106744 17380 106800 17382
rect 106824 17380 106880 17382
rect 106904 17380 106960 17382
rect 105928 16890 105984 16892
rect 106008 16890 106064 16892
rect 106088 16890 106144 16892
rect 106168 16890 106224 16892
rect 105928 16838 105974 16890
rect 105974 16838 105984 16890
rect 106008 16838 106038 16890
rect 106038 16838 106050 16890
rect 106050 16838 106064 16890
rect 106088 16838 106102 16890
rect 106102 16838 106114 16890
rect 106114 16838 106144 16890
rect 106168 16838 106178 16890
rect 106178 16838 106224 16890
rect 105928 16836 105984 16838
rect 106008 16836 106064 16838
rect 106088 16836 106144 16838
rect 106168 16836 106224 16838
rect 106664 16346 106720 16348
rect 106744 16346 106800 16348
rect 106824 16346 106880 16348
rect 106904 16346 106960 16348
rect 106664 16294 106710 16346
rect 106710 16294 106720 16346
rect 106744 16294 106774 16346
rect 106774 16294 106786 16346
rect 106786 16294 106800 16346
rect 106824 16294 106838 16346
rect 106838 16294 106850 16346
rect 106850 16294 106880 16346
rect 106904 16294 106914 16346
rect 106914 16294 106960 16346
rect 106664 16292 106720 16294
rect 106744 16292 106800 16294
rect 106824 16292 106880 16294
rect 106904 16292 106960 16294
rect 105928 15802 105984 15804
rect 106008 15802 106064 15804
rect 106088 15802 106144 15804
rect 106168 15802 106224 15804
rect 105928 15750 105974 15802
rect 105974 15750 105984 15802
rect 106008 15750 106038 15802
rect 106038 15750 106050 15802
rect 106050 15750 106064 15802
rect 106088 15750 106102 15802
rect 106102 15750 106114 15802
rect 106114 15750 106144 15802
rect 106168 15750 106178 15802
rect 106178 15750 106224 15802
rect 105928 15748 105984 15750
rect 106008 15748 106064 15750
rect 106088 15748 106144 15750
rect 106168 15748 106224 15750
rect 106664 15258 106720 15260
rect 106744 15258 106800 15260
rect 106824 15258 106880 15260
rect 106904 15258 106960 15260
rect 106664 15206 106710 15258
rect 106710 15206 106720 15258
rect 106744 15206 106774 15258
rect 106774 15206 106786 15258
rect 106786 15206 106800 15258
rect 106824 15206 106838 15258
rect 106838 15206 106850 15258
rect 106850 15206 106880 15258
rect 106904 15206 106914 15258
rect 106914 15206 106960 15258
rect 106664 15204 106720 15206
rect 106744 15204 106800 15206
rect 106824 15204 106880 15206
rect 106904 15204 106960 15206
rect 105928 14714 105984 14716
rect 106008 14714 106064 14716
rect 106088 14714 106144 14716
rect 106168 14714 106224 14716
rect 105928 14662 105974 14714
rect 105974 14662 105984 14714
rect 106008 14662 106038 14714
rect 106038 14662 106050 14714
rect 106050 14662 106064 14714
rect 106088 14662 106102 14714
rect 106102 14662 106114 14714
rect 106114 14662 106144 14714
rect 106168 14662 106178 14714
rect 106178 14662 106224 14714
rect 105928 14660 105984 14662
rect 106008 14660 106064 14662
rect 106088 14660 106144 14662
rect 106168 14660 106224 14662
rect 106664 14170 106720 14172
rect 106744 14170 106800 14172
rect 106824 14170 106880 14172
rect 106904 14170 106960 14172
rect 106664 14118 106710 14170
rect 106710 14118 106720 14170
rect 106744 14118 106774 14170
rect 106774 14118 106786 14170
rect 106786 14118 106800 14170
rect 106824 14118 106838 14170
rect 106838 14118 106850 14170
rect 106850 14118 106880 14170
rect 106904 14118 106914 14170
rect 106914 14118 106960 14170
rect 106664 14116 106720 14118
rect 106744 14116 106800 14118
rect 106824 14116 106880 14118
rect 106904 14116 106960 14118
rect 105928 13626 105984 13628
rect 106008 13626 106064 13628
rect 106088 13626 106144 13628
rect 106168 13626 106224 13628
rect 105928 13574 105974 13626
rect 105974 13574 105984 13626
rect 106008 13574 106038 13626
rect 106038 13574 106050 13626
rect 106050 13574 106064 13626
rect 106088 13574 106102 13626
rect 106102 13574 106114 13626
rect 106114 13574 106144 13626
rect 106168 13574 106178 13626
rect 106178 13574 106224 13626
rect 105928 13572 105984 13574
rect 106008 13572 106064 13574
rect 106088 13572 106144 13574
rect 106168 13572 106224 13574
rect 106664 13082 106720 13084
rect 106744 13082 106800 13084
rect 106824 13082 106880 13084
rect 106904 13082 106960 13084
rect 106664 13030 106710 13082
rect 106710 13030 106720 13082
rect 106744 13030 106774 13082
rect 106774 13030 106786 13082
rect 106786 13030 106800 13082
rect 106824 13030 106838 13082
rect 106838 13030 106850 13082
rect 106850 13030 106880 13082
rect 106904 13030 106914 13082
rect 106914 13030 106960 13082
rect 106664 13028 106720 13030
rect 106744 13028 106800 13030
rect 106824 13028 106880 13030
rect 106904 13028 106960 13030
rect 105928 12538 105984 12540
rect 106008 12538 106064 12540
rect 106088 12538 106144 12540
rect 106168 12538 106224 12540
rect 105928 12486 105974 12538
rect 105974 12486 105984 12538
rect 106008 12486 106038 12538
rect 106038 12486 106050 12538
rect 106050 12486 106064 12538
rect 106088 12486 106102 12538
rect 106102 12486 106114 12538
rect 106114 12486 106144 12538
rect 106168 12486 106178 12538
rect 106178 12486 106224 12538
rect 105928 12484 105984 12486
rect 106008 12484 106064 12486
rect 106088 12484 106144 12486
rect 106168 12484 106224 12486
rect 106664 11994 106720 11996
rect 106744 11994 106800 11996
rect 106824 11994 106880 11996
rect 106904 11994 106960 11996
rect 106664 11942 106710 11994
rect 106710 11942 106720 11994
rect 106744 11942 106774 11994
rect 106774 11942 106786 11994
rect 106786 11942 106800 11994
rect 106824 11942 106838 11994
rect 106838 11942 106850 11994
rect 106850 11942 106880 11994
rect 106904 11942 106914 11994
rect 106914 11942 106960 11994
rect 106664 11940 106720 11942
rect 106744 11940 106800 11942
rect 106824 11940 106880 11942
rect 106904 11940 106960 11942
rect 105928 11450 105984 11452
rect 106008 11450 106064 11452
rect 106088 11450 106144 11452
rect 106168 11450 106224 11452
rect 105928 11398 105974 11450
rect 105974 11398 105984 11450
rect 106008 11398 106038 11450
rect 106038 11398 106050 11450
rect 106050 11398 106064 11450
rect 106088 11398 106102 11450
rect 106102 11398 106114 11450
rect 106114 11398 106144 11450
rect 106168 11398 106178 11450
rect 106178 11398 106224 11450
rect 105928 11396 105984 11398
rect 106008 11396 106064 11398
rect 106088 11396 106144 11398
rect 106168 11396 106224 11398
rect 106664 10906 106720 10908
rect 106744 10906 106800 10908
rect 106824 10906 106880 10908
rect 106904 10906 106960 10908
rect 106664 10854 106710 10906
rect 106710 10854 106720 10906
rect 106744 10854 106774 10906
rect 106774 10854 106786 10906
rect 106786 10854 106800 10906
rect 106824 10854 106838 10906
rect 106838 10854 106850 10906
rect 106850 10854 106880 10906
rect 106904 10854 106914 10906
rect 106914 10854 106960 10906
rect 106664 10852 106720 10854
rect 106744 10852 106800 10854
rect 106824 10852 106880 10854
rect 106904 10852 106960 10854
rect 105928 10362 105984 10364
rect 106008 10362 106064 10364
rect 106088 10362 106144 10364
rect 106168 10362 106224 10364
rect 105928 10310 105974 10362
rect 105974 10310 105984 10362
rect 106008 10310 106038 10362
rect 106038 10310 106050 10362
rect 106050 10310 106064 10362
rect 106088 10310 106102 10362
rect 106102 10310 106114 10362
rect 106114 10310 106144 10362
rect 106168 10310 106178 10362
rect 106178 10310 106224 10362
rect 105928 10308 105984 10310
rect 106008 10308 106064 10310
rect 106088 10308 106144 10310
rect 106168 10308 106224 10310
rect 106664 9818 106720 9820
rect 106744 9818 106800 9820
rect 106824 9818 106880 9820
rect 106904 9818 106960 9820
rect 106664 9766 106710 9818
rect 106710 9766 106720 9818
rect 106744 9766 106774 9818
rect 106774 9766 106786 9818
rect 106786 9766 106800 9818
rect 106824 9766 106838 9818
rect 106838 9766 106850 9818
rect 106850 9766 106880 9818
rect 106904 9766 106914 9818
rect 106914 9766 106960 9818
rect 106664 9764 106720 9766
rect 106744 9764 106800 9766
rect 106824 9764 106880 9766
rect 106904 9764 106960 9766
rect 105928 9274 105984 9276
rect 106008 9274 106064 9276
rect 106088 9274 106144 9276
rect 106168 9274 106224 9276
rect 105928 9222 105974 9274
rect 105974 9222 105984 9274
rect 106008 9222 106038 9274
rect 106038 9222 106050 9274
rect 106050 9222 106064 9274
rect 106088 9222 106102 9274
rect 106102 9222 106114 9274
rect 106114 9222 106144 9274
rect 106168 9222 106178 9274
rect 106178 9222 106224 9274
rect 105928 9220 105984 9222
rect 106008 9220 106064 9222
rect 106088 9220 106144 9222
rect 106168 9220 106224 9222
rect 106664 8730 106720 8732
rect 106744 8730 106800 8732
rect 106824 8730 106880 8732
rect 106904 8730 106960 8732
rect 106664 8678 106710 8730
rect 106710 8678 106720 8730
rect 106744 8678 106774 8730
rect 106774 8678 106786 8730
rect 106786 8678 106800 8730
rect 106824 8678 106838 8730
rect 106838 8678 106850 8730
rect 106850 8678 106880 8730
rect 106904 8678 106914 8730
rect 106914 8678 106960 8730
rect 106664 8676 106720 8678
rect 106744 8676 106800 8678
rect 106824 8676 106880 8678
rect 106904 8676 106960 8678
rect 105928 8186 105984 8188
rect 106008 8186 106064 8188
rect 106088 8186 106144 8188
rect 106168 8186 106224 8188
rect 105928 8134 105974 8186
rect 105974 8134 105984 8186
rect 106008 8134 106038 8186
rect 106038 8134 106050 8186
rect 106050 8134 106064 8186
rect 106088 8134 106102 8186
rect 106102 8134 106114 8186
rect 106114 8134 106144 8186
rect 106168 8134 106178 8186
rect 106178 8134 106224 8186
rect 105928 8132 105984 8134
rect 106008 8132 106064 8134
rect 106088 8132 106144 8134
rect 106168 8132 106224 8134
rect 97040 7642 97096 7644
rect 97120 7642 97176 7644
rect 97200 7642 97256 7644
rect 97280 7642 97336 7644
rect 97040 7590 97086 7642
rect 97086 7590 97096 7642
rect 97120 7590 97150 7642
rect 97150 7590 97162 7642
rect 97162 7590 97176 7642
rect 97200 7590 97214 7642
rect 97214 7590 97226 7642
rect 97226 7590 97256 7642
rect 97280 7590 97290 7642
rect 97290 7590 97336 7642
rect 97040 7588 97096 7590
rect 97120 7588 97176 7590
rect 97200 7588 97256 7590
rect 97280 7588 97336 7590
rect 106664 7642 106720 7644
rect 106744 7642 106800 7644
rect 106824 7642 106880 7644
rect 106904 7642 106960 7644
rect 106664 7590 106710 7642
rect 106710 7590 106720 7642
rect 106744 7590 106774 7642
rect 106774 7590 106786 7642
rect 106786 7590 106800 7642
rect 106824 7590 106838 7642
rect 106838 7590 106850 7642
rect 106850 7590 106880 7642
rect 106904 7590 106914 7642
rect 106914 7590 106960 7642
rect 106664 7588 106720 7590
rect 106744 7588 106800 7590
rect 106824 7588 106880 7590
rect 106904 7588 106960 7590
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 105928 7098 105984 7100
rect 106008 7098 106064 7100
rect 106088 7098 106144 7100
rect 106168 7098 106224 7100
rect 105928 7046 105974 7098
rect 105974 7046 105984 7098
rect 106008 7046 106038 7098
rect 106038 7046 106050 7098
rect 106050 7046 106064 7098
rect 106088 7046 106102 7098
rect 106102 7046 106114 7098
rect 106114 7046 106144 7098
rect 106168 7046 106178 7098
rect 106178 7046 106224 7098
rect 105928 7044 105984 7046
rect 106008 7044 106064 7046
rect 106088 7044 106144 7046
rect 106168 7044 106224 7046
rect 66320 6554 66376 6556
rect 66400 6554 66456 6556
rect 66480 6554 66536 6556
rect 66560 6554 66616 6556
rect 66320 6502 66366 6554
rect 66366 6502 66376 6554
rect 66400 6502 66430 6554
rect 66430 6502 66442 6554
rect 66442 6502 66456 6554
rect 66480 6502 66494 6554
rect 66494 6502 66506 6554
rect 66506 6502 66536 6554
rect 66560 6502 66570 6554
rect 66570 6502 66616 6554
rect 66320 6500 66376 6502
rect 66400 6500 66456 6502
rect 66480 6500 66536 6502
rect 66560 6500 66616 6502
rect 97040 6554 97096 6556
rect 97120 6554 97176 6556
rect 97200 6554 97256 6556
rect 97280 6554 97336 6556
rect 97040 6502 97086 6554
rect 97086 6502 97096 6554
rect 97120 6502 97150 6554
rect 97150 6502 97162 6554
rect 97162 6502 97176 6554
rect 97200 6502 97214 6554
rect 97214 6502 97226 6554
rect 97226 6502 97256 6554
rect 97280 6502 97290 6554
rect 97290 6502 97336 6554
rect 97040 6500 97096 6502
rect 97120 6500 97176 6502
rect 97200 6500 97256 6502
rect 97280 6500 97336 6502
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 66320 5466 66376 5468
rect 66400 5466 66456 5468
rect 66480 5466 66536 5468
rect 66560 5466 66616 5468
rect 66320 5414 66366 5466
rect 66366 5414 66376 5466
rect 66400 5414 66430 5466
rect 66430 5414 66442 5466
rect 66442 5414 66456 5466
rect 66480 5414 66494 5466
rect 66494 5414 66506 5466
rect 66506 5414 66536 5466
rect 66560 5414 66570 5466
rect 66570 5414 66616 5466
rect 66320 5412 66376 5414
rect 66400 5412 66456 5414
rect 66480 5412 66536 5414
rect 66560 5412 66616 5414
rect 97040 5466 97096 5468
rect 97120 5466 97176 5468
rect 97200 5466 97256 5468
rect 97280 5466 97336 5468
rect 97040 5414 97086 5466
rect 97086 5414 97096 5466
rect 97120 5414 97150 5466
rect 97150 5414 97162 5466
rect 97162 5414 97176 5466
rect 97200 5414 97214 5466
rect 97214 5414 97226 5466
rect 97226 5414 97256 5466
rect 97280 5414 97290 5466
rect 97290 5414 97336 5466
rect 97040 5412 97096 5414
rect 97120 5412 97176 5414
rect 97200 5412 97256 5414
rect 97280 5412 97336 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 66320 4378 66376 4380
rect 66400 4378 66456 4380
rect 66480 4378 66536 4380
rect 66560 4378 66616 4380
rect 66320 4326 66366 4378
rect 66366 4326 66376 4378
rect 66400 4326 66430 4378
rect 66430 4326 66442 4378
rect 66442 4326 66456 4378
rect 66480 4326 66494 4378
rect 66494 4326 66506 4378
rect 66506 4326 66536 4378
rect 66560 4326 66570 4378
rect 66570 4326 66616 4378
rect 66320 4324 66376 4326
rect 66400 4324 66456 4326
rect 66480 4324 66536 4326
rect 66560 4324 66616 4326
rect 97040 4378 97096 4380
rect 97120 4378 97176 4380
rect 97200 4378 97256 4380
rect 97280 4378 97336 4380
rect 97040 4326 97086 4378
rect 97086 4326 97096 4378
rect 97120 4326 97150 4378
rect 97150 4326 97162 4378
rect 97162 4326 97176 4378
rect 97200 4326 97214 4378
rect 97214 4326 97226 4378
rect 97226 4326 97256 4378
rect 97280 4326 97290 4378
rect 97290 4326 97336 4378
rect 97040 4324 97096 4326
rect 97120 4324 97176 4326
rect 97200 4324 97256 4326
rect 97280 4324 97336 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 66320 3290 66376 3292
rect 66400 3290 66456 3292
rect 66480 3290 66536 3292
rect 66560 3290 66616 3292
rect 66320 3238 66366 3290
rect 66366 3238 66376 3290
rect 66400 3238 66430 3290
rect 66430 3238 66442 3290
rect 66442 3238 66456 3290
rect 66480 3238 66494 3290
rect 66494 3238 66506 3290
rect 66506 3238 66536 3290
rect 66560 3238 66570 3290
rect 66570 3238 66616 3290
rect 66320 3236 66376 3238
rect 66400 3236 66456 3238
rect 66480 3236 66536 3238
rect 66560 3236 66616 3238
rect 97040 3290 97096 3292
rect 97120 3290 97176 3292
rect 97200 3290 97256 3292
rect 97280 3290 97336 3292
rect 97040 3238 97086 3290
rect 97086 3238 97096 3290
rect 97120 3238 97150 3290
rect 97150 3238 97162 3290
rect 97162 3238 97176 3290
rect 97200 3238 97214 3290
rect 97214 3238 97226 3290
rect 97226 3238 97256 3290
rect 97280 3238 97290 3290
rect 97290 3238 97336 3290
rect 97040 3236 97096 3238
rect 97120 3236 97176 3238
rect 97200 3236 97256 3238
rect 97280 3236 97336 3238
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 66320 2202 66376 2204
rect 66400 2202 66456 2204
rect 66480 2202 66536 2204
rect 66560 2202 66616 2204
rect 66320 2150 66366 2202
rect 66366 2150 66376 2202
rect 66400 2150 66430 2202
rect 66430 2150 66442 2202
rect 66442 2150 66456 2202
rect 66480 2150 66494 2202
rect 66494 2150 66506 2202
rect 66506 2150 66536 2202
rect 66560 2150 66570 2202
rect 66570 2150 66616 2202
rect 66320 2148 66376 2150
rect 66400 2148 66456 2150
rect 66480 2148 66536 2150
rect 66560 2148 66616 2150
rect 97040 2202 97096 2204
rect 97120 2202 97176 2204
rect 97200 2202 97256 2204
rect 97280 2202 97336 2204
rect 97040 2150 97086 2202
rect 97086 2150 97096 2202
rect 97120 2150 97150 2202
rect 97150 2150 97162 2202
rect 97162 2150 97176 2202
rect 97200 2150 97214 2202
rect 97214 2150 97226 2202
rect 97226 2150 97256 2202
rect 97280 2150 97290 2202
rect 97290 2150 97336 2202
rect 97040 2148 97096 2150
rect 97120 2148 97176 2150
rect 97200 2148 97256 2150
rect 97280 2148 97336 2150
<< metal3 >>
rect 4210 147456 4526 147457
rect 4210 147392 4216 147456
rect 4280 147392 4296 147456
rect 4360 147392 4376 147456
rect 4440 147392 4456 147456
rect 4520 147392 4526 147456
rect 4210 147391 4526 147392
rect 34930 147456 35246 147457
rect 34930 147392 34936 147456
rect 35000 147392 35016 147456
rect 35080 147392 35096 147456
rect 35160 147392 35176 147456
rect 35240 147392 35246 147456
rect 34930 147391 35246 147392
rect 65650 147456 65966 147457
rect 65650 147392 65656 147456
rect 65720 147392 65736 147456
rect 65800 147392 65816 147456
rect 65880 147392 65896 147456
rect 65960 147392 65966 147456
rect 65650 147391 65966 147392
rect 96370 147456 96686 147457
rect 96370 147392 96376 147456
rect 96440 147392 96456 147456
rect 96520 147392 96536 147456
rect 96600 147392 96616 147456
rect 96680 147392 96686 147456
rect 96370 147391 96686 147392
rect 4870 146912 5186 146913
rect 4870 146848 4876 146912
rect 4940 146848 4956 146912
rect 5020 146848 5036 146912
rect 5100 146848 5116 146912
rect 5180 146848 5186 146912
rect 4870 146847 5186 146848
rect 35590 146912 35906 146913
rect 35590 146848 35596 146912
rect 35660 146848 35676 146912
rect 35740 146848 35756 146912
rect 35820 146848 35836 146912
rect 35900 146848 35906 146912
rect 35590 146847 35906 146848
rect 66310 146912 66626 146913
rect 66310 146848 66316 146912
rect 66380 146848 66396 146912
rect 66460 146848 66476 146912
rect 66540 146848 66556 146912
rect 66620 146848 66626 146912
rect 66310 146847 66626 146848
rect 97030 146912 97346 146913
rect 97030 146848 97036 146912
rect 97100 146848 97116 146912
rect 97180 146848 97196 146912
rect 97260 146848 97276 146912
rect 97340 146848 97346 146912
rect 97030 146847 97346 146848
rect 4210 146368 4526 146369
rect 4210 146304 4216 146368
rect 4280 146304 4296 146368
rect 4360 146304 4376 146368
rect 4440 146304 4456 146368
rect 4520 146304 4526 146368
rect 4210 146303 4526 146304
rect 34930 146368 35246 146369
rect 34930 146304 34936 146368
rect 35000 146304 35016 146368
rect 35080 146304 35096 146368
rect 35160 146304 35176 146368
rect 35240 146304 35246 146368
rect 34930 146303 35246 146304
rect 65650 146368 65966 146369
rect 65650 146304 65656 146368
rect 65720 146304 65736 146368
rect 65800 146304 65816 146368
rect 65880 146304 65896 146368
rect 65960 146304 65966 146368
rect 65650 146303 65966 146304
rect 96370 146368 96686 146369
rect 96370 146304 96376 146368
rect 96440 146304 96456 146368
rect 96520 146304 96536 146368
rect 96600 146304 96616 146368
rect 96680 146304 96686 146368
rect 96370 146303 96686 146304
rect 4870 145824 5186 145825
rect 4870 145760 4876 145824
rect 4940 145760 4956 145824
rect 5020 145760 5036 145824
rect 5100 145760 5116 145824
rect 5180 145760 5186 145824
rect 4870 145759 5186 145760
rect 35590 145824 35906 145825
rect 35590 145760 35596 145824
rect 35660 145760 35676 145824
rect 35740 145760 35756 145824
rect 35820 145760 35836 145824
rect 35900 145760 35906 145824
rect 35590 145759 35906 145760
rect 66310 145824 66626 145825
rect 66310 145760 66316 145824
rect 66380 145760 66396 145824
rect 66460 145760 66476 145824
rect 66540 145760 66556 145824
rect 66620 145760 66626 145824
rect 66310 145759 66626 145760
rect 97030 145824 97346 145825
rect 97030 145760 97036 145824
rect 97100 145760 97116 145824
rect 97180 145760 97196 145824
rect 97260 145760 97276 145824
rect 97340 145760 97346 145824
rect 97030 145759 97346 145760
rect 4210 145280 4526 145281
rect 4210 145216 4216 145280
rect 4280 145216 4296 145280
rect 4360 145216 4376 145280
rect 4440 145216 4456 145280
rect 4520 145216 4526 145280
rect 4210 145215 4526 145216
rect 34930 145280 35246 145281
rect 34930 145216 34936 145280
rect 35000 145216 35016 145280
rect 35080 145216 35096 145280
rect 35160 145216 35176 145280
rect 35240 145216 35246 145280
rect 34930 145215 35246 145216
rect 65650 145280 65966 145281
rect 65650 145216 65656 145280
rect 65720 145216 65736 145280
rect 65800 145216 65816 145280
rect 65880 145216 65896 145280
rect 65960 145216 65966 145280
rect 65650 145215 65966 145216
rect 96370 145280 96686 145281
rect 96370 145216 96376 145280
rect 96440 145216 96456 145280
rect 96520 145216 96536 145280
rect 96600 145216 96616 145280
rect 96680 145216 96686 145280
rect 96370 145215 96686 145216
rect 4870 144736 5186 144737
rect 4870 144672 4876 144736
rect 4940 144672 4956 144736
rect 5020 144672 5036 144736
rect 5100 144672 5116 144736
rect 5180 144672 5186 144736
rect 4870 144671 5186 144672
rect 35590 144736 35906 144737
rect 35590 144672 35596 144736
rect 35660 144672 35676 144736
rect 35740 144672 35756 144736
rect 35820 144672 35836 144736
rect 35900 144672 35906 144736
rect 35590 144671 35906 144672
rect 66310 144736 66626 144737
rect 66310 144672 66316 144736
rect 66380 144672 66396 144736
rect 66460 144672 66476 144736
rect 66540 144672 66556 144736
rect 66620 144672 66626 144736
rect 66310 144671 66626 144672
rect 97030 144736 97346 144737
rect 97030 144672 97036 144736
rect 97100 144672 97116 144736
rect 97180 144672 97196 144736
rect 97260 144672 97276 144736
rect 97340 144672 97346 144736
rect 97030 144671 97346 144672
rect 4210 144192 4526 144193
rect 4210 144128 4216 144192
rect 4280 144128 4296 144192
rect 4360 144128 4376 144192
rect 4440 144128 4456 144192
rect 4520 144128 4526 144192
rect 4210 144127 4526 144128
rect 34930 144192 35246 144193
rect 34930 144128 34936 144192
rect 35000 144128 35016 144192
rect 35080 144128 35096 144192
rect 35160 144128 35176 144192
rect 35240 144128 35246 144192
rect 34930 144127 35246 144128
rect 65650 144192 65966 144193
rect 65650 144128 65656 144192
rect 65720 144128 65736 144192
rect 65800 144128 65816 144192
rect 65880 144128 65896 144192
rect 65960 144128 65966 144192
rect 65650 144127 65966 144128
rect 96370 144192 96686 144193
rect 96370 144128 96376 144192
rect 96440 144128 96456 144192
rect 96520 144128 96536 144192
rect 96600 144128 96616 144192
rect 96680 144128 96686 144192
rect 96370 144127 96686 144128
rect 4870 143648 5186 143649
rect 4870 143584 4876 143648
rect 4940 143584 4956 143648
rect 5020 143584 5036 143648
rect 5100 143584 5116 143648
rect 5180 143584 5186 143648
rect 4870 143583 5186 143584
rect 35590 143648 35906 143649
rect 35590 143584 35596 143648
rect 35660 143584 35676 143648
rect 35740 143584 35756 143648
rect 35820 143584 35836 143648
rect 35900 143584 35906 143648
rect 35590 143583 35906 143584
rect 66310 143648 66626 143649
rect 66310 143584 66316 143648
rect 66380 143584 66396 143648
rect 66460 143584 66476 143648
rect 66540 143584 66556 143648
rect 66620 143584 66626 143648
rect 66310 143583 66626 143584
rect 97030 143648 97346 143649
rect 97030 143584 97036 143648
rect 97100 143584 97116 143648
rect 97180 143584 97196 143648
rect 97260 143584 97276 143648
rect 97340 143584 97346 143648
rect 97030 143583 97346 143584
rect 4210 143104 4526 143105
rect 4210 143040 4216 143104
rect 4280 143040 4296 143104
rect 4360 143040 4376 143104
rect 4440 143040 4456 143104
rect 4520 143040 4526 143104
rect 4210 143039 4526 143040
rect 34930 143104 35246 143105
rect 34930 143040 34936 143104
rect 35000 143040 35016 143104
rect 35080 143040 35096 143104
rect 35160 143040 35176 143104
rect 35240 143040 35246 143104
rect 34930 143039 35246 143040
rect 65650 143104 65966 143105
rect 65650 143040 65656 143104
rect 65720 143040 65736 143104
rect 65800 143040 65816 143104
rect 65880 143040 65896 143104
rect 65960 143040 65966 143104
rect 65650 143039 65966 143040
rect 96370 143104 96686 143105
rect 96370 143040 96376 143104
rect 96440 143040 96456 143104
rect 96520 143040 96536 143104
rect 96600 143040 96616 143104
rect 96680 143040 96686 143104
rect 96370 143039 96686 143040
rect 4870 142560 5186 142561
rect 4870 142496 4876 142560
rect 4940 142496 4956 142560
rect 5020 142496 5036 142560
rect 5100 142496 5116 142560
rect 5180 142496 5186 142560
rect 4870 142495 5186 142496
rect 35590 142560 35906 142561
rect 35590 142496 35596 142560
rect 35660 142496 35676 142560
rect 35740 142496 35756 142560
rect 35820 142496 35836 142560
rect 35900 142496 35906 142560
rect 35590 142495 35906 142496
rect 66310 142560 66626 142561
rect 66310 142496 66316 142560
rect 66380 142496 66396 142560
rect 66460 142496 66476 142560
rect 66540 142496 66556 142560
rect 66620 142496 66626 142560
rect 66310 142495 66626 142496
rect 97030 142560 97346 142561
rect 97030 142496 97036 142560
rect 97100 142496 97116 142560
rect 97180 142496 97196 142560
rect 97260 142496 97276 142560
rect 97340 142496 97346 142560
rect 97030 142495 97346 142496
rect 4210 142016 4526 142017
rect 4210 141952 4216 142016
rect 4280 141952 4296 142016
rect 4360 141952 4376 142016
rect 4440 141952 4456 142016
rect 4520 141952 4526 142016
rect 4210 141951 4526 141952
rect 34930 142016 35246 142017
rect 34930 141952 34936 142016
rect 35000 141952 35016 142016
rect 35080 141952 35096 142016
rect 35160 141952 35176 142016
rect 35240 141952 35246 142016
rect 34930 141951 35246 141952
rect 65650 142016 65966 142017
rect 65650 141952 65656 142016
rect 65720 141952 65736 142016
rect 65800 141952 65816 142016
rect 65880 141952 65896 142016
rect 65960 141952 65966 142016
rect 65650 141951 65966 141952
rect 96370 142016 96686 142017
rect 96370 141952 96376 142016
rect 96440 141952 96456 142016
rect 96520 141952 96536 142016
rect 96600 141952 96616 142016
rect 96680 141952 96686 142016
rect 96370 141951 96686 141952
rect 4870 141472 5186 141473
rect 4870 141408 4876 141472
rect 4940 141408 4956 141472
rect 5020 141408 5036 141472
rect 5100 141408 5116 141472
rect 5180 141408 5186 141472
rect 4870 141407 5186 141408
rect 35590 141472 35906 141473
rect 35590 141408 35596 141472
rect 35660 141408 35676 141472
rect 35740 141408 35756 141472
rect 35820 141408 35836 141472
rect 35900 141408 35906 141472
rect 35590 141407 35906 141408
rect 66310 141472 66626 141473
rect 66310 141408 66316 141472
rect 66380 141408 66396 141472
rect 66460 141408 66476 141472
rect 66540 141408 66556 141472
rect 66620 141408 66626 141472
rect 66310 141407 66626 141408
rect 97030 141472 97346 141473
rect 97030 141408 97036 141472
rect 97100 141408 97116 141472
rect 97180 141408 97196 141472
rect 97260 141408 97276 141472
rect 97340 141408 97346 141472
rect 97030 141407 97346 141408
rect 4210 140928 4526 140929
rect 4210 140864 4216 140928
rect 4280 140864 4296 140928
rect 4360 140864 4376 140928
rect 4440 140864 4456 140928
rect 4520 140864 4526 140928
rect 4210 140863 4526 140864
rect 34930 140928 35246 140929
rect 34930 140864 34936 140928
rect 35000 140864 35016 140928
rect 35080 140864 35096 140928
rect 35160 140864 35176 140928
rect 35240 140864 35246 140928
rect 34930 140863 35246 140864
rect 65650 140928 65966 140929
rect 65650 140864 65656 140928
rect 65720 140864 65736 140928
rect 65800 140864 65816 140928
rect 65880 140864 65896 140928
rect 65960 140864 65966 140928
rect 65650 140863 65966 140864
rect 96370 140928 96686 140929
rect 96370 140864 96376 140928
rect 96440 140864 96456 140928
rect 96520 140864 96536 140928
rect 96600 140864 96616 140928
rect 96680 140864 96686 140928
rect 96370 140863 96686 140864
rect 4870 140384 5186 140385
rect 4870 140320 4876 140384
rect 4940 140320 4956 140384
rect 5020 140320 5036 140384
rect 5100 140320 5116 140384
rect 5180 140320 5186 140384
rect 4870 140319 5186 140320
rect 35590 140384 35906 140385
rect 35590 140320 35596 140384
rect 35660 140320 35676 140384
rect 35740 140320 35756 140384
rect 35820 140320 35836 140384
rect 35900 140320 35906 140384
rect 35590 140319 35906 140320
rect 66310 140384 66626 140385
rect 66310 140320 66316 140384
rect 66380 140320 66396 140384
rect 66460 140320 66476 140384
rect 66540 140320 66556 140384
rect 66620 140320 66626 140384
rect 66310 140319 66626 140320
rect 97030 140384 97346 140385
rect 97030 140320 97036 140384
rect 97100 140320 97116 140384
rect 97180 140320 97196 140384
rect 97260 140320 97276 140384
rect 97340 140320 97346 140384
rect 97030 140319 97346 140320
rect 4210 139840 4526 139841
rect 4210 139776 4216 139840
rect 4280 139776 4296 139840
rect 4360 139776 4376 139840
rect 4440 139776 4456 139840
rect 4520 139776 4526 139840
rect 4210 139775 4526 139776
rect 34930 139840 35246 139841
rect 34930 139776 34936 139840
rect 35000 139776 35016 139840
rect 35080 139776 35096 139840
rect 35160 139776 35176 139840
rect 35240 139776 35246 139840
rect 34930 139775 35246 139776
rect 65650 139840 65966 139841
rect 65650 139776 65656 139840
rect 65720 139776 65736 139840
rect 65800 139776 65816 139840
rect 65880 139776 65896 139840
rect 65960 139776 65966 139840
rect 65650 139775 65966 139776
rect 96370 139840 96686 139841
rect 96370 139776 96376 139840
rect 96440 139776 96456 139840
rect 96520 139776 96536 139840
rect 96600 139776 96616 139840
rect 96680 139776 96686 139840
rect 96370 139775 96686 139776
rect 4870 139296 5186 139297
rect 4870 139232 4876 139296
rect 4940 139232 4956 139296
rect 5020 139232 5036 139296
rect 5100 139232 5116 139296
rect 5180 139232 5186 139296
rect 4870 139231 5186 139232
rect 35590 139296 35906 139297
rect 35590 139232 35596 139296
rect 35660 139232 35676 139296
rect 35740 139232 35756 139296
rect 35820 139232 35836 139296
rect 35900 139232 35906 139296
rect 35590 139231 35906 139232
rect 66310 139296 66626 139297
rect 66310 139232 66316 139296
rect 66380 139232 66396 139296
rect 66460 139232 66476 139296
rect 66540 139232 66556 139296
rect 66620 139232 66626 139296
rect 66310 139231 66626 139232
rect 97030 139296 97346 139297
rect 97030 139232 97036 139296
rect 97100 139232 97116 139296
rect 97180 139232 97196 139296
rect 97260 139232 97276 139296
rect 97340 139232 97346 139296
rect 97030 139231 97346 139232
rect 4210 138752 4526 138753
rect 4210 138688 4216 138752
rect 4280 138688 4296 138752
rect 4360 138688 4376 138752
rect 4440 138688 4456 138752
rect 4520 138688 4526 138752
rect 4210 138687 4526 138688
rect 34930 138752 35246 138753
rect 34930 138688 34936 138752
rect 35000 138688 35016 138752
rect 35080 138688 35096 138752
rect 35160 138688 35176 138752
rect 35240 138688 35246 138752
rect 34930 138687 35246 138688
rect 65650 138752 65966 138753
rect 65650 138688 65656 138752
rect 65720 138688 65736 138752
rect 65800 138688 65816 138752
rect 65880 138688 65896 138752
rect 65960 138688 65966 138752
rect 65650 138687 65966 138688
rect 96370 138752 96686 138753
rect 96370 138688 96376 138752
rect 96440 138688 96456 138752
rect 96520 138688 96536 138752
rect 96600 138688 96616 138752
rect 96680 138688 96686 138752
rect 96370 138687 96686 138688
rect 4870 138208 5186 138209
rect 4870 138144 4876 138208
rect 4940 138144 4956 138208
rect 5020 138144 5036 138208
rect 5100 138144 5116 138208
rect 5180 138144 5186 138208
rect 4870 138143 5186 138144
rect 35590 138208 35906 138209
rect 35590 138144 35596 138208
rect 35660 138144 35676 138208
rect 35740 138144 35756 138208
rect 35820 138144 35836 138208
rect 35900 138144 35906 138208
rect 35590 138143 35906 138144
rect 66310 138208 66626 138209
rect 66310 138144 66316 138208
rect 66380 138144 66396 138208
rect 66460 138144 66476 138208
rect 66540 138144 66556 138208
rect 66620 138144 66626 138208
rect 66310 138143 66626 138144
rect 97030 138208 97346 138209
rect 97030 138144 97036 138208
rect 97100 138144 97116 138208
rect 97180 138144 97196 138208
rect 97260 138144 97276 138208
rect 97340 138144 97346 138208
rect 97030 138143 97346 138144
rect 4210 137664 4526 137665
rect 4210 137600 4216 137664
rect 4280 137600 4296 137664
rect 4360 137600 4376 137664
rect 4440 137600 4456 137664
rect 4520 137600 4526 137664
rect 4210 137599 4526 137600
rect 34930 137664 35246 137665
rect 34930 137600 34936 137664
rect 35000 137600 35016 137664
rect 35080 137600 35096 137664
rect 35160 137600 35176 137664
rect 35240 137600 35246 137664
rect 34930 137599 35246 137600
rect 65650 137664 65966 137665
rect 65650 137600 65656 137664
rect 65720 137600 65736 137664
rect 65800 137600 65816 137664
rect 65880 137600 65896 137664
rect 65960 137600 65966 137664
rect 65650 137599 65966 137600
rect 96370 137664 96686 137665
rect 96370 137600 96376 137664
rect 96440 137600 96456 137664
rect 96520 137600 96536 137664
rect 96600 137600 96616 137664
rect 96680 137600 96686 137664
rect 96370 137599 96686 137600
rect 4870 137120 5186 137121
rect 4870 137056 4876 137120
rect 4940 137056 4956 137120
rect 5020 137056 5036 137120
rect 5100 137056 5116 137120
rect 5180 137056 5186 137120
rect 4870 137055 5186 137056
rect 35590 137120 35906 137121
rect 35590 137056 35596 137120
rect 35660 137056 35676 137120
rect 35740 137056 35756 137120
rect 35820 137056 35836 137120
rect 35900 137056 35906 137120
rect 35590 137055 35906 137056
rect 66310 137120 66626 137121
rect 66310 137056 66316 137120
rect 66380 137056 66396 137120
rect 66460 137056 66476 137120
rect 66540 137056 66556 137120
rect 66620 137056 66626 137120
rect 66310 137055 66626 137056
rect 97030 137120 97346 137121
rect 97030 137056 97036 137120
rect 97100 137056 97116 137120
rect 97180 137056 97196 137120
rect 97260 137056 97276 137120
rect 97340 137056 97346 137120
rect 97030 137055 97346 137056
rect 4210 136576 4526 136577
rect 4210 136512 4216 136576
rect 4280 136512 4296 136576
rect 4360 136512 4376 136576
rect 4440 136512 4456 136576
rect 4520 136512 4526 136576
rect 4210 136511 4526 136512
rect 34930 136576 35246 136577
rect 34930 136512 34936 136576
rect 35000 136512 35016 136576
rect 35080 136512 35096 136576
rect 35160 136512 35176 136576
rect 35240 136512 35246 136576
rect 34930 136511 35246 136512
rect 65650 136576 65966 136577
rect 65650 136512 65656 136576
rect 65720 136512 65736 136576
rect 65800 136512 65816 136576
rect 65880 136512 65896 136576
rect 65960 136512 65966 136576
rect 65650 136511 65966 136512
rect 96370 136576 96686 136577
rect 96370 136512 96376 136576
rect 96440 136512 96456 136576
rect 96520 136512 96536 136576
rect 96600 136512 96616 136576
rect 96680 136512 96686 136576
rect 96370 136511 96686 136512
rect 105918 136576 106234 136577
rect 105918 136512 105924 136576
rect 105988 136512 106004 136576
rect 106068 136512 106084 136576
rect 106148 136512 106164 136576
rect 106228 136512 106234 136576
rect 105918 136511 106234 136512
rect 4870 136032 5186 136033
rect 4870 135968 4876 136032
rect 4940 135968 4956 136032
rect 5020 135968 5036 136032
rect 5100 135968 5116 136032
rect 5180 135968 5186 136032
rect 4870 135967 5186 135968
rect 35590 136032 35906 136033
rect 35590 135968 35596 136032
rect 35660 135968 35676 136032
rect 35740 135968 35756 136032
rect 35820 135968 35836 136032
rect 35900 135968 35906 136032
rect 35590 135967 35906 135968
rect 66310 136032 66626 136033
rect 66310 135968 66316 136032
rect 66380 135968 66396 136032
rect 66460 135968 66476 136032
rect 66540 135968 66556 136032
rect 66620 135968 66626 136032
rect 66310 135967 66626 135968
rect 97030 136032 97346 136033
rect 97030 135968 97036 136032
rect 97100 135968 97116 136032
rect 97180 135968 97196 136032
rect 97260 135968 97276 136032
rect 97340 135968 97346 136032
rect 97030 135967 97346 135968
rect 106654 136032 106970 136033
rect 106654 135968 106660 136032
rect 106724 135968 106740 136032
rect 106804 135968 106820 136032
rect 106884 135968 106900 136032
rect 106964 135968 106970 136032
rect 106654 135967 106970 135968
rect 95969 135692 96035 135693
rect 95918 135690 95924 135692
rect 95878 135630 95924 135690
rect 95988 135688 96035 135692
rect 96030 135632 96035 135688
rect 95918 135628 95924 135630
rect 95988 135628 96035 135632
rect 95969 135627 96035 135628
rect 4210 135488 4526 135489
rect 4210 135424 4216 135488
rect 4280 135424 4296 135488
rect 4360 135424 4376 135488
rect 4440 135424 4456 135488
rect 4520 135424 4526 135488
rect 4210 135423 4526 135424
rect 105918 135488 106234 135489
rect 105918 135424 105924 135488
rect 105988 135424 106004 135488
rect 106068 135424 106084 135488
rect 106148 135424 106164 135488
rect 106228 135424 106234 135488
rect 105918 135423 106234 135424
rect 58566 135220 58572 135284
rect 58636 135282 58642 135284
rect 60549 135282 60615 135285
rect 58636 135280 60615 135282
rect 58636 135224 60554 135280
rect 60610 135224 60615 135280
rect 58636 135222 60615 135224
rect 58636 135220 58642 135222
rect 60549 135219 60615 135222
rect 61142 135220 61148 135284
rect 61212 135282 61218 135284
rect 63125 135282 63191 135285
rect 61212 135280 63191 135282
rect 61212 135224 63130 135280
rect 63186 135224 63191 135280
rect 61212 135222 63191 135224
rect 61212 135220 61218 135222
rect 63125 135219 63191 135222
rect 71078 135220 71084 135284
rect 71148 135282 71154 135284
rect 72693 135282 72759 135285
rect 71148 135280 72759 135282
rect 71148 135224 72698 135280
rect 72754 135224 72759 135280
rect 71148 135222 72759 135224
rect 71148 135220 71154 135222
rect 72693 135219 72759 135222
rect 63585 135148 63651 135149
rect 63534 135084 63540 135148
rect 63604 135146 63651 135148
rect 63604 135144 63696 135146
rect 63646 135088 63696 135144
rect 63604 135086 63696 135088
rect 63604 135084 63651 135086
rect 63585 135083 63651 135084
rect 4870 134944 5186 134945
rect 4870 134880 4876 134944
rect 4940 134880 4956 134944
rect 5020 134880 5036 134944
rect 5100 134880 5116 134944
rect 5180 134880 5186 134944
rect 4870 134879 5186 134880
rect 106654 134944 106970 134945
rect 106654 134880 106660 134944
rect 106724 134880 106740 134944
rect 106804 134880 106820 134944
rect 106884 134880 106900 134944
rect 106964 134880 106970 134944
rect 106654 134879 106970 134880
rect 73470 134404 73476 134468
rect 73540 134466 73546 134468
rect 77385 134466 77451 134469
rect 73540 134464 77451 134466
rect 73540 134408 77390 134464
rect 77446 134408 77451 134464
rect 73540 134406 77451 134408
rect 73540 134404 73546 134406
rect 77385 134403 77451 134406
rect 4210 134400 4526 134401
rect 4210 134336 4216 134400
rect 4280 134336 4296 134400
rect 4360 134336 4376 134400
rect 4440 134336 4456 134400
rect 4520 134336 4526 134400
rect 4210 134335 4526 134336
rect 105918 134400 106234 134401
rect 105918 134336 105924 134400
rect 105988 134336 106004 134400
rect 106068 134336 106084 134400
rect 106148 134336 106164 134400
rect 106228 134336 106234 134400
rect 105918 134335 106234 134336
rect 38745 134194 38811 134197
rect 41061 134194 41067 134196
rect 38745 134192 41067 134194
rect 38745 134136 38750 134192
rect 38806 134136 41067 134192
rect 38745 134134 41067 134136
rect 38745 134131 38811 134134
rect 41061 134132 41067 134134
rect 41131 134132 41137 134196
rect 43161 134194 43227 134197
rect 43557 134194 43563 134196
rect 43161 134192 43563 134194
rect 43161 134136 43166 134192
rect 43222 134136 43563 134192
rect 43161 134134 43563 134136
rect 43161 134131 43227 134134
rect 43557 134132 43563 134134
rect 43627 134132 43633 134196
rect 53541 134132 53547 134196
rect 53611 134194 53617 134196
rect 55397 134194 55463 134197
rect 53611 134192 55463 134194
rect 53611 134136 55402 134192
rect 55458 134136 55463 134192
rect 53611 134134 55463 134136
rect 53611 134132 53617 134134
rect 55397 134131 55463 134134
rect 56037 134132 56043 134196
rect 56107 134194 56113 134196
rect 57973 134194 58039 134197
rect 56107 134192 58039 134194
rect 56107 134136 57978 134192
rect 58034 134136 58039 134192
rect 56107 134134 58039 134136
rect 56107 134132 56113 134134
rect 57973 134131 58039 134134
rect 66021 134132 66027 134196
rect 66091 134194 66097 134196
rect 72509 134194 72575 134197
rect 66091 134192 72575 134194
rect 66091 134136 72514 134192
rect 72570 134136 72575 134192
rect 66091 134134 72575 134136
rect 66091 134132 66097 134134
rect 72509 134131 72575 134134
rect 36077 133924 36143 133925
rect 38561 133924 38627 133925
rect 46105 133924 46171 133925
rect 36069 133860 36075 133924
rect 36139 133922 36145 133924
rect 38561 133922 38571 133924
rect 36139 133862 36231 133922
rect 38479 133920 38571 133922
rect 38479 133864 38566 133920
rect 38479 133862 38571 133864
rect 36139 133860 36145 133862
rect 38561 133860 38571 133862
rect 38635 133860 38641 133924
rect 46054 133922 46060 133924
rect 46014 133862 46060 133922
rect 46124 133920 46171 133924
rect 46166 133864 46171 133920
rect 46054 133860 46060 133862
rect 46124 133860 46171 133864
rect 36077 133859 36143 133860
rect 38561 133859 38627 133860
rect 46105 133859 46171 133860
rect 48497 133924 48563 133925
rect 51073 133924 51139 133925
rect 68553 133924 68619 133925
rect 48497 133920 48544 133924
rect 48608 133922 48614 133924
rect 51045 133922 51051 133924
rect 48497 133864 48502 133920
rect 48497 133860 48544 133864
rect 48608 133862 48654 133922
rect 50982 133862 51051 133922
rect 51115 133920 51139 133924
rect 68517 133922 68523 133924
rect 51134 133864 51139 133920
rect 48608 133860 48614 133862
rect 51045 133860 51051 133862
rect 51115 133860 51139 133864
rect 68462 133862 68523 133922
rect 68587 133920 68619 133924
rect 68614 133864 68619 133920
rect 68517 133860 68523 133862
rect 68587 133860 68619 133864
rect 86136 133860 86142 133924
rect 86206 133922 86212 133924
rect 86309 133922 86375 133925
rect 87321 133924 87387 133925
rect 87304 133922 87310 133924
rect 86206 133920 86375 133922
rect 86206 133864 86314 133920
rect 86370 133864 86375 133920
rect 86206 133862 86375 133864
rect 87230 133862 87310 133922
rect 87374 133920 87387 133924
rect 87382 133864 87387 133920
rect 86206 133860 86212 133862
rect 48497 133859 48563 133860
rect 51073 133859 51139 133860
rect 68553 133859 68619 133860
rect 86309 133859 86375 133862
rect 87304 133860 87310 133862
rect 87374 133860 87387 133864
rect 87321 133859 87387 133860
rect 4870 133856 5186 133857
rect 4870 133792 4876 133856
rect 4940 133792 4956 133856
rect 5020 133792 5036 133856
rect 5100 133792 5116 133856
rect 5180 133792 5186 133856
rect 4870 133791 5186 133792
rect 106654 133856 106970 133857
rect 106654 133792 106660 133856
rect 106724 133792 106740 133856
rect 106804 133792 106820 133856
rect 106884 133792 106900 133856
rect 106964 133792 106970 133856
rect 106654 133791 106970 133792
rect 4210 133312 4526 133313
rect 4210 133248 4216 133312
rect 4280 133248 4296 133312
rect 4360 133248 4376 133312
rect 4440 133248 4456 133312
rect 4520 133248 4526 133312
rect 4210 133247 4526 133248
rect 105918 133312 106234 133313
rect 105918 133248 105924 133312
rect 105988 133248 106004 133312
rect 106068 133248 106084 133312
rect 106148 133248 106164 133312
rect 106228 133248 106234 133312
rect 105918 133247 106234 133248
rect 4870 132768 5186 132769
rect 4870 132704 4876 132768
rect 4940 132704 4956 132768
rect 5020 132704 5036 132768
rect 5100 132704 5116 132768
rect 5180 132704 5186 132768
rect 4870 132703 5186 132704
rect 106654 132768 106970 132769
rect 106654 132704 106660 132768
rect 106724 132704 106740 132768
rect 106804 132704 106820 132768
rect 106884 132704 106900 132768
rect 106964 132704 106970 132768
rect 106654 132703 106970 132704
rect 4210 132224 4526 132225
rect 4210 132160 4216 132224
rect 4280 132160 4296 132224
rect 4360 132160 4376 132224
rect 4440 132160 4456 132224
rect 4520 132160 4526 132224
rect 4210 132159 4526 132160
rect 105918 132224 106234 132225
rect 105918 132160 105924 132224
rect 105988 132160 106004 132224
rect 106068 132160 106084 132224
rect 106148 132160 106164 132224
rect 106228 132160 106234 132224
rect 105918 132159 106234 132160
rect 4870 131680 5186 131681
rect 4870 131616 4876 131680
rect 4940 131616 4956 131680
rect 5020 131616 5036 131680
rect 5100 131616 5116 131680
rect 5180 131616 5186 131680
rect 4870 131615 5186 131616
rect 106654 131680 106970 131681
rect 106654 131616 106660 131680
rect 106724 131616 106740 131680
rect 106804 131616 106820 131680
rect 106884 131616 106900 131680
rect 106964 131616 106970 131680
rect 106654 131615 106970 131616
rect 4210 131136 4526 131137
rect 4210 131072 4216 131136
rect 4280 131072 4296 131136
rect 4360 131072 4376 131136
rect 4440 131072 4456 131136
rect 4520 131072 4526 131136
rect 4210 131071 4526 131072
rect 105918 131136 106234 131137
rect 105918 131072 105924 131136
rect 105988 131072 106004 131136
rect 106068 131072 106084 131136
rect 106148 131072 106164 131136
rect 106228 131072 106234 131136
rect 105918 131071 106234 131072
rect 4870 130592 5186 130593
rect 4870 130528 4876 130592
rect 4940 130528 4956 130592
rect 5020 130528 5036 130592
rect 5100 130528 5116 130592
rect 5180 130528 5186 130592
rect 4870 130527 5186 130528
rect 106654 130592 106970 130593
rect 106654 130528 106660 130592
rect 106724 130528 106740 130592
rect 106804 130528 106820 130592
rect 106884 130528 106900 130592
rect 106964 130528 106970 130592
rect 106654 130527 106970 130528
rect 4210 130048 4526 130049
rect 4210 129984 4216 130048
rect 4280 129984 4296 130048
rect 4360 129984 4376 130048
rect 4440 129984 4456 130048
rect 4520 129984 4526 130048
rect 4210 129983 4526 129984
rect 105918 130048 106234 130049
rect 105918 129984 105924 130048
rect 105988 129984 106004 130048
rect 106068 129984 106084 130048
rect 106148 129984 106164 130048
rect 106228 129984 106234 130048
rect 105918 129983 106234 129984
rect 103881 129842 103947 129845
rect 102550 129840 103947 129842
rect 102550 129784 103886 129840
rect 103942 129784 103947 129840
rect 102550 129782 103947 129784
rect 102550 129768 102610 129782
rect 103881 129779 103947 129782
rect 101948 129708 102610 129768
rect 4870 129504 5186 129505
rect 4870 129440 4876 129504
rect 4940 129440 4956 129504
rect 5020 129440 5036 129504
rect 5100 129440 5116 129504
rect 5180 129440 5186 129504
rect 4870 129439 5186 129440
rect 106654 129504 106970 129505
rect 106654 129440 106660 129504
rect 106724 129440 106740 129504
rect 106804 129440 106820 129504
rect 106884 129440 106900 129504
rect 106964 129440 106970 129504
rect 106654 129439 106970 129440
rect 4210 128960 4526 128961
rect 4210 128896 4216 128960
rect 4280 128896 4296 128960
rect 4360 128896 4376 128960
rect 4440 128896 4456 128960
rect 4520 128896 4526 128960
rect 4210 128895 4526 128896
rect 105918 128960 106234 128961
rect 105918 128896 105924 128960
rect 105988 128896 106004 128960
rect 106068 128896 106084 128960
rect 106148 128896 106164 128960
rect 106228 128896 106234 128960
rect 105918 128895 106234 128896
rect 4870 128416 5186 128417
rect 4870 128352 4876 128416
rect 4940 128352 4956 128416
rect 5020 128352 5036 128416
rect 5100 128352 5116 128416
rect 5180 128352 5186 128416
rect 4870 128351 5186 128352
rect 106654 128416 106970 128417
rect 106654 128352 106660 128416
rect 106724 128352 106740 128416
rect 106804 128352 106820 128416
rect 106884 128352 106900 128416
rect 106964 128352 106970 128416
rect 106654 128351 106970 128352
rect 4210 127872 4526 127873
rect 4210 127808 4216 127872
rect 4280 127808 4296 127872
rect 4360 127808 4376 127872
rect 4440 127808 4456 127872
rect 4520 127808 4526 127872
rect 4210 127807 4526 127808
rect 105918 127872 106234 127873
rect 105918 127808 105924 127872
rect 105988 127808 106004 127872
rect 106068 127808 106084 127872
rect 106148 127808 106164 127872
rect 106228 127808 106234 127872
rect 105918 127807 106234 127808
rect 4870 127328 5186 127329
rect 4870 127264 4876 127328
rect 4940 127264 4956 127328
rect 5020 127264 5036 127328
rect 5100 127264 5116 127328
rect 5180 127264 5186 127328
rect 4870 127263 5186 127264
rect 106654 127328 106970 127329
rect 106654 127264 106660 127328
rect 106724 127264 106740 127328
rect 106804 127264 106820 127328
rect 106884 127264 106900 127328
rect 106964 127264 106970 127328
rect 106654 127263 106970 127264
rect 4210 126784 4526 126785
rect 4210 126720 4216 126784
rect 4280 126720 4296 126784
rect 4360 126720 4376 126784
rect 4440 126720 4456 126784
rect 4520 126720 4526 126784
rect 4210 126719 4526 126720
rect 105918 126784 106234 126785
rect 105918 126720 105924 126784
rect 105988 126720 106004 126784
rect 106068 126720 106084 126784
rect 106148 126720 106164 126784
rect 106228 126720 106234 126784
rect 105918 126719 106234 126720
rect 4870 126240 5186 126241
rect 4870 126176 4876 126240
rect 4940 126176 4956 126240
rect 5020 126176 5036 126240
rect 5100 126176 5116 126240
rect 5180 126176 5186 126240
rect 4870 126175 5186 126176
rect 106654 126240 106970 126241
rect 106654 126176 106660 126240
rect 106724 126176 106740 126240
rect 106804 126176 106820 126240
rect 106884 126176 106900 126240
rect 106964 126176 106970 126240
rect 106654 126175 106970 126176
rect 4210 125696 4526 125697
rect 4210 125632 4216 125696
rect 4280 125632 4296 125696
rect 4360 125632 4376 125696
rect 4440 125632 4456 125696
rect 4520 125632 4526 125696
rect 4210 125631 4526 125632
rect 105918 125696 106234 125697
rect 105918 125632 105924 125696
rect 105988 125632 106004 125696
rect 106068 125632 106084 125696
rect 106148 125632 106164 125696
rect 106228 125632 106234 125696
rect 105918 125631 106234 125632
rect 4870 125152 5186 125153
rect 4870 125088 4876 125152
rect 4940 125088 4956 125152
rect 5020 125088 5036 125152
rect 5100 125088 5116 125152
rect 5180 125088 5186 125152
rect 4870 125087 5186 125088
rect 106654 125152 106970 125153
rect 106654 125088 106660 125152
rect 106724 125088 106740 125152
rect 106804 125088 106820 125152
rect 106884 125088 106900 125152
rect 106964 125088 106970 125152
rect 106654 125087 106970 125088
rect 4210 124608 4526 124609
rect 4210 124544 4216 124608
rect 4280 124544 4296 124608
rect 4360 124544 4376 124608
rect 4440 124544 4456 124608
rect 4520 124544 4526 124608
rect 4210 124543 4526 124544
rect 105918 124608 106234 124609
rect 105918 124544 105924 124608
rect 105988 124544 106004 124608
rect 106068 124544 106084 124608
rect 106148 124544 106164 124608
rect 106228 124544 106234 124608
rect 105918 124543 106234 124544
rect 4870 124064 5186 124065
rect 4870 124000 4876 124064
rect 4940 124000 4956 124064
rect 5020 124000 5036 124064
rect 5100 124000 5116 124064
rect 5180 124000 5186 124064
rect 4870 123999 5186 124000
rect 106654 124064 106970 124065
rect 106654 124000 106660 124064
rect 106724 124000 106740 124064
rect 106804 124000 106820 124064
rect 106884 124000 106900 124064
rect 106964 124000 106970 124064
rect 106654 123999 106970 124000
rect 4210 123520 4526 123521
rect 4210 123456 4216 123520
rect 4280 123456 4296 123520
rect 4360 123456 4376 123520
rect 4440 123456 4456 123520
rect 4520 123456 4526 123520
rect 4210 123455 4526 123456
rect 105918 123520 106234 123521
rect 105918 123456 105924 123520
rect 105988 123456 106004 123520
rect 106068 123456 106084 123520
rect 106148 123456 106164 123520
rect 106228 123456 106234 123520
rect 105918 123455 106234 123456
rect 4870 122976 5186 122977
rect 4870 122912 4876 122976
rect 4940 122912 4956 122976
rect 5020 122912 5036 122976
rect 5100 122912 5116 122976
rect 5180 122912 5186 122976
rect 4870 122911 5186 122912
rect 106654 122976 106970 122977
rect 106654 122912 106660 122976
rect 106724 122912 106740 122976
rect 106804 122912 106820 122976
rect 106884 122912 106900 122976
rect 106964 122912 106970 122976
rect 106654 122911 106970 122912
rect 4210 122432 4526 122433
rect 4210 122368 4216 122432
rect 4280 122368 4296 122432
rect 4360 122368 4376 122432
rect 4440 122368 4456 122432
rect 4520 122368 4526 122432
rect 4210 122367 4526 122368
rect 105918 122432 106234 122433
rect 105918 122368 105924 122432
rect 105988 122368 106004 122432
rect 106068 122368 106084 122432
rect 106148 122368 106164 122432
rect 106228 122368 106234 122432
rect 105918 122367 106234 122368
rect 4870 121888 5186 121889
rect 4870 121824 4876 121888
rect 4940 121824 4956 121888
rect 5020 121824 5036 121888
rect 5100 121824 5116 121888
rect 5180 121824 5186 121888
rect 4870 121823 5186 121824
rect 106654 121888 106970 121889
rect 106654 121824 106660 121888
rect 106724 121824 106740 121888
rect 106804 121824 106820 121888
rect 106884 121824 106900 121888
rect 106964 121824 106970 121888
rect 106654 121823 106970 121824
rect 4210 121344 4526 121345
rect 4210 121280 4216 121344
rect 4280 121280 4296 121344
rect 4360 121280 4376 121344
rect 4440 121280 4456 121344
rect 4520 121280 4526 121344
rect 4210 121279 4526 121280
rect 105918 121344 106234 121345
rect 105918 121280 105924 121344
rect 105988 121280 106004 121344
rect 106068 121280 106084 121344
rect 106148 121280 106164 121344
rect 106228 121280 106234 121344
rect 105918 121279 106234 121280
rect 4870 120800 5186 120801
rect 4870 120736 4876 120800
rect 4940 120736 4956 120800
rect 5020 120736 5036 120800
rect 5100 120736 5116 120800
rect 5180 120736 5186 120800
rect 4870 120735 5186 120736
rect 106654 120800 106970 120801
rect 106654 120736 106660 120800
rect 106724 120736 106740 120800
rect 106804 120736 106820 120800
rect 106884 120736 106900 120800
rect 106964 120736 106970 120800
rect 106654 120735 106970 120736
rect 4210 120256 4526 120257
rect 4210 120192 4216 120256
rect 4280 120192 4296 120256
rect 4360 120192 4376 120256
rect 4440 120192 4456 120256
rect 4520 120192 4526 120256
rect 4210 120191 4526 120192
rect 105918 120256 106234 120257
rect 105918 120192 105924 120256
rect 105988 120192 106004 120256
rect 106068 120192 106084 120256
rect 106148 120192 106164 120256
rect 106228 120192 106234 120256
rect 105918 120191 106234 120192
rect 4870 119712 5186 119713
rect 4870 119648 4876 119712
rect 4940 119648 4956 119712
rect 5020 119648 5036 119712
rect 5100 119648 5116 119712
rect 5180 119648 5186 119712
rect 4870 119647 5186 119648
rect 106654 119712 106970 119713
rect 106654 119648 106660 119712
rect 106724 119648 106740 119712
rect 106804 119648 106820 119712
rect 106884 119648 106900 119712
rect 106964 119648 106970 119712
rect 106654 119647 106970 119648
rect 4210 119168 4526 119169
rect 4210 119104 4216 119168
rect 4280 119104 4296 119168
rect 4360 119104 4376 119168
rect 4440 119104 4456 119168
rect 4520 119104 4526 119168
rect 4210 119103 4526 119104
rect 105918 119168 106234 119169
rect 105918 119104 105924 119168
rect 105988 119104 106004 119168
rect 106068 119104 106084 119168
rect 106148 119104 106164 119168
rect 106228 119104 106234 119168
rect 105918 119103 106234 119104
rect 4870 118624 5186 118625
rect 4870 118560 4876 118624
rect 4940 118560 4956 118624
rect 5020 118560 5036 118624
rect 5100 118560 5116 118624
rect 5180 118560 5186 118624
rect 4870 118559 5186 118560
rect 106654 118624 106970 118625
rect 106654 118560 106660 118624
rect 106724 118560 106740 118624
rect 106804 118560 106820 118624
rect 106884 118560 106900 118624
rect 106964 118560 106970 118624
rect 106654 118559 106970 118560
rect 4210 118080 4526 118081
rect 4210 118016 4216 118080
rect 4280 118016 4296 118080
rect 4360 118016 4376 118080
rect 4440 118016 4456 118080
rect 4520 118016 4526 118080
rect 4210 118015 4526 118016
rect 105918 118080 106234 118081
rect 105918 118016 105924 118080
rect 105988 118016 106004 118080
rect 106068 118016 106084 118080
rect 106148 118016 106164 118080
rect 106228 118016 106234 118080
rect 105918 118015 106234 118016
rect 4870 117536 5186 117537
rect 4870 117472 4876 117536
rect 4940 117472 4956 117536
rect 5020 117472 5036 117536
rect 5100 117472 5116 117536
rect 5180 117472 5186 117536
rect 4870 117471 5186 117472
rect 106654 117536 106970 117537
rect 106654 117472 106660 117536
rect 106724 117472 106740 117536
rect 106804 117472 106820 117536
rect 106884 117472 106900 117536
rect 106964 117472 106970 117536
rect 106654 117471 106970 117472
rect 4210 116992 4526 116993
rect 4210 116928 4216 116992
rect 4280 116928 4296 116992
rect 4360 116928 4376 116992
rect 4440 116928 4456 116992
rect 4520 116928 4526 116992
rect 4210 116927 4526 116928
rect 105918 116992 106234 116993
rect 105918 116928 105924 116992
rect 105988 116928 106004 116992
rect 106068 116928 106084 116992
rect 106148 116928 106164 116992
rect 106228 116928 106234 116992
rect 105918 116927 106234 116928
rect 4870 116448 5186 116449
rect 4870 116384 4876 116448
rect 4940 116384 4956 116448
rect 5020 116384 5036 116448
rect 5100 116384 5116 116448
rect 5180 116384 5186 116448
rect 4870 116383 5186 116384
rect 106654 116448 106970 116449
rect 106654 116384 106660 116448
rect 106724 116384 106740 116448
rect 106804 116384 106820 116448
rect 106884 116384 106900 116448
rect 106964 116384 106970 116448
rect 106654 116383 106970 116384
rect 4210 115904 4526 115905
rect 4210 115840 4216 115904
rect 4280 115840 4296 115904
rect 4360 115840 4376 115904
rect 4440 115840 4456 115904
rect 4520 115840 4526 115904
rect 4210 115839 4526 115840
rect 105918 115904 106234 115905
rect 105918 115840 105924 115904
rect 105988 115840 106004 115904
rect 106068 115840 106084 115904
rect 106148 115840 106164 115904
rect 106228 115840 106234 115904
rect 105918 115839 106234 115840
rect 4870 115360 5186 115361
rect 4870 115296 4876 115360
rect 4940 115296 4956 115360
rect 5020 115296 5036 115360
rect 5100 115296 5116 115360
rect 5180 115296 5186 115360
rect 4870 115295 5186 115296
rect 106654 115360 106970 115361
rect 106654 115296 106660 115360
rect 106724 115296 106740 115360
rect 106804 115296 106820 115360
rect 106884 115296 106900 115360
rect 106964 115296 106970 115360
rect 106654 115295 106970 115296
rect 4210 114816 4526 114817
rect 4210 114752 4216 114816
rect 4280 114752 4296 114816
rect 4360 114752 4376 114816
rect 4440 114752 4456 114816
rect 4520 114752 4526 114816
rect 4210 114751 4526 114752
rect 105918 114816 106234 114817
rect 105918 114752 105924 114816
rect 105988 114752 106004 114816
rect 106068 114752 106084 114816
rect 106148 114752 106164 114816
rect 106228 114752 106234 114816
rect 105918 114751 106234 114752
rect 4870 114272 5186 114273
rect 4870 114208 4876 114272
rect 4940 114208 4956 114272
rect 5020 114208 5036 114272
rect 5100 114208 5116 114272
rect 5180 114208 5186 114272
rect 4870 114207 5186 114208
rect 106654 114272 106970 114273
rect 106654 114208 106660 114272
rect 106724 114208 106740 114272
rect 106804 114208 106820 114272
rect 106884 114208 106900 114272
rect 106964 114208 106970 114272
rect 106654 114207 106970 114208
rect 4210 113728 4526 113729
rect 4210 113664 4216 113728
rect 4280 113664 4296 113728
rect 4360 113664 4376 113728
rect 4440 113664 4456 113728
rect 4520 113664 4526 113728
rect 4210 113663 4526 113664
rect 105918 113728 106234 113729
rect 105918 113664 105924 113728
rect 105988 113664 106004 113728
rect 106068 113664 106084 113728
rect 106148 113664 106164 113728
rect 106228 113664 106234 113728
rect 105918 113663 106234 113664
rect 4870 113184 5186 113185
rect 4870 113120 4876 113184
rect 4940 113120 4956 113184
rect 5020 113120 5036 113184
rect 5100 113120 5116 113184
rect 5180 113120 5186 113184
rect 4870 113119 5186 113120
rect 106654 113184 106970 113185
rect 106654 113120 106660 113184
rect 106724 113120 106740 113184
rect 106804 113120 106820 113184
rect 106884 113120 106900 113184
rect 106964 113120 106970 113184
rect 106654 113119 106970 113120
rect 4210 112640 4526 112641
rect 4210 112576 4216 112640
rect 4280 112576 4296 112640
rect 4360 112576 4376 112640
rect 4440 112576 4456 112640
rect 4520 112576 4526 112640
rect 4210 112575 4526 112576
rect 105918 112640 106234 112641
rect 105918 112576 105924 112640
rect 105988 112576 106004 112640
rect 106068 112576 106084 112640
rect 106148 112576 106164 112640
rect 106228 112576 106234 112640
rect 105918 112575 106234 112576
rect 4870 112096 5186 112097
rect 4870 112032 4876 112096
rect 4940 112032 4956 112096
rect 5020 112032 5036 112096
rect 5100 112032 5116 112096
rect 5180 112032 5186 112096
rect 4870 112031 5186 112032
rect 106654 112096 106970 112097
rect 106654 112032 106660 112096
rect 106724 112032 106740 112096
rect 106804 112032 106820 112096
rect 106884 112032 106900 112096
rect 106964 112032 106970 112096
rect 106654 112031 106970 112032
rect 4210 111552 4526 111553
rect 4210 111488 4216 111552
rect 4280 111488 4296 111552
rect 4360 111488 4376 111552
rect 4440 111488 4456 111552
rect 4520 111488 4526 111552
rect 4210 111487 4526 111488
rect 105918 111552 106234 111553
rect 105918 111488 105924 111552
rect 105988 111488 106004 111552
rect 106068 111488 106084 111552
rect 106148 111488 106164 111552
rect 106228 111488 106234 111552
rect 105918 111487 106234 111488
rect 9489 111254 9555 111257
rect 9489 111252 10028 111254
rect 9489 111196 9494 111252
rect 9550 111196 10028 111252
rect 9489 111194 10028 111196
rect 9489 111191 9555 111194
rect 4870 111008 5186 111009
rect 0 110938 800 110968
rect 4870 110944 4876 111008
rect 4940 110944 4956 111008
rect 5020 110944 5036 111008
rect 5100 110944 5116 111008
rect 5180 110944 5186 111008
rect 4870 110943 5186 110944
rect 106654 111008 106970 111009
rect 106654 110944 106660 111008
rect 106724 110944 106740 111008
rect 106804 110944 106820 111008
rect 106884 110944 106900 111008
rect 106964 110944 106970 111008
rect 106654 110943 106970 110944
rect 1301 110938 1367 110941
rect 0 110936 1367 110938
rect 0 110880 1306 110936
rect 1362 110880 1367 110936
rect 0 110878 1367 110880
rect 0 110848 800 110878
rect 1301 110875 1367 110878
rect 4210 110464 4526 110465
rect 4210 110400 4216 110464
rect 4280 110400 4296 110464
rect 4360 110400 4376 110464
rect 4440 110400 4456 110464
rect 4520 110400 4526 110464
rect 4210 110399 4526 110400
rect 105918 110464 106234 110465
rect 105918 110400 105924 110464
rect 105988 110400 106004 110464
rect 106068 110400 106084 110464
rect 106148 110400 106164 110464
rect 106228 110400 106234 110464
rect 105918 110399 106234 110400
rect 4870 109920 5186 109921
rect 4870 109856 4876 109920
rect 4940 109856 4956 109920
rect 5020 109856 5036 109920
rect 5100 109856 5116 109920
rect 5180 109856 5186 109920
rect 4870 109855 5186 109856
rect 106654 109920 106970 109921
rect 106654 109856 106660 109920
rect 106724 109856 106740 109920
rect 106804 109856 106820 109920
rect 106884 109856 106900 109920
rect 106964 109856 106970 109920
rect 106654 109855 106970 109856
rect 0 109578 800 109608
rect 1301 109578 1367 109581
rect 0 109576 1367 109578
rect 0 109520 1306 109576
rect 1362 109520 1367 109576
rect 0 109518 1367 109520
rect 0 109488 800 109518
rect 1301 109515 1367 109518
rect 9489 109554 9555 109557
rect 9489 109552 10028 109554
rect 9489 109496 9494 109552
rect 9550 109496 10028 109552
rect 9489 109494 10028 109496
rect 9489 109491 9555 109494
rect 4210 109376 4526 109377
rect 4210 109312 4216 109376
rect 4280 109312 4296 109376
rect 4360 109312 4376 109376
rect 4440 109312 4456 109376
rect 4520 109312 4526 109376
rect 4210 109311 4526 109312
rect 105918 109376 106234 109377
rect 105918 109312 105924 109376
rect 105988 109312 106004 109376
rect 106068 109312 106084 109376
rect 106148 109312 106164 109376
rect 106228 109312 106234 109376
rect 105918 109311 106234 109312
rect 4870 108832 5186 108833
rect 4870 108768 4876 108832
rect 4940 108768 4956 108832
rect 5020 108768 5036 108832
rect 5100 108768 5116 108832
rect 5180 108768 5186 108832
rect 4870 108767 5186 108768
rect 106654 108832 106970 108833
rect 106654 108768 106660 108832
rect 106724 108768 106740 108832
rect 106804 108768 106820 108832
rect 106884 108768 106900 108832
rect 106964 108768 106970 108832
rect 106654 108767 106970 108768
rect 9489 108426 9555 108429
rect 9489 108424 10028 108426
rect 9489 108368 9494 108424
rect 9550 108368 10028 108424
rect 9489 108366 10028 108368
rect 9489 108363 9555 108366
rect 4210 108288 4526 108289
rect 0 108218 800 108248
rect 4210 108224 4216 108288
rect 4280 108224 4296 108288
rect 4360 108224 4376 108288
rect 4440 108224 4456 108288
rect 4520 108224 4526 108288
rect 4210 108223 4526 108224
rect 105918 108288 106234 108289
rect 105918 108224 105924 108288
rect 105988 108224 106004 108288
rect 106068 108224 106084 108288
rect 106148 108224 106164 108288
rect 106228 108224 106234 108288
rect 105918 108223 106234 108224
rect 1301 108218 1367 108221
rect 0 108216 1367 108218
rect 0 108160 1306 108216
rect 1362 108160 1367 108216
rect 0 108158 1367 108160
rect 0 108128 800 108158
rect 1301 108155 1367 108158
rect 4870 107744 5186 107745
rect 4870 107680 4876 107744
rect 4940 107680 4956 107744
rect 5020 107680 5036 107744
rect 5100 107680 5116 107744
rect 5180 107680 5186 107744
rect 4870 107679 5186 107680
rect 106654 107744 106970 107745
rect 106654 107680 106660 107744
rect 106724 107680 106740 107744
rect 106804 107680 106820 107744
rect 106884 107680 106900 107744
rect 106964 107680 106970 107744
rect 106654 107679 106970 107680
rect 4210 107200 4526 107201
rect 4210 107136 4216 107200
rect 4280 107136 4296 107200
rect 4360 107136 4376 107200
rect 4440 107136 4456 107200
rect 4520 107136 4526 107200
rect 4210 107135 4526 107136
rect 105918 107200 106234 107201
rect 105918 107136 105924 107200
rect 105988 107136 106004 107200
rect 106068 107136 106084 107200
rect 106148 107136 106164 107200
rect 106228 107136 106234 107200
rect 105918 107135 106234 107136
rect 0 106858 800 106888
rect 1209 106858 1275 106861
rect 0 106856 1275 106858
rect 0 106800 1214 106856
rect 1270 106800 1275 106856
rect 0 106798 1275 106800
rect 0 106768 800 106798
rect 1209 106795 1275 106798
rect 9489 106726 9555 106729
rect 9489 106724 10028 106726
rect 9489 106668 9494 106724
rect 9550 106668 10028 106724
rect 9489 106666 10028 106668
rect 9489 106663 9555 106666
rect 4870 106656 5186 106657
rect 4870 106592 4876 106656
rect 4940 106592 4956 106656
rect 5020 106592 5036 106656
rect 5100 106592 5116 106656
rect 5180 106592 5186 106656
rect 4870 106591 5186 106592
rect 106654 106656 106970 106657
rect 106654 106592 106660 106656
rect 106724 106592 106740 106656
rect 106804 106592 106820 106656
rect 106884 106592 106900 106656
rect 106964 106592 106970 106656
rect 106654 106591 106970 106592
rect 4210 106112 4526 106113
rect 4210 106048 4216 106112
rect 4280 106048 4296 106112
rect 4360 106048 4376 106112
rect 4440 106048 4456 106112
rect 4520 106048 4526 106112
rect 4210 106047 4526 106048
rect 105918 106112 106234 106113
rect 105918 106048 105924 106112
rect 105988 106048 106004 106112
rect 106068 106048 106084 106112
rect 106148 106048 106164 106112
rect 106228 106048 106234 106112
rect 105918 106047 106234 106048
rect 9489 105643 9555 105646
rect 9489 105641 10028 105643
rect 9489 105585 9494 105641
rect 9550 105585 10028 105641
rect 9489 105583 10028 105585
rect 9489 105580 9555 105583
rect 4870 105568 5186 105569
rect 0 105498 800 105528
rect 4870 105504 4876 105568
rect 4940 105504 4956 105568
rect 5020 105504 5036 105568
rect 5100 105504 5116 105568
rect 5180 105504 5186 105568
rect 4870 105503 5186 105504
rect 106654 105568 106970 105569
rect 106654 105504 106660 105568
rect 106724 105504 106740 105568
rect 106804 105504 106820 105568
rect 106884 105504 106900 105568
rect 106964 105504 106970 105568
rect 106654 105503 106970 105504
rect 1301 105498 1367 105501
rect 0 105496 1367 105498
rect 0 105440 1306 105496
rect 1362 105440 1367 105496
rect 0 105438 1367 105440
rect 0 105408 800 105438
rect 1301 105435 1367 105438
rect 4210 105024 4526 105025
rect 4210 104960 4216 105024
rect 4280 104960 4296 105024
rect 4360 104960 4376 105024
rect 4440 104960 4456 105024
rect 4520 104960 4526 105024
rect 4210 104959 4526 104960
rect 105918 105024 106234 105025
rect 105918 104960 105924 105024
rect 105988 104960 106004 105024
rect 106068 104960 106084 105024
rect 106148 104960 106164 105024
rect 106228 104960 106234 105024
rect 105918 104959 106234 104960
rect 4870 104480 5186 104481
rect 4870 104416 4876 104480
rect 4940 104416 4956 104480
rect 5020 104416 5036 104480
rect 5100 104416 5116 104480
rect 5180 104416 5186 104480
rect 4870 104415 5186 104416
rect 106654 104480 106970 104481
rect 106654 104416 106660 104480
rect 106724 104416 106740 104480
rect 106804 104416 106820 104480
rect 106884 104416 106900 104480
rect 106964 104416 106970 104480
rect 106654 104415 106970 104416
rect 0 104138 800 104168
rect 1301 104138 1367 104141
rect 0 104136 1367 104138
rect 0 104080 1306 104136
rect 1362 104080 1367 104136
rect 0 104078 1367 104080
rect 0 104048 800 104078
rect 1301 104075 1367 104078
rect 9489 103963 9555 103966
rect 9489 103961 10028 103963
rect 4210 103936 4526 103937
rect 4210 103872 4216 103936
rect 4280 103872 4296 103936
rect 4360 103872 4376 103936
rect 4440 103872 4456 103936
rect 4520 103872 4526 103936
rect 9489 103905 9494 103961
rect 9550 103905 10028 103961
rect 9489 103903 10028 103905
rect 105918 103936 106234 103937
rect 9489 103900 9555 103903
rect 4210 103871 4526 103872
rect 105918 103872 105924 103936
rect 105988 103872 106004 103936
rect 106068 103872 106084 103936
rect 106148 103872 106164 103936
rect 106228 103872 106234 103936
rect 105918 103871 106234 103872
rect 4870 103392 5186 103393
rect 4870 103328 4876 103392
rect 4940 103328 4956 103392
rect 5020 103328 5036 103392
rect 5100 103328 5116 103392
rect 5180 103328 5186 103392
rect 4870 103327 5186 103328
rect 106654 103392 106970 103393
rect 106654 103328 106660 103392
rect 106724 103328 106740 103392
rect 106804 103328 106820 103392
rect 106884 103328 106900 103392
rect 106964 103328 106970 103392
rect 106654 103327 106970 103328
rect 4210 102848 4526 102849
rect 4210 102784 4216 102848
rect 4280 102784 4296 102848
rect 4360 102784 4376 102848
rect 4440 102784 4456 102848
rect 4520 102784 4526 102848
rect 4210 102783 4526 102784
rect 105918 102848 106234 102849
rect 105918 102784 105924 102848
rect 105988 102784 106004 102848
rect 106068 102784 106084 102848
rect 106148 102784 106164 102848
rect 106228 102784 106234 102848
rect 105918 102783 106234 102784
rect 4870 102304 5186 102305
rect 4870 102240 4876 102304
rect 4940 102240 4956 102304
rect 5020 102240 5036 102304
rect 5100 102240 5116 102304
rect 5180 102240 5186 102304
rect 4870 102239 5186 102240
rect 106654 102304 106970 102305
rect 106654 102240 106660 102304
rect 106724 102240 106740 102304
rect 106804 102240 106820 102304
rect 106884 102240 106900 102304
rect 106964 102240 106970 102304
rect 106654 102239 106970 102240
rect 4210 101760 4526 101761
rect 4210 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4526 101760
rect 4210 101695 4526 101696
rect 105918 101760 106234 101761
rect 105918 101696 105924 101760
rect 105988 101696 106004 101760
rect 106068 101696 106084 101760
rect 106148 101696 106164 101760
rect 106228 101696 106234 101760
rect 105918 101695 106234 101696
rect 4870 101216 5186 101217
rect 4870 101152 4876 101216
rect 4940 101152 4956 101216
rect 5020 101152 5036 101216
rect 5100 101152 5116 101216
rect 5180 101152 5186 101216
rect 4870 101151 5186 101152
rect 106654 101216 106970 101217
rect 106654 101152 106660 101216
rect 106724 101152 106740 101216
rect 106804 101152 106820 101216
rect 106884 101152 106900 101216
rect 106964 101152 106970 101216
rect 106654 101151 106970 101152
rect 4210 100672 4526 100673
rect 4210 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4526 100672
rect 4210 100607 4526 100608
rect 105918 100672 106234 100673
rect 105918 100608 105924 100672
rect 105988 100608 106004 100672
rect 106068 100608 106084 100672
rect 106148 100608 106164 100672
rect 106228 100608 106234 100672
rect 105918 100607 106234 100608
rect 4870 100128 5186 100129
rect 4870 100064 4876 100128
rect 4940 100064 4956 100128
rect 5020 100064 5036 100128
rect 5100 100064 5116 100128
rect 5180 100064 5186 100128
rect 4870 100063 5186 100064
rect 106654 100128 106970 100129
rect 106654 100064 106660 100128
rect 106724 100064 106740 100128
rect 106804 100064 106820 100128
rect 106884 100064 106900 100128
rect 106964 100064 106970 100128
rect 106654 100063 106970 100064
rect 4210 99584 4526 99585
rect 4210 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4526 99584
rect 4210 99519 4526 99520
rect 105918 99584 106234 99585
rect 105918 99520 105924 99584
rect 105988 99520 106004 99584
rect 106068 99520 106084 99584
rect 106148 99520 106164 99584
rect 106228 99520 106234 99584
rect 105918 99519 106234 99520
rect 4870 99040 5186 99041
rect 4870 98976 4876 99040
rect 4940 98976 4956 99040
rect 5020 98976 5036 99040
rect 5100 98976 5116 99040
rect 5180 98976 5186 99040
rect 4870 98975 5186 98976
rect 106654 99040 106970 99041
rect 106654 98976 106660 99040
rect 106724 98976 106740 99040
rect 106804 98976 106820 99040
rect 106884 98976 106900 99040
rect 106964 98976 106970 99040
rect 106654 98975 106970 98976
rect 4210 98496 4526 98497
rect 4210 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4526 98496
rect 4210 98431 4526 98432
rect 105918 98496 106234 98497
rect 105918 98432 105924 98496
rect 105988 98432 106004 98496
rect 106068 98432 106084 98496
rect 106148 98432 106164 98496
rect 106228 98432 106234 98496
rect 105918 98431 106234 98432
rect 4870 97952 5186 97953
rect 4870 97888 4876 97952
rect 4940 97888 4956 97952
rect 5020 97888 5036 97952
rect 5100 97888 5116 97952
rect 5180 97888 5186 97952
rect 4870 97887 5186 97888
rect 106654 97952 106970 97953
rect 106654 97888 106660 97952
rect 106724 97888 106740 97952
rect 106804 97888 106820 97952
rect 106884 97888 106900 97952
rect 106964 97888 106970 97952
rect 106654 97887 106970 97888
rect 4210 97408 4526 97409
rect 4210 97344 4216 97408
rect 4280 97344 4296 97408
rect 4360 97344 4376 97408
rect 4440 97344 4456 97408
rect 4520 97344 4526 97408
rect 4210 97343 4526 97344
rect 105918 97408 106234 97409
rect 105918 97344 105924 97408
rect 105988 97344 106004 97408
rect 106068 97344 106084 97408
rect 106148 97344 106164 97408
rect 106228 97344 106234 97408
rect 105918 97343 106234 97344
rect 4870 96864 5186 96865
rect 4870 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5186 96864
rect 4870 96799 5186 96800
rect 106654 96864 106970 96865
rect 106654 96800 106660 96864
rect 106724 96800 106740 96864
rect 106804 96800 106820 96864
rect 106884 96800 106900 96864
rect 106964 96800 106970 96864
rect 106654 96799 106970 96800
rect 4210 96320 4526 96321
rect 4210 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4526 96320
rect 4210 96255 4526 96256
rect 105918 96320 106234 96321
rect 105918 96256 105924 96320
rect 105988 96256 106004 96320
rect 106068 96256 106084 96320
rect 106148 96256 106164 96320
rect 106228 96256 106234 96320
rect 105918 96255 106234 96256
rect 4870 95776 5186 95777
rect 4870 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5186 95776
rect 4870 95711 5186 95712
rect 106654 95776 106970 95777
rect 106654 95712 106660 95776
rect 106724 95712 106740 95776
rect 106804 95712 106820 95776
rect 106884 95712 106900 95776
rect 106964 95712 106970 95776
rect 106654 95711 106970 95712
rect 4210 95232 4526 95233
rect 4210 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4526 95232
rect 4210 95167 4526 95168
rect 105918 95232 106234 95233
rect 105918 95168 105924 95232
rect 105988 95168 106004 95232
rect 106068 95168 106084 95232
rect 106148 95168 106164 95232
rect 106228 95168 106234 95232
rect 105918 95167 106234 95168
rect 102501 95090 102567 95093
rect 101948 95088 102567 95090
rect 101948 95032 102506 95088
rect 102562 95032 102567 95088
rect 101948 95030 102567 95032
rect 102501 95027 102567 95030
rect 4870 94688 5186 94689
rect 4870 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5186 94688
rect 4870 94623 5186 94624
rect 106654 94688 106970 94689
rect 106654 94624 106660 94688
rect 106724 94624 106740 94688
rect 106804 94624 106820 94688
rect 106884 94624 106900 94688
rect 106964 94624 106970 94688
rect 106654 94623 106970 94624
rect 4210 94144 4526 94145
rect 4210 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4526 94144
rect 4210 94079 4526 94080
rect 105918 94144 106234 94145
rect 105918 94080 105924 94144
rect 105988 94080 106004 94144
rect 106068 94080 106084 94144
rect 106148 94080 106164 94144
rect 106228 94080 106234 94144
rect 105918 94079 106234 94080
rect 4870 93600 5186 93601
rect 4870 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5186 93600
rect 4870 93535 5186 93536
rect 106654 93600 106970 93601
rect 106654 93536 106660 93600
rect 106724 93536 106740 93600
rect 106804 93536 106820 93600
rect 106884 93536 106900 93600
rect 106964 93536 106970 93600
rect 106654 93535 106970 93536
rect 102174 93390 102180 93392
rect 101948 93330 102180 93390
rect 102174 93328 102180 93330
rect 102244 93390 102250 93392
rect 102409 93390 102475 93393
rect 102244 93388 102475 93390
rect 102244 93332 102414 93388
rect 102470 93332 102475 93388
rect 102244 93330 102475 93332
rect 102244 93328 102250 93330
rect 102409 93327 102475 93330
rect 4210 93056 4526 93057
rect 4210 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4526 93056
rect 4210 92991 4526 92992
rect 105918 93056 106234 93057
rect 105918 92992 105924 93056
rect 105988 92992 106004 93056
rect 106068 92992 106084 93056
rect 106148 92992 106164 93056
rect 106228 92992 106234 93056
rect 105918 92991 106234 92992
rect 4870 92512 5186 92513
rect 4870 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5186 92512
rect 4870 92447 5186 92448
rect 106654 92512 106970 92513
rect 106654 92448 106660 92512
rect 106724 92448 106740 92512
rect 106804 92448 106820 92512
rect 106884 92448 106900 92512
rect 106964 92448 106970 92512
rect 106654 92447 106970 92448
rect 103881 92306 103947 92309
rect 102550 92304 103947 92306
rect 102041 92262 102107 92265
rect 102550 92262 103886 92304
rect 101948 92260 103886 92262
rect 101948 92204 102046 92260
rect 102102 92248 103886 92260
rect 103942 92248 103947 92304
rect 102102 92246 103947 92248
rect 102102 92204 102610 92246
rect 103881 92243 103947 92246
rect 101948 92202 102610 92204
rect 102041 92199 102107 92202
rect 4210 91968 4526 91969
rect 4210 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4526 91968
rect 4210 91903 4526 91904
rect 105918 91968 106234 91969
rect 105918 91904 105924 91968
rect 105988 91904 106004 91968
rect 106068 91904 106084 91968
rect 106148 91904 106164 91968
rect 106228 91904 106234 91968
rect 105918 91903 106234 91904
rect 4870 91424 5186 91425
rect 4870 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5186 91424
rect 4870 91359 5186 91360
rect 106654 91424 106970 91425
rect 106654 91360 106660 91424
rect 106724 91360 106740 91424
rect 106804 91360 106820 91424
rect 106884 91360 106900 91424
rect 106964 91360 106970 91424
rect 106654 91359 106970 91360
rect 4210 90880 4526 90881
rect 4210 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4526 90880
rect 4210 90815 4526 90816
rect 105918 90880 106234 90881
rect 105918 90816 105924 90880
rect 105988 90816 106004 90880
rect 106068 90816 106084 90880
rect 106148 90816 106164 90880
rect 106228 90816 106234 90880
rect 105918 90815 106234 90816
rect 4870 90336 5186 90337
rect 4870 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5186 90336
rect 4870 90271 5186 90272
rect 106654 90336 106970 90337
rect 106654 90272 106660 90336
rect 106724 90272 106740 90336
rect 106804 90272 106820 90336
rect 106884 90272 106900 90336
rect 106964 90272 106970 90336
rect 106654 90271 106970 90272
rect 4210 89792 4526 89793
rect 4210 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4526 89792
rect 4210 89727 4526 89728
rect 105918 89792 106234 89793
rect 105918 89728 105924 89792
rect 105988 89728 106004 89792
rect 106068 89728 106084 89792
rect 106148 89728 106164 89792
rect 106228 89728 106234 89792
rect 105918 89727 106234 89728
rect 4870 89248 5186 89249
rect 4870 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5186 89248
rect 4870 89183 5186 89184
rect 106654 89248 106970 89249
rect 106654 89184 106660 89248
rect 106724 89184 106740 89248
rect 106804 89184 106820 89248
rect 106884 89184 106900 89248
rect 106964 89184 106970 89248
rect 106654 89183 106970 89184
rect 4210 88704 4526 88705
rect 4210 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4526 88704
rect 4210 88639 4526 88640
rect 105918 88704 106234 88705
rect 105918 88640 105924 88704
rect 105988 88640 106004 88704
rect 106068 88640 106084 88704
rect 106148 88640 106164 88704
rect 106228 88640 106234 88704
rect 105918 88639 106234 88640
rect 0 88498 800 88528
rect 1301 88498 1367 88501
rect 0 88496 1367 88498
rect 0 88440 1306 88496
rect 1362 88440 1367 88496
rect 0 88438 1367 88440
rect 0 88408 800 88438
rect 1301 88435 1367 88438
rect 4870 88160 5186 88161
rect 4870 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5186 88160
rect 4870 88095 5186 88096
rect 106654 88160 106970 88161
rect 106654 88096 106660 88160
rect 106724 88096 106740 88160
rect 106804 88096 106820 88160
rect 106884 88096 106900 88160
rect 106964 88096 106970 88160
rect 106654 88095 106970 88096
rect 0 87818 800 87848
rect 1209 87818 1275 87821
rect 0 87816 1275 87818
rect 0 87760 1214 87816
rect 1270 87760 1275 87816
rect 0 87758 1275 87760
rect 0 87728 800 87758
rect 1209 87755 1275 87758
rect 4210 87616 4526 87617
rect 4210 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4526 87616
rect 4210 87551 4526 87552
rect 105918 87616 106234 87617
rect 105918 87552 105924 87616
rect 105988 87552 106004 87616
rect 106068 87552 106084 87616
rect 106148 87552 106164 87616
rect 106228 87552 106234 87616
rect 105918 87551 106234 87552
rect 0 87138 800 87168
rect 1209 87138 1275 87141
rect 0 87136 1275 87138
rect 0 87080 1214 87136
rect 1270 87080 1275 87136
rect 0 87078 1275 87080
rect 0 87048 800 87078
rect 1209 87075 1275 87078
rect 4870 87072 5186 87073
rect 4870 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5186 87072
rect 4870 87007 5186 87008
rect 106654 87072 106970 87073
rect 106654 87008 106660 87072
rect 106724 87008 106740 87072
rect 106804 87008 106820 87072
rect 106884 87008 106900 87072
rect 106964 87008 106970 87072
rect 106654 87007 106970 87008
rect 4210 86528 4526 86529
rect 0 86458 800 86488
rect 4210 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4526 86528
rect 4210 86463 4526 86464
rect 105918 86528 106234 86529
rect 105918 86464 105924 86528
rect 105988 86464 106004 86528
rect 106068 86464 106084 86528
rect 106148 86464 106164 86528
rect 106228 86464 106234 86528
rect 105918 86463 106234 86464
rect 1301 86458 1367 86461
rect 0 86456 1367 86458
rect 0 86400 1306 86456
rect 1362 86400 1367 86456
rect 0 86398 1367 86400
rect 0 86368 800 86398
rect 1301 86395 1367 86398
rect 4870 85984 5186 85985
rect 4870 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5186 85984
rect 4870 85919 5186 85920
rect 106654 85984 106970 85985
rect 106654 85920 106660 85984
rect 106724 85920 106740 85984
rect 106804 85920 106820 85984
rect 106884 85920 106900 85984
rect 106964 85920 106970 85984
rect 106654 85919 106970 85920
rect 0 85778 800 85808
rect 1301 85778 1367 85781
rect 0 85776 1367 85778
rect 0 85720 1306 85776
rect 1362 85720 1367 85776
rect 0 85718 1367 85720
rect 0 85688 800 85718
rect 1301 85715 1367 85718
rect 5533 85506 5599 85509
rect 5533 85504 9506 85506
rect 5533 85448 5538 85504
rect 5594 85483 9506 85504
rect 5594 85448 10028 85483
rect 5533 85446 10028 85448
rect 5533 85443 5599 85446
rect 4210 85440 4526 85441
rect 4210 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4526 85440
rect 9446 85423 10028 85446
rect 105918 85440 106234 85441
rect 4210 85375 4526 85376
rect 105918 85376 105924 85440
rect 105988 85376 106004 85440
rect 106068 85376 106084 85440
rect 106148 85376 106164 85440
rect 106228 85376 106234 85440
rect 105918 85375 106234 85376
rect 0 85098 800 85128
rect 1209 85098 1275 85101
rect 0 85096 1275 85098
rect 0 85040 1214 85096
rect 1270 85040 1275 85096
rect 0 85038 1275 85040
rect 0 85008 800 85038
rect 1209 85035 1275 85038
rect 4870 84896 5186 84897
rect 4870 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5186 84896
rect 4870 84831 5186 84832
rect 106654 84896 106970 84897
rect 106654 84832 106660 84896
rect 106724 84832 106740 84896
rect 106804 84832 106820 84896
rect 106884 84832 106900 84896
rect 106964 84832 106970 84896
rect 106654 84831 106970 84832
rect 0 84418 800 84448
rect 1301 84418 1367 84421
rect 0 84416 1367 84418
rect 0 84360 1306 84416
rect 1362 84360 1367 84416
rect 0 84358 1367 84360
rect 0 84328 800 84358
rect 1301 84355 1367 84358
rect 4210 84352 4526 84353
rect 4210 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4526 84352
rect 4210 84287 4526 84288
rect 105918 84352 106234 84353
rect 105918 84288 105924 84352
rect 105988 84288 106004 84352
rect 106068 84288 106084 84352
rect 106148 84288 106164 84352
rect 106228 84288 106234 84352
rect 105918 84287 106234 84288
rect 4870 83808 5186 83809
rect 0 83738 800 83768
rect 4870 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5186 83808
rect 4870 83743 5186 83744
rect 106654 83808 106970 83809
rect 106654 83744 106660 83808
rect 106724 83744 106740 83808
rect 106804 83744 106820 83808
rect 106884 83744 106900 83808
rect 106964 83744 106970 83808
rect 106654 83743 106970 83744
rect 1301 83738 1367 83741
rect 0 83736 1367 83738
rect 0 83680 1306 83736
rect 1362 83680 1367 83736
rect 0 83678 1367 83680
rect 0 83648 800 83678
rect 1301 83675 1367 83678
rect 4210 83264 4526 83265
rect 4210 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4526 83264
rect 4210 83199 4526 83200
rect 105918 83264 106234 83265
rect 105918 83200 105924 83264
rect 105988 83200 106004 83264
rect 106068 83200 106084 83264
rect 106148 83200 106164 83264
rect 106228 83200 106234 83264
rect 105918 83199 106234 83200
rect 0 83058 800 83088
rect 1301 83058 1367 83061
rect 0 83056 1367 83058
rect 0 83000 1306 83056
rect 1362 83000 1367 83056
rect 0 82998 1367 83000
rect 0 82968 800 82998
rect 1301 82995 1367 82998
rect 4870 82720 5186 82721
rect 4870 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5186 82720
rect 4870 82655 5186 82656
rect 106654 82720 106970 82721
rect 106654 82656 106660 82720
rect 106724 82656 106740 82720
rect 106804 82656 106820 82720
rect 106884 82656 106900 82720
rect 106964 82656 106970 82720
rect 106654 82655 106970 82656
rect 0 82378 800 82408
rect 1209 82378 1275 82381
rect 0 82376 1275 82378
rect 0 82320 1214 82376
rect 1270 82320 1275 82376
rect 0 82318 1275 82320
rect 0 82288 800 82318
rect 1209 82315 1275 82318
rect 4210 82176 4526 82177
rect 4210 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4526 82176
rect 4210 82111 4526 82112
rect 105918 82176 106234 82177
rect 105918 82112 105924 82176
rect 105988 82112 106004 82176
rect 106068 82112 106084 82176
rect 106148 82112 106164 82176
rect 106228 82112 106234 82176
rect 105918 82111 106234 82112
rect 0 81698 800 81728
rect 1209 81698 1275 81701
rect 0 81696 1275 81698
rect 0 81640 1214 81696
rect 1270 81640 1275 81696
rect 0 81638 1275 81640
rect 0 81608 800 81638
rect 1209 81635 1275 81638
rect 4870 81632 5186 81633
rect 4870 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5186 81632
rect 4870 81567 5186 81568
rect 106654 81632 106970 81633
rect 106654 81568 106660 81632
rect 106724 81568 106740 81632
rect 106804 81568 106820 81632
rect 106884 81568 106900 81632
rect 106964 81568 106970 81632
rect 106654 81567 106970 81568
rect 4210 81088 4526 81089
rect 0 81018 800 81048
rect 4210 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4526 81088
rect 4210 81023 4526 81024
rect 105918 81088 106234 81089
rect 105918 81024 105924 81088
rect 105988 81024 106004 81088
rect 106068 81024 106084 81088
rect 106148 81024 106164 81088
rect 106228 81024 106234 81088
rect 105918 81023 106234 81024
rect 1301 81018 1367 81021
rect 0 81016 1367 81018
rect 0 80960 1306 81016
rect 1362 80960 1367 81016
rect 0 80958 1367 80960
rect 0 80928 800 80958
rect 1301 80955 1367 80958
rect 4870 80544 5186 80545
rect 4870 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5186 80544
rect 4870 80479 5186 80480
rect 106654 80544 106970 80545
rect 106654 80480 106660 80544
rect 106724 80480 106740 80544
rect 106804 80480 106820 80544
rect 106884 80480 106900 80544
rect 106964 80480 106970 80544
rect 106654 80479 106970 80480
rect 0 80338 800 80368
rect 1301 80338 1367 80341
rect 0 80336 1367 80338
rect 0 80280 1306 80336
rect 1362 80280 1367 80336
rect 0 80278 1367 80280
rect 0 80248 800 80278
rect 1301 80275 1367 80278
rect 108481 80338 108547 80341
rect 109200 80338 110000 80368
rect 108481 80336 110000 80338
rect 108481 80280 108486 80336
rect 108542 80280 110000 80336
rect 108481 80278 110000 80280
rect 108481 80275 108547 80278
rect 109200 80248 110000 80278
rect 4210 80000 4526 80001
rect 4210 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4526 80000
rect 4210 79935 4526 79936
rect 105918 80000 106234 80001
rect 105918 79936 105924 80000
rect 105988 79936 106004 80000
rect 106068 79936 106084 80000
rect 106148 79936 106164 80000
rect 106228 79936 106234 80000
rect 105918 79935 106234 79936
rect 7465 79930 7531 79933
rect 16113 79932 16179 79933
rect 23473 79932 23539 79933
rect 16062 79930 16068 79932
rect 7465 79928 16068 79930
rect 16132 79928 16179 79932
rect 23432 79930 23438 79932
rect 7465 79872 7470 79928
rect 7526 79872 16068 79928
rect 16174 79872 16179 79928
rect 7465 79870 16068 79872
rect 7465 79867 7531 79870
rect 16062 79868 16068 79870
rect 16132 79868 16179 79872
rect 23382 79870 23438 79930
rect 23502 79928 23539 79932
rect 23534 79872 23539 79928
rect 23432 79868 23438 79870
rect 23502 79868 23539 79872
rect 16113 79867 16179 79868
rect 23473 79867 23539 79868
rect 36261 79932 36327 79933
rect 39757 79932 39823 79933
rect 40953 79932 41019 79933
rect 43253 79932 43319 79933
rect 36261 79928 36286 79932
rect 36350 79930 36356 79932
rect 36261 79872 36266 79928
rect 36261 79868 36286 79872
rect 36350 79870 36418 79930
rect 39757 79928 39790 79932
rect 39854 79930 39860 79932
rect 39757 79872 39762 79928
rect 36350 79868 36356 79870
rect 39757 79868 39790 79872
rect 39854 79870 39914 79930
rect 39854 79868 39860 79870
rect 40952 79868 40958 79932
rect 41022 79930 41028 79932
rect 41022 79870 41110 79930
rect 43253 79928 43294 79932
rect 43358 79930 43364 79932
rect 43253 79872 43258 79928
rect 41022 79868 41028 79870
rect 43253 79868 43294 79872
rect 43358 79870 43410 79930
rect 43358 79868 43364 79870
rect 36261 79867 36327 79868
rect 39757 79867 39823 79868
rect 40953 79867 41019 79868
rect 43253 79867 43319 79868
rect 9581 79794 9647 79797
rect 38653 79796 38719 79797
rect 32776 79794 32782 79796
rect 9581 79792 32782 79794
rect 9581 79736 9586 79792
rect 9642 79736 32782 79792
rect 9581 79734 32782 79736
rect 9581 79731 9647 79734
rect 32776 79732 32782 79734
rect 32846 79732 32852 79796
rect 38616 79794 38622 79796
rect 38562 79734 38622 79794
rect 38686 79792 38719 79796
rect 38714 79736 38719 79792
rect 38616 79732 38622 79734
rect 38686 79732 38719 79736
rect 38653 79731 38719 79732
rect 0 79658 800 79688
rect 1209 79658 1275 79661
rect 0 79656 1275 79658
rect 0 79600 1214 79656
rect 1270 79600 1275 79656
rect 0 79598 1275 79600
rect 0 79568 800 79598
rect 1209 79595 1275 79598
rect 8385 79658 8451 79661
rect 30465 79660 30531 79661
rect 31661 79660 31727 79661
rect 37457 79660 37523 79661
rect 30440 79658 30446 79660
rect 8385 79656 30446 79658
rect 30510 79658 30531 79660
rect 31610 79658 31616 79660
rect 30510 79656 30638 79658
rect 8385 79600 8390 79656
rect 8446 79600 30446 79656
rect 30526 79600 30638 79656
rect 8385 79598 30446 79600
rect 8385 79595 8451 79598
rect 30440 79596 30446 79598
rect 30510 79598 30638 79600
rect 31570 79598 31616 79658
rect 31680 79656 31727 79660
rect 37448 79658 37454 79660
rect 31722 79600 31727 79656
rect 30510 79596 30531 79598
rect 31610 79596 31616 79598
rect 31680 79596 31727 79600
rect 37366 79598 37454 79658
rect 37448 79596 37454 79598
rect 37518 79596 37524 79660
rect 108389 79658 108455 79661
rect 109200 79658 110000 79688
rect 108389 79656 110000 79658
rect 108389 79600 108394 79656
rect 108450 79600 110000 79656
rect 108389 79598 110000 79600
rect 30465 79595 30531 79596
rect 31661 79595 31727 79596
rect 37457 79595 37523 79596
rect 108389 79595 108455 79598
rect 109200 79568 110000 79598
rect 5533 79522 5599 79525
rect 24669 79524 24735 79525
rect 24618 79522 24624 79524
rect 5533 79520 24624 79522
rect 24688 79520 24735 79524
rect 5533 79464 5538 79520
rect 5594 79464 24624 79520
rect 24730 79464 24735 79520
rect 5533 79462 24624 79464
rect 5533 79459 5599 79462
rect 24618 79460 24624 79462
rect 24688 79460 24735 79464
rect 25768 79460 25774 79524
rect 25838 79522 25844 79524
rect 26049 79522 26115 79525
rect 26969 79524 27035 79525
rect 28165 79524 28231 79525
rect 26936 79522 26942 79524
rect 25838 79520 26115 79522
rect 25838 79464 26054 79520
rect 26110 79464 26115 79520
rect 25838 79462 26115 79464
rect 26878 79462 26942 79522
rect 27006 79520 27035 79524
rect 28114 79522 28120 79524
rect 27030 79464 27035 79520
rect 25838 79460 25844 79462
rect 24669 79459 24735 79460
rect 26049 79459 26115 79462
rect 26936 79460 26942 79462
rect 27006 79460 27035 79464
rect 28074 79462 28120 79522
rect 28184 79520 28231 79524
rect 28226 79464 28231 79520
rect 28114 79460 28120 79462
rect 28184 79460 28231 79464
rect 29272 79460 29278 79524
rect 29342 79522 29348 79524
rect 29545 79522 29611 79525
rect 33961 79524 34027 79525
rect 33944 79522 33950 79524
rect 29342 79520 29611 79522
rect 29342 79464 29550 79520
rect 29606 79464 29611 79520
rect 29342 79462 29611 79464
rect 33870 79462 33950 79522
rect 34014 79520 34027 79524
rect 34022 79464 34027 79520
rect 29342 79460 29348 79462
rect 26969 79459 27035 79460
rect 28165 79459 28231 79460
rect 29545 79459 29611 79462
rect 33944 79460 33950 79462
rect 34014 79460 34027 79464
rect 35112 79460 35118 79524
rect 35182 79522 35188 79524
rect 35341 79522 35407 79525
rect 42149 79524 42215 79525
rect 42120 79522 42126 79524
rect 35182 79520 35407 79522
rect 35182 79464 35346 79520
rect 35402 79464 35407 79520
rect 35182 79462 35407 79464
rect 42058 79462 42126 79522
rect 42190 79520 42215 79524
rect 42210 79464 42215 79520
rect 35182 79460 35188 79462
rect 33961 79459 34027 79460
rect 35341 79459 35407 79462
rect 42120 79460 42126 79462
rect 42190 79460 42215 79464
rect 42149 79459 42215 79460
rect 4870 79456 5186 79457
rect 4870 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5186 79456
rect 4870 79391 5186 79392
rect 106654 79456 106970 79457
rect 106654 79392 106660 79456
rect 106724 79392 106740 79456
rect 106804 79392 106820 79456
rect 106884 79392 106900 79456
rect 106964 79392 106970 79456
rect 106654 79391 106970 79392
rect 9305 79250 9371 79253
rect 26969 79250 27035 79253
rect 9305 79248 27035 79250
rect 9305 79192 9310 79248
rect 9366 79192 26974 79248
rect 27030 79192 27035 79248
rect 9305 79190 27035 79192
rect 9305 79187 9371 79190
rect 26969 79187 27035 79190
rect 9213 79114 9279 79117
rect 28165 79114 28231 79117
rect 32857 79116 32923 79117
rect 32806 79114 32812 79116
rect 9213 79112 28231 79114
rect 9213 79056 9218 79112
rect 9274 79056 28170 79112
rect 28226 79056 28231 79112
rect 9213 79054 28231 79056
rect 32766 79054 32812 79114
rect 32876 79112 32923 79116
rect 32918 79056 32923 79112
rect 9213 79051 9279 79054
rect 28165 79051 28231 79054
rect 32806 79052 32812 79054
rect 32876 79052 32923 79056
rect 32857 79051 32923 79052
rect 0 78978 800 79008
rect 1301 78978 1367 78981
rect 0 78976 1367 78978
rect 0 78920 1306 78976
rect 1362 78920 1367 78976
rect 0 78918 1367 78920
rect 0 78888 800 78918
rect 1301 78915 1367 78918
rect 108389 78978 108455 78981
rect 109200 78978 110000 79008
rect 108389 78976 110000 78978
rect 108389 78920 108394 78976
rect 108450 78920 110000 78976
rect 108389 78918 110000 78920
rect 108389 78915 108455 78918
rect 4210 78912 4526 78913
rect 4210 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4526 78912
rect 4210 78847 4526 78848
rect 105918 78912 106234 78913
rect 105918 78848 105924 78912
rect 105988 78848 106004 78912
rect 106068 78848 106084 78912
rect 106148 78848 106164 78912
rect 106228 78848 106234 78912
rect 109200 78888 110000 78918
rect 105918 78847 106234 78848
rect 4870 78368 5186 78369
rect 0 78298 800 78328
rect 4870 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5186 78368
rect 4870 78303 5186 78304
rect 106654 78368 106970 78369
rect 106654 78304 106660 78368
rect 106724 78304 106740 78368
rect 106804 78304 106820 78368
rect 106884 78304 106900 78368
rect 106964 78304 106970 78368
rect 106654 78303 106970 78304
rect 1301 78298 1367 78301
rect 0 78296 1367 78298
rect 0 78240 1306 78296
rect 1362 78240 1367 78296
rect 0 78238 1367 78240
rect 0 78208 800 78238
rect 1301 78235 1367 78238
rect 108389 78298 108455 78301
rect 109200 78298 110000 78328
rect 108389 78296 110000 78298
rect 108389 78240 108394 78296
rect 108450 78240 110000 78296
rect 108389 78238 110000 78240
rect 108389 78235 108455 78238
rect 109200 78208 110000 78238
rect 4210 77824 4526 77825
rect 4210 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4526 77824
rect 4210 77759 4526 77760
rect 34930 77824 35246 77825
rect 34930 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35246 77824
rect 34930 77759 35246 77760
rect 65650 77824 65966 77825
rect 65650 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65966 77824
rect 65650 77759 65966 77760
rect 96370 77824 96686 77825
rect 96370 77760 96376 77824
rect 96440 77760 96456 77824
rect 96520 77760 96536 77824
rect 96600 77760 96616 77824
rect 96680 77760 96686 77824
rect 96370 77759 96686 77760
rect 105918 77824 106234 77825
rect 105918 77760 105924 77824
rect 105988 77760 106004 77824
rect 106068 77760 106084 77824
rect 106148 77760 106164 77824
rect 106228 77760 106234 77824
rect 105918 77759 106234 77760
rect 90398 77692 90404 77756
rect 90468 77754 90474 77756
rect 91461 77754 91527 77757
rect 90468 77752 91527 77754
rect 90468 77696 91466 77752
rect 91522 77696 91527 77752
rect 90468 77694 91527 77696
rect 90468 77692 90474 77694
rect 91461 77691 91527 77694
rect 0 77618 800 77648
rect 1301 77618 1367 77621
rect 0 77616 1367 77618
rect 0 77560 1306 77616
rect 1362 77560 1367 77616
rect 0 77558 1367 77560
rect 0 77528 800 77558
rect 1301 77555 1367 77558
rect 90950 77556 90956 77620
rect 91020 77618 91026 77620
rect 92197 77618 92263 77621
rect 91020 77616 92263 77618
rect 91020 77560 92202 77616
rect 92258 77560 92263 77616
rect 91020 77558 92263 77560
rect 91020 77556 91026 77558
rect 92197 77555 92263 77558
rect 108389 77618 108455 77621
rect 109200 77618 110000 77648
rect 108389 77616 110000 77618
rect 108389 77560 108394 77616
rect 108450 77560 110000 77616
rect 108389 77558 110000 77560
rect 108389 77555 108455 77558
rect 109200 77528 110000 77558
rect 90766 77420 90772 77484
rect 90836 77482 90842 77484
rect 91553 77482 91619 77485
rect 90836 77480 91619 77482
rect 90836 77424 91558 77480
rect 91614 77424 91619 77480
rect 90836 77422 91619 77424
rect 90836 77420 90842 77422
rect 91553 77419 91619 77422
rect 4870 77280 5186 77281
rect 4870 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5186 77280
rect 4870 77215 5186 77216
rect 35590 77280 35906 77281
rect 35590 77216 35596 77280
rect 35660 77216 35676 77280
rect 35740 77216 35756 77280
rect 35820 77216 35836 77280
rect 35900 77216 35906 77280
rect 35590 77215 35906 77216
rect 66310 77280 66626 77281
rect 66310 77216 66316 77280
rect 66380 77216 66396 77280
rect 66460 77216 66476 77280
rect 66540 77216 66556 77280
rect 66620 77216 66626 77280
rect 66310 77215 66626 77216
rect 97030 77280 97346 77281
rect 97030 77216 97036 77280
rect 97100 77216 97116 77280
rect 97180 77216 97196 77280
rect 97260 77216 97276 77280
rect 97340 77216 97346 77280
rect 97030 77215 97346 77216
rect 106654 77280 106970 77281
rect 106654 77216 106660 77280
rect 106724 77216 106740 77280
rect 106804 77216 106820 77280
rect 106884 77216 106900 77280
rect 106964 77216 106970 77280
rect 106654 77215 106970 77216
rect 67909 77074 67975 77077
rect 103605 77074 103671 77077
rect 67909 77072 103671 77074
rect 67909 77016 67914 77072
rect 67970 77016 103610 77072
rect 103666 77016 103671 77072
rect 67909 77014 103671 77016
rect 67909 77011 67975 77014
rect 103605 77011 103671 77014
rect 0 76938 800 76968
rect 1209 76938 1275 76941
rect 0 76936 1275 76938
rect 0 76880 1214 76936
rect 1270 76880 1275 76936
rect 0 76878 1275 76880
rect 0 76848 800 76878
rect 1209 76875 1275 76878
rect 65977 76938 66043 76941
rect 103789 76938 103855 76941
rect 65977 76936 103855 76938
rect 65977 76880 65982 76936
rect 66038 76880 103794 76936
rect 103850 76880 103855 76936
rect 65977 76878 103855 76880
rect 65977 76875 66043 76878
rect 103789 76875 103855 76878
rect 108389 76938 108455 76941
rect 109200 76938 110000 76968
rect 108389 76936 110000 76938
rect 108389 76880 108394 76936
rect 108450 76880 110000 76936
rect 108389 76878 110000 76880
rect 108389 76875 108455 76878
rect 109200 76848 110000 76878
rect 4210 76736 4526 76737
rect 4210 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4526 76736
rect 4210 76671 4526 76672
rect 34930 76736 35246 76737
rect 34930 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35246 76736
rect 34930 76671 35246 76672
rect 65650 76736 65966 76737
rect 65650 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65966 76736
rect 65650 76671 65966 76672
rect 96370 76736 96686 76737
rect 96370 76672 96376 76736
rect 96440 76672 96456 76736
rect 96520 76672 96536 76736
rect 96600 76672 96616 76736
rect 96680 76672 96686 76736
rect 96370 76671 96686 76672
rect 63125 76530 63191 76533
rect 102225 76530 102291 76533
rect 63125 76528 102291 76530
rect 63125 76472 63130 76528
rect 63186 76472 102230 76528
rect 102286 76472 102291 76528
rect 63125 76470 102291 76472
rect 63125 76467 63191 76470
rect 102225 76467 102291 76470
rect 841 76394 907 76397
rect 798 76392 907 76394
rect 798 76336 846 76392
rect 902 76336 907 76392
rect 798 76331 907 76336
rect 61009 76394 61075 76397
rect 103697 76394 103763 76397
rect 61009 76392 103763 76394
rect 61009 76336 61014 76392
rect 61070 76336 103702 76392
rect 103758 76336 103763 76392
rect 61009 76334 103763 76336
rect 61009 76331 61075 76334
rect 103697 76331 103763 76334
rect 798 76288 858 76331
rect 0 76198 858 76288
rect 108389 76258 108455 76261
rect 109200 76258 110000 76288
rect 108389 76256 110000 76258
rect 108389 76200 108394 76256
rect 108450 76200 110000 76256
rect 108389 76198 110000 76200
rect 0 76168 800 76198
rect 108389 76195 108455 76198
rect 4870 76192 5186 76193
rect 4870 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5186 76192
rect 4870 76127 5186 76128
rect 35590 76192 35906 76193
rect 35590 76128 35596 76192
rect 35660 76128 35676 76192
rect 35740 76128 35756 76192
rect 35820 76128 35836 76192
rect 35900 76128 35906 76192
rect 35590 76127 35906 76128
rect 66310 76192 66626 76193
rect 66310 76128 66316 76192
rect 66380 76128 66396 76192
rect 66460 76128 66476 76192
rect 66540 76128 66556 76192
rect 66620 76128 66626 76192
rect 66310 76127 66626 76128
rect 97030 76192 97346 76193
rect 97030 76128 97036 76192
rect 97100 76128 97116 76192
rect 97180 76128 97196 76192
rect 97260 76128 97276 76192
rect 97340 76128 97346 76192
rect 109200 76168 110000 76198
rect 97030 76127 97346 76128
rect 84837 75986 84903 75989
rect 103513 75986 103579 75989
rect 84837 75984 103579 75986
rect 84837 75928 84842 75984
rect 84898 75928 103518 75984
rect 103574 75928 103579 75984
rect 84837 75926 103579 75928
rect 84837 75923 84903 75926
rect 103513 75923 103579 75926
rect 4210 75648 4526 75649
rect 0 75578 800 75608
rect 4210 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4526 75648
rect 4210 75583 4526 75584
rect 34930 75648 35246 75649
rect 34930 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35246 75648
rect 34930 75583 35246 75584
rect 65650 75648 65966 75649
rect 65650 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65966 75648
rect 65650 75583 65966 75584
rect 96370 75648 96686 75649
rect 96370 75584 96376 75648
rect 96440 75584 96456 75648
rect 96520 75584 96536 75648
rect 96600 75584 96616 75648
rect 96680 75584 96686 75648
rect 96370 75583 96686 75584
rect 1485 75578 1551 75581
rect 0 75576 1551 75578
rect 0 75520 1490 75576
rect 1546 75520 1551 75576
rect 0 75518 1551 75520
rect 0 75488 800 75518
rect 1485 75515 1551 75518
rect 108389 75578 108455 75581
rect 109200 75578 110000 75608
rect 108389 75576 110000 75578
rect 108389 75520 108394 75576
rect 108450 75520 110000 75576
rect 108389 75518 110000 75520
rect 108389 75515 108455 75518
rect 109200 75488 110000 75518
rect 4870 75104 5186 75105
rect 4870 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5186 75104
rect 4870 75039 5186 75040
rect 35590 75104 35906 75105
rect 35590 75040 35596 75104
rect 35660 75040 35676 75104
rect 35740 75040 35756 75104
rect 35820 75040 35836 75104
rect 35900 75040 35906 75104
rect 35590 75039 35906 75040
rect 66310 75104 66626 75105
rect 66310 75040 66316 75104
rect 66380 75040 66396 75104
rect 66460 75040 66476 75104
rect 66540 75040 66556 75104
rect 66620 75040 66626 75104
rect 66310 75039 66626 75040
rect 97030 75104 97346 75105
rect 97030 75040 97036 75104
rect 97100 75040 97116 75104
rect 97180 75040 97196 75104
rect 97260 75040 97276 75104
rect 97340 75040 97346 75104
rect 97030 75039 97346 75040
rect 841 75034 907 75037
rect 798 75032 907 75034
rect 798 74976 846 75032
rect 902 74976 907 75032
rect 798 74971 907 74976
rect 798 74928 858 74971
rect 0 74838 858 74928
rect 108389 74898 108455 74901
rect 109200 74898 110000 74928
rect 108389 74896 110000 74898
rect 108389 74840 108394 74896
rect 108450 74840 110000 74896
rect 108389 74838 110000 74840
rect 0 74808 800 74838
rect 108389 74835 108455 74838
rect 109200 74808 110000 74838
rect 4210 74560 4526 74561
rect 4210 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4526 74560
rect 4210 74495 4526 74496
rect 34930 74560 35246 74561
rect 34930 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35246 74560
rect 34930 74495 35246 74496
rect 65650 74560 65966 74561
rect 65650 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65966 74560
rect 65650 74495 65966 74496
rect 96370 74560 96686 74561
rect 96370 74496 96376 74560
rect 96440 74496 96456 74560
rect 96520 74496 96536 74560
rect 96600 74496 96616 74560
rect 96680 74496 96686 74560
rect 96370 74495 96686 74496
rect 99465 74490 99531 74493
rect 100385 74490 100451 74493
rect 99465 74488 100451 74490
rect 99465 74432 99470 74488
rect 99526 74432 100390 74488
rect 100446 74432 100451 74488
rect 99465 74430 100451 74432
rect 99465 74427 99531 74430
rect 100385 74427 100451 74430
rect 841 74354 907 74357
rect 798 74352 907 74354
rect 798 74296 846 74352
rect 902 74296 907 74352
rect 798 74291 907 74296
rect 798 74248 858 74291
rect 0 74158 858 74248
rect 98821 74218 98887 74221
rect 100201 74218 100267 74221
rect 100569 74218 100635 74221
rect 98821 74216 100635 74218
rect 98821 74160 98826 74216
rect 98882 74160 100206 74216
rect 100262 74160 100574 74216
rect 100630 74160 100635 74216
rect 98821 74158 100635 74160
rect 0 74128 800 74158
rect 98821 74155 98887 74158
rect 100201 74155 100267 74158
rect 100569 74155 100635 74158
rect 108389 74218 108455 74221
rect 109200 74218 110000 74248
rect 108389 74216 110000 74218
rect 108389 74160 108394 74216
rect 108450 74160 110000 74216
rect 108389 74158 110000 74160
rect 108389 74155 108455 74158
rect 109200 74128 110000 74158
rect 4870 74016 5186 74017
rect 4870 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5186 74016
rect 4870 73951 5186 73952
rect 35590 74016 35906 74017
rect 35590 73952 35596 74016
rect 35660 73952 35676 74016
rect 35740 73952 35756 74016
rect 35820 73952 35836 74016
rect 35900 73952 35906 74016
rect 35590 73951 35906 73952
rect 66310 74016 66626 74017
rect 66310 73952 66316 74016
rect 66380 73952 66396 74016
rect 66460 73952 66476 74016
rect 66540 73952 66556 74016
rect 66620 73952 66626 74016
rect 66310 73951 66626 73952
rect 97030 74016 97346 74017
rect 97030 73952 97036 74016
rect 97100 73952 97116 74016
rect 97180 73952 97196 74016
rect 97260 73952 97276 74016
rect 97340 73952 97346 74016
rect 97030 73951 97346 73952
rect 102501 73810 102567 73813
rect 104709 73810 104775 73813
rect 102501 73808 104775 73810
rect 102501 73752 102506 73808
rect 102562 73752 104714 73808
rect 104770 73752 104775 73808
rect 102501 73750 104775 73752
rect 102501 73747 102567 73750
rect 104709 73747 104775 73750
rect 841 73674 907 73677
rect 798 73672 907 73674
rect 798 73616 846 73672
rect 902 73616 907 73672
rect 798 73611 907 73616
rect 798 73568 858 73611
rect 0 73478 858 73568
rect 108481 73538 108547 73541
rect 109200 73538 110000 73568
rect 108481 73536 110000 73538
rect 108481 73480 108486 73536
rect 108542 73480 110000 73536
rect 108481 73478 110000 73480
rect 0 73448 800 73478
rect 108481 73475 108547 73478
rect 4210 73472 4526 73473
rect 4210 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4526 73472
rect 4210 73407 4526 73408
rect 34930 73472 35246 73473
rect 34930 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35246 73472
rect 34930 73407 35246 73408
rect 65650 73472 65966 73473
rect 65650 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65966 73472
rect 65650 73407 65966 73408
rect 96370 73472 96686 73473
rect 96370 73408 96376 73472
rect 96440 73408 96456 73472
rect 96520 73408 96536 73472
rect 96600 73408 96616 73472
rect 96680 73408 96686 73472
rect 109200 73448 110000 73478
rect 96370 73407 96686 73408
rect 98545 73402 98611 73405
rect 99465 73402 99531 73405
rect 98545 73400 99531 73402
rect 98545 73344 98550 73400
rect 98606 73344 99470 73400
rect 99526 73344 99531 73400
rect 98545 73342 99531 73344
rect 98545 73339 98611 73342
rect 99465 73339 99531 73342
rect 99097 73266 99163 73269
rect 99649 73266 99715 73269
rect 99097 73264 99715 73266
rect 99097 73208 99102 73264
rect 99158 73208 99654 73264
rect 99710 73208 99715 73264
rect 99097 73206 99715 73208
rect 99097 73203 99163 73206
rect 99649 73203 99715 73206
rect 841 72994 907 72997
rect 798 72992 907 72994
rect 798 72936 846 72992
rect 902 72936 907 72992
rect 798 72931 907 72936
rect 798 72888 858 72931
rect 0 72798 858 72888
rect 4870 72928 5186 72929
rect 4870 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5186 72928
rect 4870 72863 5186 72864
rect 35590 72928 35906 72929
rect 35590 72864 35596 72928
rect 35660 72864 35676 72928
rect 35740 72864 35756 72928
rect 35820 72864 35836 72928
rect 35900 72864 35906 72928
rect 35590 72863 35906 72864
rect 66310 72928 66626 72929
rect 66310 72864 66316 72928
rect 66380 72864 66396 72928
rect 66460 72864 66476 72928
rect 66540 72864 66556 72928
rect 66620 72864 66626 72928
rect 66310 72863 66626 72864
rect 97030 72928 97346 72929
rect 97030 72864 97036 72928
rect 97100 72864 97116 72928
rect 97180 72864 97196 72928
rect 97260 72864 97276 72928
rect 97340 72864 97346 72928
rect 97030 72863 97346 72864
rect 108481 72858 108547 72861
rect 109200 72858 110000 72888
rect 108481 72856 110000 72858
rect 108481 72800 108486 72856
rect 108542 72800 110000 72856
rect 108481 72798 110000 72800
rect 0 72768 800 72798
rect 108481 72795 108547 72798
rect 109200 72768 110000 72798
rect 86166 72524 86172 72588
rect 86236 72586 86242 72588
rect 88977 72586 89043 72589
rect 86236 72584 89043 72586
rect 86236 72528 88982 72584
rect 89038 72528 89043 72584
rect 86236 72526 89043 72528
rect 86236 72524 86242 72526
rect 88977 72523 89043 72526
rect 4210 72384 4526 72385
rect 4210 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4526 72384
rect 4210 72319 4526 72320
rect 34930 72384 35246 72385
rect 34930 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35246 72384
rect 34930 72319 35246 72320
rect 65650 72384 65966 72385
rect 65650 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65966 72384
rect 65650 72319 65966 72320
rect 96370 72384 96686 72385
rect 96370 72320 96376 72384
rect 96440 72320 96456 72384
rect 96520 72320 96536 72384
rect 96600 72320 96616 72384
rect 96680 72320 96686 72384
rect 96370 72319 96686 72320
rect 841 72314 907 72317
rect 798 72312 907 72314
rect 798 72256 846 72312
rect 902 72256 907 72312
rect 798 72251 907 72256
rect 798 72208 858 72251
rect 0 72118 858 72208
rect 108481 72178 108547 72181
rect 109200 72178 110000 72208
rect 108481 72176 110000 72178
rect 108481 72120 108486 72176
rect 108542 72120 110000 72176
rect 108481 72118 110000 72120
rect 0 72088 800 72118
rect 108481 72115 108547 72118
rect 109200 72088 110000 72118
rect 4870 71840 5186 71841
rect 4870 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5186 71840
rect 4870 71775 5186 71776
rect 35590 71840 35906 71841
rect 35590 71776 35596 71840
rect 35660 71776 35676 71840
rect 35740 71776 35756 71840
rect 35820 71776 35836 71840
rect 35900 71776 35906 71840
rect 35590 71775 35906 71776
rect 66310 71840 66626 71841
rect 66310 71776 66316 71840
rect 66380 71776 66396 71840
rect 66460 71776 66476 71840
rect 66540 71776 66556 71840
rect 66620 71776 66626 71840
rect 66310 71775 66626 71776
rect 97030 71840 97346 71841
rect 97030 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97346 71840
rect 97030 71775 97346 71776
rect 0 71498 800 71528
rect 1209 71498 1275 71501
rect 0 71496 1275 71498
rect 0 71440 1214 71496
rect 1270 71440 1275 71496
rect 0 71438 1275 71440
rect 0 71408 800 71438
rect 1209 71435 1275 71438
rect 108481 71498 108547 71501
rect 109200 71498 110000 71528
rect 108481 71496 110000 71498
rect 108481 71440 108486 71496
rect 108542 71440 110000 71496
rect 108481 71438 110000 71440
rect 108481 71435 108547 71438
rect 109200 71408 110000 71438
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 34930 71296 35246 71297
rect 34930 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35246 71296
rect 34930 71231 35246 71232
rect 65650 71296 65966 71297
rect 65650 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65966 71296
rect 65650 71231 65966 71232
rect 96370 71296 96686 71297
rect 96370 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96686 71296
rect 96370 71231 96686 71232
rect 97717 71090 97783 71093
rect 98177 71090 98243 71093
rect 97717 71088 98243 71090
rect 97717 71032 97722 71088
rect 97778 71032 98182 71088
rect 98238 71032 98243 71088
rect 97717 71030 98243 71032
rect 97717 71027 97783 71030
rect 98177 71027 98243 71030
rect 98821 70954 98887 70957
rect 101029 70954 101095 70957
rect 103513 70954 103579 70957
rect 98821 70952 103579 70954
rect 98821 70896 98826 70952
rect 98882 70896 101034 70952
rect 101090 70896 103518 70952
rect 103574 70896 103579 70952
rect 98821 70894 103579 70896
rect 98821 70891 98887 70894
rect 101029 70891 101095 70894
rect 103513 70891 103579 70894
rect 108481 70818 108547 70821
rect 109200 70818 110000 70848
rect 108481 70816 110000 70818
rect 108481 70760 108486 70816
rect 108542 70760 110000 70816
rect 108481 70758 110000 70760
rect 108481 70755 108547 70758
rect 4870 70752 5186 70753
rect 4870 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5186 70752
rect 4870 70687 5186 70688
rect 35590 70752 35906 70753
rect 35590 70688 35596 70752
rect 35660 70688 35676 70752
rect 35740 70688 35756 70752
rect 35820 70688 35836 70752
rect 35900 70688 35906 70752
rect 35590 70687 35906 70688
rect 66310 70752 66626 70753
rect 66310 70688 66316 70752
rect 66380 70688 66396 70752
rect 66460 70688 66476 70752
rect 66540 70688 66556 70752
rect 66620 70688 66626 70752
rect 66310 70687 66626 70688
rect 97030 70752 97346 70753
rect 97030 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97346 70752
rect 109200 70728 110000 70758
rect 97030 70687 97346 70688
rect 4210 70208 4526 70209
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 34930 70208 35246 70209
rect 34930 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35246 70208
rect 34930 70143 35246 70144
rect 65650 70208 65966 70209
rect 65650 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65966 70208
rect 65650 70143 65966 70144
rect 96370 70208 96686 70209
rect 96370 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96686 70208
rect 96370 70143 96686 70144
rect 108481 70138 108547 70141
rect 109200 70138 110000 70168
rect 108481 70136 110000 70138
rect 108481 70080 108486 70136
rect 108542 70080 110000 70136
rect 108481 70078 110000 70080
rect 108481 70075 108547 70078
rect 109200 70048 110000 70078
rect 97533 70002 97599 70005
rect 100017 70002 100083 70005
rect 97533 70000 100083 70002
rect 97533 69944 97538 70000
rect 97594 69944 100022 70000
rect 100078 69944 100083 70000
rect 97533 69942 100083 69944
rect 97533 69939 97599 69942
rect 100017 69939 100083 69942
rect 63534 69804 63540 69868
rect 63604 69866 63610 69868
rect 72693 69866 72759 69869
rect 63604 69864 72759 69866
rect 63604 69808 72698 69864
rect 72754 69808 72759 69864
rect 63604 69806 72759 69808
rect 63604 69804 63610 69806
rect 72693 69803 72759 69806
rect 73654 69804 73660 69868
rect 73724 69866 73730 69868
rect 79317 69866 79383 69869
rect 73724 69864 79383 69866
rect 73724 69808 79322 69864
rect 79378 69808 79383 69864
rect 73724 69806 79383 69808
rect 73724 69804 73730 69806
rect 79317 69803 79383 69806
rect 4870 69664 5186 69665
rect 4870 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5186 69664
rect 4870 69599 5186 69600
rect 35590 69664 35906 69665
rect 35590 69600 35596 69664
rect 35660 69600 35676 69664
rect 35740 69600 35756 69664
rect 35820 69600 35836 69664
rect 35900 69600 35906 69664
rect 35590 69599 35906 69600
rect 66310 69664 66626 69665
rect 66310 69600 66316 69664
rect 66380 69600 66396 69664
rect 66460 69600 66476 69664
rect 66540 69600 66556 69664
rect 66620 69600 66626 69664
rect 66310 69599 66626 69600
rect 97030 69664 97346 69665
rect 97030 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97346 69664
rect 97030 69599 97346 69600
rect 108481 69458 108547 69461
rect 109200 69458 110000 69488
rect 108481 69456 110000 69458
rect 108481 69400 108486 69456
rect 108542 69400 110000 69456
rect 108481 69398 110000 69400
rect 108481 69395 108547 69398
rect 109200 69368 110000 69398
rect 61142 69260 61148 69324
rect 61212 69322 61218 69324
rect 66437 69322 66503 69325
rect 61212 69320 66503 69322
rect 61212 69264 66442 69320
rect 66498 69264 66503 69320
rect 61212 69262 66503 69264
rect 61212 69260 61218 69262
rect 66437 69259 66503 69262
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 34930 69120 35246 69121
rect 34930 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35246 69120
rect 34930 69055 35246 69056
rect 65650 69120 65966 69121
rect 65650 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65966 69120
rect 65650 69055 65966 69056
rect 96370 69120 96686 69121
rect 96370 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96686 69120
rect 96370 69055 96686 69056
rect 100293 68914 100359 68917
rect 102726 68914 102732 68916
rect 100293 68912 102732 68914
rect 100293 68856 100298 68912
rect 100354 68856 102732 68912
rect 100293 68854 102732 68856
rect 100293 68851 100359 68854
rect 102726 68852 102732 68854
rect 102796 68852 102802 68916
rect 53598 68716 53604 68780
rect 53668 68778 53674 68780
rect 58709 68778 58775 68781
rect 53668 68776 58775 68778
rect 53668 68720 58714 68776
rect 58770 68720 58775 68776
rect 53668 68718 58775 68720
rect 53668 68716 53674 68718
rect 58709 68715 58775 68718
rect 56174 68580 56180 68644
rect 56244 68642 56250 68644
rect 61469 68642 61535 68645
rect 56244 68640 61535 68642
rect 56244 68584 61474 68640
rect 61530 68584 61535 68640
rect 56244 68582 61535 68584
rect 56244 68580 56250 68582
rect 61469 68579 61535 68582
rect 4870 68576 5186 68577
rect 4870 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5186 68576
rect 4870 68511 5186 68512
rect 35590 68576 35906 68577
rect 35590 68512 35596 68576
rect 35660 68512 35676 68576
rect 35740 68512 35756 68576
rect 35820 68512 35836 68576
rect 35900 68512 35906 68576
rect 35590 68511 35906 68512
rect 66310 68576 66626 68577
rect 66310 68512 66316 68576
rect 66380 68512 66396 68576
rect 66460 68512 66476 68576
rect 66540 68512 66556 68576
rect 66620 68512 66626 68576
rect 66310 68511 66626 68512
rect 97030 68576 97346 68577
rect 97030 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97346 68576
rect 97030 68511 97346 68512
rect 100845 68370 100911 68373
rect 104893 68370 104959 68373
rect 100845 68368 104959 68370
rect 100845 68312 100850 68368
rect 100906 68312 104898 68368
rect 104954 68312 104959 68368
rect 100845 68310 104959 68312
rect 100845 68307 100911 68310
rect 104893 68307 104959 68310
rect 43713 68234 43779 68237
rect 48630 68234 48636 68236
rect 43713 68232 48636 68234
rect 43713 68176 43718 68232
rect 43774 68176 48636 68232
rect 43713 68174 48636 68176
rect 43713 68171 43779 68174
rect 48630 68172 48636 68174
rect 48700 68172 48706 68236
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 34930 68032 35246 68033
rect 34930 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35246 68032
rect 34930 67967 35246 67968
rect 65650 68032 65966 68033
rect 65650 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65966 68032
rect 65650 67967 65966 67968
rect 96370 68032 96686 68033
rect 96370 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96686 68032
rect 96370 67967 96686 67968
rect 102133 67826 102199 67829
rect 102961 67826 103027 67829
rect 102133 67824 103027 67826
rect 102133 67768 102138 67824
rect 102194 67768 102966 67824
rect 103022 67768 103027 67824
rect 102133 67766 103027 67768
rect 102133 67763 102199 67766
rect 102961 67763 103027 67766
rect 97533 67690 97599 67693
rect 100845 67690 100911 67693
rect 97533 67688 100911 67690
rect 97533 67632 97538 67688
rect 97594 67632 100850 67688
rect 100906 67632 100911 67688
rect 97533 67630 100911 67632
rect 97533 67627 97599 67630
rect 100845 67627 100911 67630
rect 4870 67488 5186 67489
rect 4870 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5186 67488
rect 4870 67423 5186 67424
rect 35590 67488 35906 67489
rect 35590 67424 35596 67488
rect 35660 67424 35676 67488
rect 35740 67424 35756 67488
rect 35820 67424 35836 67488
rect 35900 67424 35906 67488
rect 35590 67423 35906 67424
rect 66310 67488 66626 67489
rect 66310 67424 66316 67488
rect 66380 67424 66396 67488
rect 66460 67424 66476 67488
rect 66540 67424 66556 67488
rect 66620 67424 66626 67488
rect 66310 67423 66626 67424
rect 97030 67488 97346 67489
rect 97030 67424 97036 67488
rect 97100 67424 97116 67488
rect 97180 67424 97196 67488
rect 97260 67424 97276 67488
rect 97340 67424 97346 67488
rect 97030 67423 97346 67424
rect 108481 67418 108547 67421
rect 109200 67418 110000 67448
rect 108481 67416 110000 67418
rect 108481 67360 108486 67416
rect 108542 67360 110000 67416
rect 108481 67358 110000 67360
rect 108481 67355 108547 67358
rect 109200 67328 110000 67358
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 96370 66944 96686 66945
rect 96370 66880 96376 66944
rect 96440 66880 96456 66944
rect 96520 66880 96536 66944
rect 96600 66880 96616 66944
rect 96680 66880 96686 66944
rect 96370 66879 96686 66880
rect 4870 66400 5186 66401
rect 4870 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5186 66400
rect 4870 66335 5186 66336
rect 35590 66400 35906 66401
rect 35590 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35906 66400
rect 35590 66335 35906 66336
rect 66310 66400 66626 66401
rect 66310 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66626 66400
rect 66310 66335 66626 66336
rect 97030 66400 97346 66401
rect 97030 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97346 66400
rect 97030 66335 97346 66336
rect 106654 66400 106970 66401
rect 106654 66336 106660 66400
rect 106724 66336 106740 66400
rect 106804 66336 106820 66400
rect 106884 66336 106900 66400
rect 106964 66336 106970 66400
rect 106654 66335 106970 66336
rect 68502 66132 68508 66196
rect 68572 66194 68578 66196
rect 68645 66194 68711 66197
rect 68572 66192 68711 66194
rect 68572 66136 68650 66192
rect 68706 66136 68711 66192
rect 68572 66134 68711 66136
rect 68572 66132 68578 66134
rect 68645 66131 68711 66134
rect 87270 65860 87276 65924
rect 87340 65922 87346 65924
rect 88241 65922 88307 65925
rect 87340 65920 88307 65922
rect 87340 65864 88246 65920
rect 88302 65864 88307 65920
rect 87340 65862 88307 65864
rect 87340 65860 87346 65862
rect 88241 65859 88307 65862
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 96370 65856 96686 65857
rect 96370 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96686 65856
rect 96370 65791 96686 65792
rect 105918 65856 106234 65857
rect 105918 65792 105924 65856
rect 105988 65792 106004 65856
rect 106068 65792 106084 65856
rect 106148 65792 106164 65856
rect 106228 65792 106234 65856
rect 105918 65791 106234 65792
rect 34513 65650 34579 65653
rect 36118 65650 36124 65652
rect 34513 65648 36124 65650
rect 34513 65592 34518 65648
rect 34574 65592 36124 65648
rect 34513 65590 36124 65592
rect 34513 65587 34579 65590
rect 36118 65588 36124 65590
rect 36188 65588 36194 65652
rect 45093 65650 45159 65653
rect 46054 65650 46060 65652
rect 45093 65648 46060 65650
rect 45093 65592 45098 65648
rect 45154 65592 46060 65648
rect 45093 65590 46060 65592
rect 45093 65587 45159 65590
rect 46054 65588 46060 65590
rect 46124 65588 46130 65652
rect 31661 65514 31727 65517
rect 38510 65514 38516 65516
rect 31661 65512 38516 65514
rect 31661 65456 31666 65512
rect 31722 65456 38516 65512
rect 31661 65454 38516 65456
rect 31661 65451 31727 65454
rect 38510 65452 38516 65454
rect 38580 65452 38586 65516
rect 4870 65312 5186 65313
rect 4870 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5186 65312
rect 4870 65247 5186 65248
rect 106654 65312 106970 65313
rect 106654 65248 106660 65312
rect 106724 65248 106740 65312
rect 106804 65248 106820 65312
rect 106884 65248 106900 65312
rect 106964 65248 106970 65312
rect 106654 65247 106970 65248
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 105918 64768 106234 64769
rect 105918 64704 105924 64768
rect 105988 64704 106004 64768
rect 106068 64704 106084 64768
rect 106148 64704 106164 64768
rect 106228 64704 106234 64768
rect 105918 64703 106234 64704
rect 41137 64292 41203 64293
rect 41086 64290 41092 64292
rect 41046 64230 41092 64290
rect 41156 64288 41203 64292
rect 41198 64232 41203 64288
rect 41086 64228 41092 64230
rect 41156 64228 41203 64232
rect 41137 64227 41203 64228
rect 4870 64224 5186 64225
rect 4870 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5186 64224
rect 4870 64159 5186 64160
rect 106654 64224 106970 64225
rect 106654 64160 106660 64224
rect 106724 64160 106740 64224
rect 106804 64160 106820 64224
rect 106884 64160 106900 64224
rect 106964 64160 106970 64224
rect 106654 64159 106970 64160
rect 39941 64154 40007 64157
rect 43557 64154 43563 64156
rect 39941 64152 43563 64154
rect 39941 64096 39946 64152
rect 40002 64096 43563 64152
rect 39941 64094 43563 64096
rect 39941 64091 40007 64094
rect 43557 64092 43563 64094
rect 43627 64092 43633 64156
rect 46473 64154 46539 64157
rect 51045 64154 51051 64156
rect 46473 64152 51051 64154
rect 46473 64096 46478 64152
rect 46534 64096 51051 64152
rect 46473 64094 51051 64096
rect 46473 64091 46539 64094
rect 51045 64092 51051 64094
rect 51115 64092 51121 64156
rect 58533 64092 58539 64156
rect 58603 64154 58609 64156
rect 66069 64154 66135 64157
rect 95877 64156 95943 64157
rect 95852 64154 95858 64156
rect 58603 64152 66135 64154
rect 58603 64096 66074 64152
rect 66130 64096 66135 64152
rect 58603 64094 66135 64096
rect 95786 64094 95858 64154
rect 95922 64152 95943 64156
rect 95938 64096 95943 64152
rect 58603 64092 58609 64094
rect 66069 64091 66135 64094
rect 95852 64092 95858 64094
rect 95922 64092 95943 64096
rect 95877 64091 95943 64092
rect 66021 63956 66027 64020
rect 66091 64018 66097 64020
rect 72417 64018 72483 64021
rect 66091 64016 72483 64018
rect 66091 63960 72422 64016
rect 72478 63960 72483 64016
rect 66091 63958 72483 63960
rect 66091 63956 66097 63958
rect 72417 63955 72483 63958
rect 71013 63820 71019 63884
rect 71083 63882 71089 63884
rect 77845 63882 77911 63885
rect 71083 63880 77911 63882
rect 71083 63824 77850 63880
rect 77906 63824 77911 63880
rect 71083 63822 77911 63824
rect 71083 63820 71089 63822
rect 77845 63819 77911 63822
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 105918 63680 106234 63681
rect 105918 63616 105924 63680
rect 105988 63616 106004 63680
rect 106068 63616 106084 63680
rect 106148 63616 106164 63680
rect 106228 63616 106234 63680
rect 105918 63615 106234 63616
rect 4870 63136 5186 63137
rect 4870 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5186 63136
rect 4870 63071 5186 63072
rect 106654 63136 106970 63137
rect 106654 63072 106660 63136
rect 106724 63072 106740 63136
rect 106804 63072 106820 63136
rect 106884 63072 106900 63136
rect 106964 63072 106970 63136
rect 106654 63071 106970 63072
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 105918 62592 106234 62593
rect 105918 62528 105924 62592
rect 105988 62528 106004 62592
rect 106068 62528 106084 62592
rect 106148 62528 106164 62592
rect 106228 62528 106234 62592
rect 105918 62527 106234 62528
rect 4870 62048 5186 62049
rect 4870 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5186 62048
rect 4870 61983 5186 61984
rect 106654 62048 106970 62049
rect 106654 61984 106660 62048
rect 106724 61984 106740 62048
rect 106804 61984 106820 62048
rect 106884 61984 106900 62048
rect 106964 61984 106970 62048
rect 106654 61983 106970 61984
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 105918 61504 106234 61505
rect 105918 61440 105924 61504
rect 105988 61440 106004 61504
rect 106068 61440 106084 61504
rect 106148 61440 106164 61504
rect 106228 61440 106234 61504
rect 105918 61439 106234 61440
rect 4870 60960 5186 60961
rect 4870 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5186 60960
rect 4870 60895 5186 60896
rect 106654 60960 106970 60961
rect 106654 60896 106660 60960
rect 106724 60896 106740 60960
rect 106804 60896 106820 60960
rect 106884 60896 106900 60960
rect 106964 60896 106970 60960
rect 106654 60895 106970 60896
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 105918 60416 106234 60417
rect 105918 60352 105924 60416
rect 105988 60352 106004 60416
rect 106068 60352 106084 60416
rect 106148 60352 106164 60416
rect 106228 60352 106234 60416
rect 105918 60351 106234 60352
rect 4870 59872 5186 59873
rect 4870 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5186 59872
rect 4870 59807 5186 59808
rect 106654 59872 106970 59873
rect 106654 59808 106660 59872
rect 106724 59808 106740 59872
rect 106804 59808 106820 59872
rect 106884 59808 106900 59872
rect 106964 59808 106970 59872
rect 106654 59807 106970 59808
rect 104341 59802 104407 59805
rect 102550 59800 104407 59802
rect 102550 59768 104346 59800
rect 101948 59744 104346 59768
rect 104402 59744 104407 59800
rect 101948 59742 104407 59744
rect 101948 59708 102610 59742
rect 104341 59739 104407 59742
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 105918 59328 106234 59329
rect 105918 59264 105924 59328
rect 105988 59264 106004 59328
rect 106068 59264 106084 59328
rect 106148 59264 106164 59328
rect 106228 59264 106234 59328
rect 105918 59263 106234 59264
rect 4870 58784 5186 58785
rect 4870 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5186 58784
rect 4870 58719 5186 58720
rect 106654 58784 106970 58785
rect 106654 58720 106660 58784
rect 106724 58720 106740 58784
rect 106804 58720 106820 58784
rect 106884 58720 106900 58784
rect 106964 58720 106970 58784
rect 106654 58719 106970 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 105918 58240 106234 58241
rect 105918 58176 105924 58240
rect 105988 58176 106004 58240
rect 106068 58176 106084 58240
rect 106148 58176 106164 58240
rect 106228 58176 106234 58240
rect 105918 58175 106234 58176
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 106654 57696 106970 57697
rect 106654 57632 106660 57696
rect 106724 57632 106740 57696
rect 106804 57632 106820 57696
rect 106884 57632 106900 57696
rect 106964 57632 106970 57696
rect 106654 57631 106970 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 105918 57152 106234 57153
rect 105918 57088 105924 57152
rect 105988 57088 106004 57152
rect 106068 57088 106084 57152
rect 106148 57088 106164 57152
rect 106228 57088 106234 57152
rect 105918 57087 106234 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 106654 56608 106970 56609
rect 106654 56544 106660 56608
rect 106724 56544 106740 56608
rect 106804 56544 106820 56608
rect 106884 56544 106900 56608
rect 106964 56544 106970 56608
rect 106654 56543 106970 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 105918 56064 106234 56065
rect 105918 56000 105924 56064
rect 105988 56000 106004 56064
rect 106068 56000 106084 56064
rect 106148 56000 106164 56064
rect 106228 56000 106234 56064
rect 105918 55999 106234 56000
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 106654 55520 106970 55521
rect 106654 55456 106660 55520
rect 106724 55456 106740 55520
rect 106804 55456 106820 55520
rect 106884 55456 106900 55520
rect 106964 55456 106970 55520
rect 106654 55455 106970 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 105918 54976 106234 54977
rect 105918 54912 105924 54976
rect 105988 54912 106004 54976
rect 106068 54912 106084 54976
rect 106148 54912 106164 54976
rect 106228 54912 106234 54976
rect 105918 54911 106234 54912
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 106654 54432 106970 54433
rect 106654 54368 106660 54432
rect 106724 54368 106740 54432
rect 106804 54368 106820 54432
rect 106884 54368 106900 54432
rect 106964 54368 106970 54432
rect 106654 54367 106970 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 105918 53888 106234 53889
rect 105918 53824 105924 53888
rect 105988 53824 106004 53888
rect 106068 53824 106084 53888
rect 106148 53824 106164 53888
rect 106228 53824 106234 53888
rect 105918 53823 106234 53824
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 106654 53344 106970 53345
rect 106654 53280 106660 53344
rect 106724 53280 106740 53344
rect 106804 53280 106820 53344
rect 106884 53280 106900 53344
rect 106964 53280 106970 53344
rect 106654 53279 106970 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 105918 52800 106234 52801
rect 105918 52736 105924 52800
rect 105988 52736 106004 52800
rect 106068 52736 106084 52800
rect 106148 52736 106164 52800
rect 106228 52736 106234 52800
rect 105918 52735 106234 52736
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 106654 52256 106970 52257
rect 106654 52192 106660 52256
rect 106724 52192 106740 52256
rect 106804 52192 106820 52256
rect 106884 52192 106900 52256
rect 106964 52192 106970 52256
rect 106654 52191 106970 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 105918 51712 106234 51713
rect 105918 51648 105924 51712
rect 105988 51648 106004 51712
rect 106068 51648 106084 51712
rect 106148 51648 106164 51712
rect 106228 51648 106234 51712
rect 105918 51647 106234 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 106654 51168 106970 51169
rect 106654 51104 106660 51168
rect 106724 51104 106740 51168
rect 106804 51104 106820 51168
rect 106884 51104 106900 51168
rect 106964 51104 106970 51168
rect 106654 51103 106970 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 105918 50624 106234 50625
rect 105918 50560 105924 50624
rect 105988 50560 106004 50624
rect 106068 50560 106084 50624
rect 106148 50560 106164 50624
rect 106228 50560 106234 50624
rect 105918 50559 106234 50560
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 106654 50080 106970 50081
rect 106654 50016 106660 50080
rect 106724 50016 106740 50080
rect 106804 50016 106820 50080
rect 106884 50016 106900 50080
rect 106964 50016 106970 50080
rect 106654 50015 106970 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 105918 49536 106234 49537
rect 105918 49472 105924 49536
rect 105988 49472 106004 49536
rect 106068 49472 106084 49536
rect 106148 49472 106164 49536
rect 106228 49472 106234 49536
rect 105918 49471 106234 49472
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 106654 48992 106970 48993
rect 106654 48928 106660 48992
rect 106724 48928 106740 48992
rect 106804 48928 106820 48992
rect 106884 48928 106900 48992
rect 106964 48928 106970 48992
rect 106654 48927 106970 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 105918 48448 106234 48449
rect 105918 48384 105924 48448
rect 105988 48384 106004 48448
rect 106068 48384 106084 48448
rect 106148 48384 106164 48448
rect 106228 48384 106234 48448
rect 105918 48383 106234 48384
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 106654 47904 106970 47905
rect 106654 47840 106660 47904
rect 106724 47840 106740 47904
rect 106804 47840 106820 47904
rect 106884 47840 106900 47904
rect 106964 47840 106970 47904
rect 106654 47839 106970 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 105918 47360 106234 47361
rect 105918 47296 105924 47360
rect 105988 47296 106004 47360
rect 106068 47296 106084 47360
rect 106148 47296 106164 47360
rect 106228 47296 106234 47360
rect 105918 47295 106234 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 106654 46816 106970 46817
rect 106654 46752 106660 46816
rect 106724 46752 106740 46816
rect 106804 46752 106820 46816
rect 106884 46752 106900 46816
rect 106964 46752 106970 46816
rect 106654 46751 106970 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 105918 46272 106234 46273
rect 105918 46208 105924 46272
rect 105988 46208 106004 46272
rect 106068 46208 106084 46272
rect 106148 46208 106164 46272
rect 106228 46208 106234 46272
rect 105918 46207 106234 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 106654 45728 106970 45729
rect 106654 45664 106660 45728
rect 106724 45664 106740 45728
rect 106804 45664 106820 45728
rect 106884 45664 106900 45728
rect 106964 45664 106970 45728
rect 106654 45663 106970 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 105918 45184 106234 45185
rect 105918 45120 105924 45184
rect 105988 45120 106004 45184
rect 106068 45120 106084 45184
rect 106148 45120 106164 45184
rect 106228 45120 106234 45184
rect 105918 45119 106234 45120
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 106654 44640 106970 44641
rect 106654 44576 106660 44640
rect 106724 44576 106740 44640
rect 106804 44576 106820 44640
rect 106884 44576 106900 44640
rect 106964 44576 106970 44640
rect 106654 44575 106970 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 105918 44096 106234 44097
rect 105918 44032 105924 44096
rect 105988 44032 106004 44096
rect 106068 44032 106084 44096
rect 106148 44032 106164 44096
rect 106228 44032 106234 44096
rect 105918 44031 106234 44032
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 106654 43552 106970 43553
rect 106654 43488 106660 43552
rect 106724 43488 106740 43552
rect 106804 43488 106820 43552
rect 106884 43488 106900 43552
rect 106964 43488 106970 43552
rect 106654 43487 106970 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 105918 43008 106234 43009
rect 105918 42944 105924 43008
rect 105988 42944 106004 43008
rect 106068 42944 106084 43008
rect 106148 42944 106164 43008
rect 106228 42944 106234 43008
rect 105918 42943 106234 42944
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 106654 42464 106970 42465
rect 106654 42400 106660 42464
rect 106724 42400 106740 42464
rect 106804 42400 106820 42464
rect 106884 42400 106900 42464
rect 106964 42400 106970 42464
rect 106654 42399 106970 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 105918 41920 106234 41921
rect 105918 41856 105924 41920
rect 105988 41856 106004 41920
rect 106068 41856 106084 41920
rect 106148 41856 106164 41920
rect 106228 41856 106234 41920
rect 105918 41855 106234 41856
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 106654 41376 106970 41377
rect 106654 41312 106660 41376
rect 106724 41312 106740 41376
rect 106804 41312 106820 41376
rect 106884 41312 106900 41376
rect 106964 41312 106970 41376
rect 106654 41311 106970 41312
rect 7557 41306 7623 41309
rect 7557 41304 9506 41306
rect 7557 41248 7562 41304
rect 7618 41254 9506 41304
rect 7618 41248 10028 41254
rect 7557 41246 10028 41248
rect 7557 41243 7623 41246
rect 9446 41194 10028 41246
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 105918 40832 106234 40833
rect 105918 40768 105924 40832
rect 105988 40768 106004 40832
rect 106068 40768 106084 40832
rect 106148 40768 106164 40832
rect 106228 40768 106234 40832
rect 105918 40767 106234 40768
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 106654 40288 106970 40289
rect 106654 40224 106660 40288
rect 106724 40224 106740 40288
rect 106804 40224 106820 40288
rect 106884 40224 106900 40288
rect 106964 40224 106970 40288
rect 106654 40223 106970 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 105918 39744 106234 39745
rect 105918 39680 105924 39744
rect 105988 39680 106004 39744
rect 106068 39680 106084 39744
rect 106148 39680 106164 39744
rect 106228 39680 106234 39744
rect 105918 39679 106234 39680
rect 7281 39538 7347 39541
rect 9446 39538 10028 39554
rect 7281 39536 10028 39538
rect 7281 39480 7286 39536
rect 7342 39494 10028 39536
rect 7342 39480 9506 39494
rect 7281 39478 9506 39480
rect 7281 39475 7347 39478
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 106654 39200 106970 39201
rect 106654 39136 106660 39200
rect 106724 39136 106740 39200
rect 106804 39136 106820 39200
rect 106884 39136 106900 39200
rect 106964 39136 106970 39200
rect 106654 39135 106970 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 105918 38656 106234 38657
rect 105918 38592 105924 38656
rect 105988 38592 106004 38656
rect 106068 38592 106084 38656
rect 106148 38592 106164 38656
rect 106228 38592 106234 38656
rect 105918 38591 106234 38592
rect 7557 38450 7623 38453
rect 7557 38448 9506 38450
rect 7557 38392 7562 38448
rect 7618 38426 9506 38448
rect 7618 38392 10028 38426
rect 7557 38390 10028 38392
rect 7557 38387 7623 38390
rect 9446 38366 10028 38390
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 106654 38112 106970 38113
rect 106654 38048 106660 38112
rect 106724 38048 106740 38112
rect 106804 38048 106820 38112
rect 106884 38048 106900 38112
rect 106964 38048 106970 38112
rect 106654 38047 106970 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 105918 37568 106234 37569
rect 105918 37504 105924 37568
rect 105988 37504 106004 37568
rect 106068 37504 106084 37568
rect 106148 37504 106164 37568
rect 106228 37504 106234 37568
rect 105918 37503 106234 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 106654 37024 106970 37025
rect 106654 36960 106660 37024
rect 106724 36960 106740 37024
rect 106804 36960 106820 37024
rect 106884 36960 106900 37024
rect 106964 36960 106970 37024
rect 106654 36959 106970 36960
rect 7557 36682 7623 36685
rect 9446 36682 10028 36726
rect 7557 36680 10028 36682
rect 7557 36624 7562 36680
rect 7618 36666 10028 36680
rect 7618 36624 9506 36666
rect 7557 36622 9506 36624
rect 7557 36619 7623 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 105918 36480 106234 36481
rect 105918 36416 105924 36480
rect 105988 36416 106004 36480
rect 106068 36416 106084 36480
rect 106148 36416 106164 36480
rect 106228 36416 106234 36480
rect 105918 36415 106234 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 106654 35936 106970 35937
rect 106654 35872 106660 35936
rect 106724 35872 106740 35936
rect 106804 35872 106820 35936
rect 106884 35872 106900 35936
rect 106964 35872 106970 35936
rect 106654 35871 106970 35872
rect 7465 35594 7531 35597
rect 9446 35594 10028 35643
rect 7465 35592 10028 35594
rect 7465 35536 7470 35592
rect 7526 35583 10028 35592
rect 7526 35536 9506 35583
rect 7465 35534 9506 35536
rect 7465 35531 7531 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 105918 35392 106234 35393
rect 105918 35328 105924 35392
rect 105988 35328 106004 35392
rect 106068 35328 106084 35392
rect 106148 35328 106164 35392
rect 106228 35328 106234 35392
rect 105918 35327 106234 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 106654 34848 106970 34849
rect 106654 34784 106660 34848
rect 106724 34784 106740 34848
rect 106804 34784 106820 34848
rect 106884 34784 106900 34848
rect 106964 34784 106970 34848
rect 106654 34783 106970 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 105918 34304 106234 34305
rect 105918 34240 105924 34304
rect 105988 34240 106004 34304
rect 106068 34240 106084 34304
rect 106148 34240 106164 34304
rect 106228 34240 106234 34304
rect 105918 34239 106234 34240
rect 7557 33962 7623 33965
rect 9446 33962 10028 33963
rect 7557 33960 10028 33962
rect 7557 33904 7562 33960
rect 7618 33904 10028 33960
rect 7557 33903 10028 33904
rect 7557 33902 9506 33903
rect 7557 33899 7623 33902
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 106654 33760 106970 33761
rect 106654 33696 106660 33760
rect 106724 33696 106740 33760
rect 106804 33696 106820 33760
rect 106884 33696 106900 33760
rect 106964 33696 106970 33760
rect 106654 33695 106970 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 105918 33216 106234 33217
rect 105918 33152 105924 33216
rect 105988 33152 106004 33216
rect 106068 33152 106084 33216
rect 106148 33152 106164 33216
rect 106228 33152 106234 33216
rect 105918 33151 106234 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 106654 32672 106970 32673
rect 106654 32608 106660 32672
rect 106724 32608 106740 32672
rect 106804 32608 106820 32672
rect 106884 32608 106900 32672
rect 106964 32608 106970 32672
rect 106654 32607 106970 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 105918 32128 106234 32129
rect 105918 32064 105924 32128
rect 105988 32064 106004 32128
rect 106068 32064 106084 32128
rect 106148 32064 106164 32128
rect 106228 32064 106234 32128
rect 105918 32063 106234 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 106654 31584 106970 31585
rect 106654 31520 106660 31584
rect 106724 31520 106740 31584
rect 106804 31520 106820 31584
rect 106884 31520 106900 31584
rect 106964 31520 106970 31584
rect 106654 31519 106970 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 105918 31040 106234 31041
rect 105918 30976 105924 31040
rect 105988 30976 106004 31040
rect 106068 30976 106084 31040
rect 106148 30976 106164 31040
rect 106228 30976 106234 31040
rect 105918 30975 106234 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 106654 30496 106970 30497
rect 106654 30432 106660 30496
rect 106724 30432 106740 30496
rect 106804 30432 106820 30496
rect 106884 30432 106900 30496
rect 106964 30432 106970 30496
rect 106654 30431 106970 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 105918 29952 106234 29953
rect 105918 29888 105924 29952
rect 105988 29888 106004 29952
rect 106068 29888 106084 29952
rect 106148 29888 106164 29952
rect 106228 29888 106234 29952
rect 105918 29887 106234 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 106654 29408 106970 29409
rect 106654 29344 106660 29408
rect 106724 29344 106740 29408
rect 106804 29344 106820 29408
rect 106884 29344 106900 29408
rect 106964 29344 106970 29408
rect 106654 29343 106970 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 105918 28864 106234 28865
rect 105918 28800 105924 28864
rect 105988 28800 106004 28864
rect 106068 28800 106084 28864
rect 106148 28800 106164 28864
rect 106228 28800 106234 28864
rect 105918 28799 106234 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 106654 28320 106970 28321
rect 106654 28256 106660 28320
rect 106724 28256 106740 28320
rect 106804 28256 106820 28320
rect 106884 28256 106900 28320
rect 106964 28256 106970 28320
rect 106654 28255 106970 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 105918 27776 106234 27777
rect 105918 27712 105924 27776
rect 105988 27712 106004 27776
rect 106068 27712 106084 27776
rect 106148 27712 106164 27776
rect 106228 27712 106234 27776
rect 105918 27711 106234 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 106654 27232 106970 27233
rect 106654 27168 106660 27232
rect 106724 27168 106740 27232
rect 106804 27168 106820 27232
rect 106884 27168 106900 27232
rect 106964 27168 106970 27232
rect 106654 27167 106970 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 105918 26688 106234 26689
rect 105918 26624 105924 26688
rect 105988 26624 106004 26688
rect 106068 26624 106084 26688
rect 106148 26624 106164 26688
rect 106228 26624 106234 26688
rect 105918 26623 106234 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 106654 26144 106970 26145
rect 106654 26080 106660 26144
rect 106724 26080 106740 26144
rect 106804 26080 106820 26144
rect 106884 26080 106900 26144
rect 106964 26080 106970 26144
rect 106654 26079 106970 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 105918 25600 106234 25601
rect 105918 25536 105924 25600
rect 105988 25536 106004 25600
rect 106068 25536 106084 25600
rect 106148 25536 106164 25600
rect 106228 25536 106234 25600
rect 105918 25535 106234 25536
rect 102593 25122 102659 25125
rect 102550 25120 102659 25122
rect 102225 25090 102291 25093
rect 102550 25090 102598 25120
rect 101948 25088 102598 25090
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 101948 25032 102230 25088
rect 102286 25064 102598 25088
rect 102654 25064 102659 25120
rect 102286 25059 102659 25064
rect 102286 25032 102610 25059
rect 101948 25030 102610 25032
rect 106654 25056 106970 25057
rect 102225 25027 102291 25030
rect 4870 24991 5186 24992
rect 106654 24992 106660 25056
rect 106724 24992 106740 25056
rect 106804 24992 106820 25056
rect 106884 24992 106900 25056
rect 106964 24992 106970 25056
rect 106654 24991 106970 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 105918 24512 106234 24513
rect 105918 24448 105924 24512
rect 105988 24448 106004 24512
rect 106068 24448 106084 24512
rect 106148 24448 106164 24512
rect 106228 24448 106234 24512
rect 105918 24447 106234 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 106654 23968 106970 23969
rect 106654 23904 106660 23968
rect 106724 23904 106740 23968
rect 106804 23904 106820 23968
rect 106884 23904 106900 23968
rect 106964 23904 106970 23968
rect 106654 23903 106970 23904
rect 102777 23492 102843 23493
rect 102726 23490 102732 23492
rect 102182 23430 102732 23490
rect 102796 23490 102843 23492
rect 102796 23488 102924 23490
rect 102838 23432 102924 23488
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 102182 23390 102242 23430
rect 102726 23428 102732 23430
rect 102796 23430 102924 23432
rect 102796 23428 102843 23430
rect 102777 23427 102843 23428
rect 4210 23359 4526 23360
rect 101948 23330 102242 23390
rect 105918 23424 106234 23425
rect 105918 23360 105924 23424
rect 105988 23360 106004 23424
rect 106068 23360 106084 23424
rect 106148 23360 106164 23424
rect 106228 23360 106234 23424
rect 105918 23359 106234 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 106654 22880 106970 22881
rect 106654 22816 106660 22880
rect 106724 22816 106740 22880
rect 106804 22816 106820 22880
rect 106884 22816 106900 22880
rect 106964 22816 106970 22880
rect 106654 22815 106970 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 105918 22336 106234 22337
rect 105918 22272 105924 22336
rect 105988 22272 106004 22336
rect 106068 22272 106084 22336
rect 106148 22272 106164 22336
rect 106228 22272 106234 22336
rect 105918 22271 106234 22272
rect 102133 22262 102199 22265
rect 101948 22260 102199 22262
rect 101948 22204 102138 22260
rect 102194 22204 102199 22260
rect 101948 22202 102199 22204
rect 102133 22199 102199 22202
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 106654 21792 106970 21793
rect 106654 21728 106660 21792
rect 106724 21728 106740 21792
rect 106804 21728 106820 21792
rect 106884 21728 106900 21792
rect 106964 21728 106970 21792
rect 106654 21727 106970 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 105918 21248 106234 21249
rect 105918 21184 105924 21248
rect 105988 21184 106004 21248
rect 106068 21184 106084 21248
rect 106148 21184 106164 21248
rect 106228 21184 106234 21248
rect 105918 21183 106234 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 106654 20704 106970 20705
rect 106654 20640 106660 20704
rect 106724 20640 106740 20704
rect 106804 20640 106820 20704
rect 106884 20640 106900 20704
rect 106964 20640 106970 20704
rect 106654 20639 106970 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 105918 20160 106234 20161
rect 105918 20096 105924 20160
rect 105988 20096 106004 20160
rect 106068 20096 106084 20160
rect 106148 20096 106164 20160
rect 106228 20096 106234 20160
rect 105918 20095 106234 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 106654 19616 106970 19617
rect 106654 19552 106660 19616
rect 106724 19552 106740 19616
rect 106804 19552 106820 19616
rect 106884 19552 106900 19616
rect 106964 19552 106970 19616
rect 106654 19551 106970 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 105918 19072 106234 19073
rect 105918 19008 105924 19072
rect 105988 19008 106004 19072
rect 106068 19008 106084 19072
rect 106148 19008 106164 19072
rect 106228 19008 106234 19072
rect 105918 19007 106234 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 106654 18528 106970 18529
rect 106654 18464 106660 18528
rect 106724 18464 106740 18528
rect 106804 18464 106820 18528
rect 106884 18464 106900 18528
rect 106964 18464 106970 18528
rect 106654 18463 106970 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 105918 17984 106234 17985
rect 105918 17920 105924 17984
rect 105988 17920 106004 17984
rect 106068 17920 106084 17984
rect 106148 17920 106164 17984
rect 106228 17920 106234 17984
rect 105918 17919 106234 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 106654 17440 106970 17441
rect 106654 17376 106660 17440
rect 106724 17376 106740 17440
rect 106804 17376 106820 17440
rect 106884 17376 106900 17440
rect 106964 17376 106970 17440
rect 106654 17375 106970 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 105918 16896 106234 16897
rect 105918 16832 105924 16896
rect 105988 16832 106004 16896
rect 106068 16832 106084 16896
rect 106148 16832 106164 16896
rect 106228 16832 106234 16896
rect 105918 16831 106234 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 106654 16352 106970 16353
rect 106654 16288 106660 16352
rect 106724 16288 106740 16352
rect 106804 16288 106820 16352
rect 106884 16288 106900 16352
rect 106964 16288 106970 16352
rect 106654 16287 106970 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 105918 15808 106234 15809
rect 105918 15744 105924 15808
rect 105988 15744 106004 15808
rect 106068 15744 106084 15808
rect 106148 15744 106164 15808
rect 106228 15744 106234 15808
rect 105918 15743 106234 15744
rect 7465 15466 7531 15469
rect 9446 15466 10028 15483
rect 7465 15464 10028 15466
rect 7465 15408 7470 15464
rect 7526 15423 10028 15464
rect 7526 15408 9506 15423
rect 7465 15406 9506 15408
rect 7465 15403 7531 15406
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 106654 15264 106970 15265
rect 106654 15200 106660 15264
rect 106724 15200 106740 15264
rect 106804 15200 106820 15264
rect 106884 15200 106900 15264
rect 106964 15200 106970 15264
rect 106654 15199 106970 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 105918 14720 106234 14721
rect 105918 14656 105924 14720
rect 105988 14656 106004 14720
rect 106068 14656 106084 14720
rect 106148 14656 106164 14720
rect 106228 14656 106234 14720
rect 105918 14655 106234 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 106654 14176 106970 14177
rect 106654 14112 106660 14176
rect 106724 14112 106740 14176
rect 106804 14112 106820 14176
rect 106884 14112 106900 14176
rect 106964 14112 106970 14176
rect 106654 14111 106970 14112
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 105918 13632 106234 13633
rect 105918 13568 105924 13632
rect 105988 13568 106004 13632
rect 106068 13568 106084 13632
rect 106148 13568 106164 13632
rect 106228 13568 106234 13632
rect 105918 13567 106234 13568
rect 4870 13088 5186 13089
rect 0 13018 800 13048
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 106654 13088 106970 13089
rect 106654 13024 106660 13088
rect 106724 13024 106740 13088
rect 106804 13024 106820 13088
rect 106884 13024 106900 13088
rect 106964 13024 106970 13088
rect 106654 13023 106970 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 105918 12544 106234 12545
rect 105918 12480 105924 12544
rect 105988 12480 106004 12544
rect 106068 12480 106084 12544
rect 106148 12480 106164 12544
rect 106228 12480 106234 12544
rect 105918 12479 106234 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 106654 12000 106970 12001
rect 106654 11936 106660 12000
rect 106724 11936 106740 12000
rect 106804 11936 106820 12000
rect 106884 11936 106900 12000
rect 106964 11936 106970 12000
rect 106654 11935 106970 11936
rect 0 11658 800 11688
rect 1209 11658 1275 11661
rect 0 11656 1275 11658
rect 0 11600 1214 11656
rect 1270 11600 1275 11656
rect 0 11598 1275 11600
rect 0 11568 800 11598
rect 1209 11595 1275 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 105918 11456 106234 11457
rect 105918 11392 105924 11456
rect 105988 11392 106004 11456
rect 106068 11392 106084 11456
rect 106148 11392 106164 11456
rect 106228 11392 106234 11456
rect 105918 11391 106234 11392
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 106654 10912 106970 10913
rect 106654 10848 106660 10912
rect 106724 10848 106740 10912
rect 106804 10848 106820 10912
rect 106884 10848 106900 10912
rect 106964 10848 106970 10912
rect 106654 10847 106970 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 105918 10368 106234 10369
rect 105918 10304 105924 10368
rect 105988 10304 106004 10368
rect 106068 10304 106084 10368
rect 106148 10304 106164 10368
rect 106228 10304 106234 10368
rect 105918 10303 106234 10304
rect 1301 10298 1367 10301
rect 0 10296 1367 10298
rect 0 10240 1306 10296
rect 1362 10240 1367 10296
rect 0 10238 1367 10240
rect 0 10208 800 10238
rect 1301 10235 1367 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 106654 9824 106970 9825
rect 106654 9760 106660 9824
rect 106724 9760 106740 9824
rect 106804 9760 106820 9824
rect 106884 9760 106900 9824
rect 106964 9760 106970 9824
rect 106654 9759 106970 9760
rect 23473 9756 23539 9757
rect 25773 9756 25839 9757
rect 28165 9756 28231 9757
rect 23432 9692 23438 9756
rect 23502 9754 23539 9756
rect 25768 9754 25774 9756
rect 23502 9752 23594 9754
rect 23534 9696 23594 9752
rect 23502 9694 23594 9696
rect 25686 9694 25774 9754
rect 23502 9692 23539 9694
rect 25768 9692 25774 9694
rect 25838 9692 25844 9756
rect 28114 9692 28120 9756
rect 28184 9754 28231 9756
rect 28184 9752 28276 9754
rect 28226 9696 28276 9752
rect 28184 9694 28276 9696
rect 28184 9692 28231 9694
rect 29272 9692 29278 9756
rect 29342 9754 29348 9756
rect 29545 9754 29611 9757
rect 30465 9756 30531 9757
rect 29342 9752 29611 9754
rect 29342 9696 29550 9752
rect 29606 9696 29611 9752
rect 29342 9694 29611 9696
rect 29342 9692 29348 9694
rect 23473 9691 23539 9692
rect 25773 9691 25839 9692
rect 28165 9691 28231 9692
rect 29545 9691 29611 9694
rect 30440 9692 30446 9756
rect 30510 9754 30531 9756
rect 30510 9752 30602 9754
rect 30526 9696 30602 9752
rect 30510 9694 30602 9696
rect 30510 9692 30531 9694
rect 30465 9691 30531 9692
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 16021 9620 16087 9621
rect 24669 9620 24735 9621
rect 16021 9616 16058 9620
rect 16122 9618 16128 9620
rect 24618 9618 24624 9620
rect 16021 9560 16026 9616
rect 16021 9556 16058 9560
rect 16122 9558 16178 9618
rect 24578 9558 24624 9618
rect 24688 9616 24735 9620
rect 90633 9620 90699 9621
rect 90817 9620 90883 9621
rect 90633 9618 90665 9620
rect 24730 9560 24735 9616
rect 16122 9556 16128 9558
rect 24618 9556 24624 9558
rect 24688 9556 24735 9560
rect 90573 9616 90665 9618
rect 90573 9560 90638 9616
rect 90573 9558 90665 9560
rect 16021 9555 16087 9556
rect 24669 9555 24735 9556
rect 90633 9556 90665 9558
rect 90729 9556 90735 9620
rect 90808 9556 90814 9620
rect 90878 9618 90884 9620
rect 90878 9558 90970 9618
rect 90878 9556 90884 9558
rect 90633 9555 90699 9556
rect 90817 9555 90883 9556
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 105918 9280 106234 9281
rect 105918 9216 105924 9280
rect 105988 9216 106004 9280
rect 106068 9216 106084 9280
rect 106148 9216 106164 9280
rect 106228 9216 106234 9280
rect 105918 9215 106234 9216
rect 0 8938 800 8968
rect 1209 8938 1275 8941
rect 0 8936 1275 8938
rect 0 8880 1214 8936
rect 1270 8880 1275 8936
rect 0 8878 1275 8880
rect 0 8848 800 8878
rect 1209 8875 1275 8878
rect 26693 8938 26759 8941
rect 26918 8938 26924 8940
rect 26693 8936 26924 8938
rect 26693 8880 26698 8936
rect 26754 8880 26924 8936
rect 26693 8878 26924 8880
rect 26693 8875 26759 8878
rect 26918 8876 26924 8878
rect 26988 8876 26994 8940
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 106654 8736 106970 8737
rect 106654 8672 106660 8736
rect 106724 8672 106740 8736
rect 106804 8672 106820 8736
rect 106884 8672 106900 8736
rect 106964 8672 106970 8736
rect 106654 8671 106970 8672
rect 90398 8332 90404 8396
rect 90468 8394 90474 8396
rect 90541 8394 90607 8397
rect 90468 8392 90607 8394
rect 90468 8336 90546 8392
rect 90602 8336 90607 8392
rect 90468 8334 90607 8336
rect 90468 8332 90474 8334
rect 90541 8331 90607 8334
rect 0 8258 800 8288
rect 1945 8258 2011 8261
rect 31661 8260 31727 8261
rect 31661 8258 31708 8260
rect 0 8256 2011 8258
rect 0 8200 1950 8256
rect 2006 8200 2011 8256
rect 0 8198 2011 8200
rect 31616 8256 31708 8258
rect 31616 8200 31666 8256
rect 31616 8198 31708 8200
rect 0 8168 800 8198
rect 1945 8195 2011 8198
rect 31661 8196 31708 8198
rect 31772 8196 31778 8260
rect 32806 8196 32812 8260
rect 32876 8258 32882 8260
rect 32949 8258 33015 8261
rect 32876 8256 33015 8258
rect 32876 8200 32954 8256
rect 33010 8200 33015 8256
rect 32876 8198 33015 8200
rect 32876 8196 32882 8198
rect 31661 8195 31727 8196
rect 32949 8195 33015 8198
rect 33910 8196 33916 8260
rect 33980 8258 33986 8260
rect 34237 8258 34303 8261
rect 33980 8256 34303 8258
rect 33980 8200 34242 8256
rect 34298 8200 34303 8256
rect 33980 8198 34303 8200
rect 33980 8196 33986 8198
rect 34237 8195 34303 8198
rect 35198 8196 35204 8260
rect 35268 8258 35274 8260
rect 35433 8258 35499 8261
rect 36353 8260 36419 8261
rect 37457 8260 37523 8261
rect 38745 8260 38811 8261
rect 36302 8258 36308 8260
rect 35268 8256 35499 8258
rect 35268 8200 35438 8256
rect 35494 8200 35499 8256
rect 35268 8198 35499 8200
rect 36262 8198 36308 8258
rect 36372 8256 36419 8260
rect 37406 8258 37412 8260
rect 36414 8200 36419 8256
rect 35268 8196 35274 8198
rect 35433 8195 35499 8198
rect 36302 8196 36308 8198
rect 36372 8196 36419 8200
rect 37366 8198 37412 8258
rect 37476 8256 37523 8260
rect 38694 8258 38700 8260
rect 37518 8200 37523 8256
rect 37406 8196 37412 8198
rect 37476 8196 37523 8200
rect 38654 8198 38700 8258
rect 38764 8256 38811 8260
rect 38806 8200 38811 8256
rect 38694 8196 38700 8198
rect 38764 8196 38811 8200
rect 40902 8196 40908 8260
rect 40972 8258 40978 8260
rect 41321 8258 41387 8261
rect 40972 8256 41387 8258
rect 40972 8200 41326 8256
rect 41382 8200 41387 8256
rect 40972 8198 41387 8200
rect 40972 8196 40978 8198
rect 36353 8195 36419 8196
rect 37457 8195 37523 8196
rect 38745 8195 38811 8196
rect 41321 8195 41387 8198
rect 42149 8260 42215 8261
rect 42149 8256 42196 8260
rect 42260 8258 42266 8260
rect 42149 8200 42154 8256
rect 42149 8196 42196 8200
rect 42260 8198 42306 8258
rect 42260 8196 42266 8198
rect 43294 8196 43300 8260
rect 43364 8258 43370 8260
rect 43437 8258 43503 8261
rect 43364 8256 43503 8258
rect 43364 8200 43442 8256
rect 43498 8200 43503 8256
rect 43364 8198 43503 8200
rect 43364 8196 43370 8198
rect 42149 8195 42215 8196
rect 43437 8195 43503 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 105918 8192 106234 8193
rect 105918 8128 105924 8192
rect 105988 8128 106004 8192
rect 106068 8128 106084 8192
rect 106148 8128 106164 8192
rect 106228 8128 106234 8192
rect 105918 8127 106234 8128
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 66310 7648 66626 7649
rect 66310 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66626 7648
rect 66310 7583 66626 7584
rect 97030 7648 97346 7649
rect 97030 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97346 7648
rect 97030 7583 97346 7584
rect 106654 7648 106970 7649
rect 106654 7584 106660 7648
rect 106724 7584 106740 7648
rect 106804 7584 106820 7648
rect 106884 7584 106900 7648
rect 106964 7584 106970 7648
rect 106654 7583 106970 7584
rect 1301 7578 1367 7581
rect 0 7576 1367 7578
rect 0 7520 1306 7576
rect 1362 7520 1367 7576
rect 0 7518 1367 7520
rect 0 7488 800 7518
rect 1301 7515 1367 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 96370 7104 96686 7105
rect 96370 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96686 7104
rect 96370 7039 96686 7040
rect 105918 7104 106234 7105
rect 105918 7040 105924 7104
rect 105988 7040 106004 7104
rect 106068 7040 106084 7104
rect 106148 7040 106164 7104
rect 106228 7040 106234 7104
rect 105918 7039 106234 7040
rect 0 6898 800 6928
rect 1301 6898 1367 6901
rect 0 6896 1367 6898
rect 0 6840 1306 6896
rect 1362 6840 1367 6896
rect 0 6838 1367 6840
rect 0 6808 800 6838
rect 1301 6835 1367 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 66310 6560 66626 6561
rect 66310 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66626 6560
rect 66310 6495 66626 6496
rect 97030 6560 97346 6561
rect 97030 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97346 6560
rect 97030 6495 97346 6496
rect 0 6218 800 6248
rect 1209 6218 1275 6221
rect 0 6216 1275 6218
rect 0 6160 1214 6216
rect 1270 6160 1275 6216
rect 0 6158 1275 6160
rect 0 6128 800 6158
rect 1209 6155 1275 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 96370 6016 96686 6017
rect 96370 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96686 6016
rect 96370 5951 96686 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 66310 5472 66626 5473
rect 66310 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66626 5472
rect 66310 5407 66626 5408
rect 97030 5472 97346 5473
rect 97030 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97346 5472
rect 97030 5407 97346 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 96370 4928 96686 4929
rect 96370 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96686 4928
rect 96370 4863 96686 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 39798 4524 39804 4588
rect 39868 4586 39874 4588
rect 39941 4586 40007 4589
rect 39868 4584 40007 4586
rect 39868 4528 39946 4584
rect 40002 4528 40007 4584
rect 39868 4526 40007 4528
rect 39868 4524 39874 4526
rect 39941 4523 40007 4526
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 66310 4384 66626 4385
rect 66310 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66626 4384
rect 66310 4319 66626 4320
rect 97030 4384 97346 4385
rect 97030 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97346 4384
rect 97030 4319 97346 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 96370 3840 96686 3841
rect 96370 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96686 3840
rect 96370 3775 96686 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 66310 3296 66626 3297
rect 66310 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66626 3296
rect 66310 3231 66626 3232
rect 97030 3296 97346 3297
rect 97030 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97346 3296
rect 97030 3231 97346 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 96370 2752 96686 2753
rect 96370 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96686 2752
rect 96370 2687 96686 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 66310 2208 66626 2209
rect 66310 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66626 2208
rect 66310 2143 66626 2144
rect 97030 2208 97346 2209
rect 97030 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97346 2208
rect 97030 2143 97346 2144
<< via3 >>
rect 4216 147452 4280 147456
rect 4216 147396 4220 147452
rect 4220 147396 4276 147452
rect 4276 147396 4280 147452
rect 4216 147392 4280 147396
rect 4296 147452 4360 147456
rect 4296 147396 4300 147452
rect 4300 147396 4356 147452
rect 4356 147396 4360 147452
rect 4296 147392 4360 147396
rect 4376 147452 4440 147456
rect 4376 147396 4380 147452
rect 4380 147396 4436 147452
rect 4436 147396 4440 147452
rect 4376 147392 4440 147396
rect 4456 147452 4520 147456
rect 4456 147396 4460 147452
rect 4460 147396 4516 147452
rect 4516 147396 4520 147452
rect 4456 147392 4520 147396
rect 34936 147452 35000 147456
rect 34936 147396 34940 147452
rect 34940 147396 34996 147452
rect 34996 147396 35000 147452
rect 34936 147392 35000 147396
rect 35016 147452 35080 147456
rect 35016 147396 35020 147452
rect 35020 147396 35076 147452
rect 35076 147396 35080 147452
rect 35016 147392 35080 147396
rect 35096 147452 35160 147456
rect 35096 147396 35100 147452
rect 35100 147396 35156 147452
rect 35156 147396 35160 147452
rect 35096 147392 35160 147396
rect 35176 147452 35240 147456
rect 35176 147396 35180 147452
rect 35180 147396 35236 147452
rect 35236 147396 35240 147452
rect 35176 147392 35240 147396
rect 65656 147452 65720 147456
rect 65656 147396 65660 147452
rect 65660 147396 65716 147452
rect 65716 147396 65720 147452
rect 65656 147392 65720 147396
rect 65736 147452 65800 147456
rect 65736 147396 65740 147452
rect 65740 147396 65796 147452
rect 65796 147396 65800 147452
rect 65736 147392 65800 147396
rect 65816 147452 65880 147456
rect 65816 147396 65820 147452
rect 65820 147396 65876 147452
rect 65876 147396 65880 147452
rect 65816 147392 65880 147396
rect 65896 147452 65960 147456
rect 65896 147396 65900 147452
rect 65900 147396 65956 147452
rect 65956 147396 65960 147452
rect 65896 147392 65960 147396
rect 96376 147452 96440 147456
rect 96376 147396 96380 147452
rect 96380 147396 96436 147452
rect 96436 147396 96440 147452
rect 96376 147392 96440 147396
rect 96456 147452 96520 147456
rect 96456 147396 96460 147452
rect 96460 147396 96516 147452
rect 96516 147396 96520 147452
rect 96456 147392 96520 147396
rect 96536 147452 96600 147456
rect 96536 147396 96540 147452
rect 96540 147396 96596 147452
rect 96596 147396 96600 147452
rect 96536 147392 96600 147396
rect 96616 147452 96680 147456
rect 96616 147396 96620 147452
rect 96620 147396 96676 147452
rect 96676 147396 96680 147452
rect 96616 147392 96680 147396
rect 4876 146908 4940 146912
rect 4876 146852 4880 146908
rect 4880 146852 4936 146908
rect 4936 146852 4940 146908
rect 4876 146848 4940 146852
rect 4956 146908 5020 146912
rect 4956 146852 4960 146908
rect 4960 146852 5016 146908
rect 5016 146852 5020 146908
rect 4956 146848 5020 146852
rect 5036 146908 5100 146912
rect 5036 146852 5040 146908
rect 5040 146852 5096 146908
rect 5096 146852 5100 146908
rect 5036 146848 5100 146852
rect 5116 146908 5180 146912
rect 5116 146852 5120 146908
rect 5120 146852 5176 146908
rect 5176 146852 5180 146908
rect 5116 146848 5180 146852
rect 35596 146908 35660 146912
rect 35596 146852 35600 146908
rect 35600 146852 35656 146908
rect 35656 146852 35660 146908
rect 35596 146848 35660 146852
rect 35676 146908 35740 146912
rect 35676 146852 35680 146908
rect 35680 146852 35736 146908
rect 35736 146852 35740 146908
rect 35676 146848 35740 146852
rect 35756 146908 35820 146912
rect 35756 146852 35760 146908
rect 35760 146852 35816 146908
rect 35816 146852 35820 146908
rect 35756 146848 35820 146852
rect 35836 146908 35900 146912
rect 35836 146852 35840 146908
rect 35840 146852 35896 146908
rect 35896 146852 35900 146908
rect 35836 146848 35900 146852
rect 66316 146908 66380 146912
rect 66316 146852 66320 146908
rect 66320 146852 66376 146908
rect 66376 146852 66380 146908
rect 66316 146848 66380 146852
rect 66396 146908 66460 146912
rect 66396 146852 66400 146908
rect 66400 146852 66456 146908
rect 66456 146852 66460 146908
rect 66396 146848 66460 146852
rect 66476 146908 66540 146912
rect 66476 146852 66480 146908
rect 66480 146852 66536 146908
rect 66536 146852 66540 146908
rect 66476 146848 66540 146852
rect 66556 146908 66620 146912
rect 66556 146852 66560 146908
rect 66560 146852 66616 146908
rect 66616 146852 66620 146908
rect 66556 146848 66620 146852
rect 97036 146908 97100 146912
rect 97036 146852 97040 146908
rect 97040 146852 97096 146908
rect 97096 146852 97100 146908
rect 97036 146848 97100 146852
rect 97116 146908 97180 146912
rect 97116 146852 97120 146908
rect 97120 146852 97176 146908
rect 97176 146852 97180 146908
rect 97116 146848 97180 146852
rect 97196 146908 97260 146912
rect 97196 146852 97200 146908
rect 97200 146852 97256 146908
rect 97256 146852 97260 146908
rect 97196 146848 97260 146852
rect 97276 146908 97340 146912
rect 97276 146852 97280 146908
rect 97280 146852 97336 146908
rect 97336 146852 97340 146908
rect 97276 146848 97340 146852
rect 4216 146364 4280 146368
rect 4216 146308 4220 146364
rect 4220 146308 4276 146364
rect 4276 146308 4280 146364
rect 4216 146304 4280 146308
rect 4296 146364 4360 146368
rect 4296 146308 4300 146364
rect 4300 146308 4356 146364
rect 4356 146308 4360 146364
rect 4296 146304 4360 146308
rect 4376 146364 4440 146368
rect 4376 146308 4380 146364
rect 4380 146308 4436 146364
rect 4436 146308 4440 146364
rect 4376 146304 4440 146308
rect 4456 146364 4520 146368
rect 4456 146308 4460 146364
rect 4460 146308 4516 146364
rect 4516 146308 4520 146364
rect 4456 146304 4520 146308
rect 34936 146364 35000 146368
rect 34936 146308 34940 146364
rect 34940 146308 34996 146364
rect 34996 146308 35000 146364
rect 34936 146304 35000 146308
rect 35016 146364 35080 146368
rect 35016 146308 35020 146364
rect 35020 146308 35076 146364
rect 35076 146308 35080 146364
rect 35016 146304 35080 146308
rect 35096 146364 35160 146368
rect 35096 146308 35100 146364
rect 35100 146308 35156 146364
rect 35156 146308 35160 146364
rect 35096 146304 35160 146308
rect 35176 146364 35240 146368
rect 35176 146308 35180 146364
rect 35180 146308 35236 146364
rect 35236 146308 35240 146364
rect 35176 146304 35240 146308
rect 65656 146364 65720 146368
rect 65656 146308 65660 146364
rect 65660 146308 65716 146364
rect 65716 146308 65720 146364
rect 65656 146304 65720 146308
rect 65736 146364 65800 146368
rect 65736 146308 65740 146364
rect 65740 146308 65796 146364
rect 65796 146308 65800 146364
rect 65736 146304 65800 146308
rect 65816 146364 65880 146368
rect 65816 146308 65820 146364
rect 65820 146308 65876 146364
rect 65876 146308 65880 146364
rect 65816 146304 65880 146308
rect 65896 146364 65960 146368
rect 65896 146308 65900 146364
rect 65900 146308 65956 146364
rect 65956 146308 65960 146364
rect 65896 146304 65960 146308
rect 96376 146364 96440 146368
rect 96376 146308 96380 146364
rect 96380 146308 96436 146364
rect 96436 146308 96440 146364
rect 96376 146304 96440 146308
rect 96456 146364 96520 146368
rect 96456 146308 96460 146364
rect 96460 146308 96516 146364
rect 96516 146308 96520 146364
rect 96456 146304 96520 146308
rect 96536 146364 96600 146368
rect 96536 146308 96540 146364
rect 96540 146308 96596 146364
rect 96596 146308 96600 146364
rect 96536 146304 96600 146308
rect 96616 146364 96680 146368
rect 96616 146308 96620 146364
rect 96620 146308 96676 146364
rect 96676 146308 96680 146364
rect 96616 146304 96680 146308
rect 4876 145820 4940 145824
rect 4876 145764 4880 145820
rect 4880 145764 4936 145820
rect 4936 145764 4940 145820
rect 4876 145760 4940 145764
rect 4956 145820 5020 145824
rect 4956 145764 4960 145820
rect 4960 145764 5016 145820
rect 5016 145764 5020 145820
rect 4956 145760 5020 145764
rect 5036 145820 5100 145824
rect 5036 145764 5040 145820
rect 5040 145764 5096 145820
rect 5096 145764 5100 145820
rect 5036 145760 5100 145764
rect 5116 145820 5180 145824
rect 5116 145764 5120 145820
rect 5120 145764 5176 145820
rect 5176 145764 5180 145820
rect 5116 145760 5180 145764
rect 35596 145820 35660 145824
rect 35596 145764 35600 145820
rect 35600 145764 35656 145820
rect 35656 145764 35660 145820
rect 35596 145760 35660 145764
rect 35676 145820 35740 145824
rect 35676 145764 35680 145820
rect 35680 145764 35736 145820
rect 35736 145764 35740 145820
rect 35676 145760 35740 145764
rect 35756 145820 35820 145824
rect 35756 145764 35760 145820
rect 35760 145764 35816 145820
rect 35816 145764 35820 145820
rect 35756 145760 35820 145764
rect 35836 145820 35900 145824
rect 35836 145764 35840 145820
rect 35840 145764 35896 145820
rect 35896 145764 35900 145820
rect 35836 145760 35900 145764
rect 66316 145820 66380 145824
rect 66316 145764 66320 145820
rect 66320 145764 66376 145820
rect 66376 145764 66380 145820
rect 66316 145760 66380 145764
rect 66396 145820 66460 145824
rect 66396 145764 66400 145820
rect 66400 145764 66456 145820
rect 66456 145764 66460 145820
rect 66396 145760 66460 145764
rect 66476 145820 66540 145824
rect 66476 145764 66480 145820
rect 66480 145764 66536 145820
rect 66536 145764 66540 145820
rect 66476 145760 66540 145764
rect 66556 145820 66620 145824
rect 66556 145764 66560 145820
rect 66560 145764 66616 145820
rect 66616 145764 66620 145820
rect 66556 145760 66620 145764
rect 97036 145820 97100 145824
rect 97036 145764 97040 145820
rect 97040 145764 97096 145820
rect 97096 145764 97100 145820
rect 97036 145760 97100 145764
rect 97116 145820 97180 145824
rect 97116 145764 97120 145820
rect 97120 145764 97176 145820
rect 97176 145764 97180 145820
rect 97116 145760 97180 145764
rect 97196 145820 97260 145824
rect 97196 145764 97200 145820
rect 97200 145764 97256 145820
rect 97256 145764 97260 145820
rect 97196 145760 97260 145764
rect 97276 145820 97340 145824
rect 97276 145764 97280 145820
rect 97280 145764 97336 145820
rect 97336 145764 97340 145820
rect 97276 145760 97340 145764
rect 4216 145276 4280 145280
rect 4216 145220 4220 145276
rect 4220 145220 4276 145276
rect 4276 145220 4280 145276
rect 4216 145216 4280 145220
rect 4296 145276 4360 145280
rect 4296 145220 4300 145276
rect 4300 145220 4356 145276
rect 4356 145220 4360 145276
rect 4296 145216 4360 145220
rect 4376 145276 4440 145280
rect 4376 145220 4380 145276
rect 4380 145220 4436 145276
rect 4436 145220 4440 145276
rect 4376 145216 4440 145220
rect 4456 145276 4520 145280
rect 4456 145220 4460 145276
rect 4460 145220 4516 145276
rect 4516 145220 4520 145276
rect 4456 145216 4520 145220
rect 34936 145276 35000 145280
rect 34936 145220 34940 145276
rect 34940 145220 34996 145276
rect 34996 145220 35000 145276
rect 34936 145216 35000 145220
rect 35016 145276 35080 145280
rect 35016 145220 35020 145276
rect 35020 145220 35076 145276
rect 35076 145220 35080 145276
rect 35016 145216 35080 145220
rect 35096 145276 35160 145280
rect 35096 145220 35100 145276
rect 35100 145220 35156 145276
rect 35156 145220 35160 145276
rect 35096 145216 35160 145220
rect 35176 145276 35240 145280
rect 35176 145220 35180 145276
rect 35180 145220 35236 145276
rect 35236 145220 35240 145276
rect 35176 145216 35240 145220
rect 65656 145276 65720 145280
rect 65656 145220 65660 145276
rect 65660 145220 65716 145276
rect 65716 145220 65720 145276
rect 65656 145216 65720 145220
rect 65736 145276 65800 145280
rect 65736 145220 65740 145276
rect 65740 145220 65796 145276
rect 65796 145220 65800 145276
rect 65736 145216 65800 145220
rect 65816 145276 65880 145280
rect 65816 145220 65820 145276
rect 65820 145220 65876 145276
rect 65876 145220 65880 145276
rect 65816 145216 65880 145220
rect 65896 145276 65960 145280
rect 65896 145220 65900 145276
rect 65900 145220 65956 145276
rect 65956 145220 65960 145276
rect 65896 145216 65960 145220
rect 96376 145276 96440 145280
rect 96376 145220 96380 145276
rect 96380 145220 96436 145276
rect 96436 145220 96440 145276
rect 96376 145216 96440 145220
rect 96456 145276 96520 145280
rect 96456 145220 96460 145276
rect 96460 145220 96516 145276
rect 96516 145220 96520 145276
rect 96456 145216 96520 145220
rect 96536 145276 96600 145280
rect 96536 145220 96540 145276
rect 96540 145220 96596 145276
rect 96596 145220 96600 145276
rect 96536 145216 96600 145220
rect 96616 145276 96680 145280
rect 96616 145220 96620 145276
rect 96620 145220 96676 145276
rect 96676 145220 96680 145276
rect 96616 145216 96680 145220
rect 4876 144732 4940 144736
rect 4876 144676 4880 144732
rect 4880 144676 4936 144732
rect 4936 144676 4940 144732
rect 4876 144672 4940 144676
rect 4956 144732 5020 144736
rect 4956 144676 4960 144732
rect 4960 144676 5016 144732
rect 5016 144676 5020 144732
rect 4956 144672 5020 144676
rect 5036 144732 5100 144736
rect 5036 144676 5040 144732
rect 5040 144676 5096 144732
rect 5096 144676 5100 144732
rect 5036 144672 5100 144676
rect 5116 144732 5180 144736
rect 5116 144676 5120 144732
rect 5120 144676 5176 144732
rect 5176 144676 5180 144732
rect 5116 144672 5180 144676
rect 35596 144732 35660 144736
rect 35596 144676 35600 144732
rect 35600 144676 35656 144732
rect 35656 144676 35660 144732
rect 35596 144672 35660 144676
rect 35676 144732 35740 144736
rect 35676 144676 35680 144732
rect 35680 144676 35736 144732
rect 35736 144676 35740 144732
rect 35676 144672 35740 144676
rect 35756 144732 35820 144736
rect 35756 144676 35760 144732
rect 35760 144676 35816 144732
rect 35816 144676 35820 144732
rect 35756 144672 35820 144676
rect 35836 144732 35900 144736
rect 35836 144676 35840 144732
rect 35840 144676 35896 144732
rect 35896 144676 35900 144732
rect 35836 144672 35900 144676
rect 66316 144732 66380 144736
rect 66316 144676 66320 144732
rect 66320 144676 66376 144732
rect 66376 144676 66380 144732
rect 66316 144672 66380 144676
rect 66396 144732 66460 144736
rect 66396 144676 66400 144732
rect 66400 144676 66456 144732
rect 66456 144676 66460 144732
rect 66396 144672 66460 144676
rect 66476 144732 66540 144736
rect 66476 144676 66480 144732
rect 66480 144676 66536 144732
rect 66536 144676 66540 144732
rect 66476 144672 66540 144676
rect 66556 144732 66620 144736
rect 66556 144676 66560 144732
rect 66560 144676 66616 144732
rect 66616 144676 66620 144732
rect 66556 144672 66620 144676
rect 97036 144732 97100 144736
rect 97036 144676 97040 144732
rect 97040 144676 97096 144732
rect 97096 144676 97100 144732
rect 97036 144672 97100 144676
rect 97116 144732 97180 144736
rect 97116 144676 97120 144732
rect 97120 144676 97176 144732
rect 97176 144676 97180 144732
rect 97116 144672 97180 144676
rect 97196 144732 97260 144736
rect 97196 144676 97200 144732
rect 97200 144676 97256 144732
rect 97256 144676 97260 144732
rect 97196 144672 97260 144676
rect 97276 144732 97340 144736
rect 97276 144676 97280 144732
rect 97280 144676 97336 144732
rect 97336 144676 97340 144732
rect 97276 144672 97340 144676
rect 4216 144188 4280 144192
rect 4216 144132 4220 144188
rect 4220 144132 4276 144188
rect 4276 144132 4280 144188
rect 4216 144128 4280 144132
rect 4296 144188 4360 144192
rect 4296 144132 4300 144188
rect 4300 144132 4356 144188
rect 4356 144132 4360 144188
rect 4296 144128 4360 144132
rect 4376 144188 4440 144192
rect 4376 144132 4380 144188
rect 4380 144132 4436 144188
rect 4436 144132 4440 144188
rect 4376 144128 4440 144132
rect 4456 144188 4520 144192
rect 4456 144132 4460 144188
rect 4460 144132 4516 144188
rect 4516 144132 4520 144188
rect 4456 144128 4520 144132
rect 34936 144188 35000 144192
rect 34936 144132 34940 144188
rect 34940 144132 34996 144188
rect 34996 144132 35000 144188
rect 34936 144128 35000 144132
rect 35016 144188 35080 144192
rect 35016 144132 35020 144188
rect 35020 144132 35076 144188
rect 35076 144132 35080 144188
rect 35016 144128 35080 144132
rect 35096 144188 35160 144192
rect 35096 144132 35100 144188
rect 35100 144132 35156 144188
rect 35156 144132 35160 144188
rect 35096 144128 35160 144132
rect 35176 144188 35240 144192
rect 35176 144132 35180 144188
rect 35180 144132 35236 144188
rect 35236 144132 35240 144188
rect 35176 144128 35240 144132
rect 65656 144188 65720 144192
rect 65656 144132 65660 144188
rect 65660 144132 65716 144188
rect 65716 144132 65720 144188
rect 65656 144128 65720 144132
rect 65736 144188 65800 144192
rect 65736 144132 65740 144188
rect 65740 144132 65796 144188
rect 65796 144132 65800 144188
rect 65736 144128 65800 144132
rect 65816 144188 65880 144192
rect 65816 144132 65820 144188
rect 65820 144132 65876 144188
rect 65876 144132 65880 144188
rect 65816 144128 65880 144132
rect 65896 144188 65960 144192
rect 65896 144132 65900 144188
rect 65900 144132 65956 144188
rect 65956 144132 65960 144188
rect 65896 144128 65960 144132
rect 96376 144188 96440 144192
rect 96376 144132 96380 144188
rect 96380 144132 96436 144188
rect 96436 144132 96440 144188
rect 96376 144128 96440 144132
rect 96456 144188 96520 144192
rect 96456 144132 96460 144188
rect 96460 144132 96516 144188
rect 96516 144132 96520 144188
rect 96456 144128 96520 144132
rect 96536 144188 96600 144192
rect 96536 144132 96540 144188
rect 96540 144132 96596 144188
rect 96596 144132 96600 144188
rect 96536 144128 96600 144132
rect 96616 144188 96680 144192
rect 96616 144132 96620 144188
rect 96620 144132 96676 144188
rect 96676 144132 96680 144188
rect 96616 144128 96680 144132
rect 4876 143644 4940 143648
rect 4876 143588 4880 143644
rect 4880 143588 4936 143644
rect 4936 143588 4940 143644
rect 4876 143584 4940 143588
rect 4956 143644 5020 143648
rect 4956 143588 4960 143644
rect 4960 143588 5016 143644
rect 5016 143588 5020 143644
rect 4956 143584 5020 143588
rect 5036 143644 5100 143648
rect 5036 143588 5040 143644
rect 5040 143588 5096 143644
rect 5096 143588 5100 143644
rect 5036 143584 5100 143588
rect 5116 143644 5180 143648
rect 5116 143588 5120 143644
rect 5120 143588 5176 143644
rect 5176 143588 5180 143644
rect 5116 143584 5180 143588
rect 35596 143644 35660 143648
rect 35596 143588 35600 143644
rect 35600 143588 35656 143644
rect 35656 143588 35660 143644
rect 35596 143584 35660 143588
rect 35676 143644 35740 143648
rect 35676 143588 35680 143644
rect 35680 143588 35736 143644
rect 35736 143588 35740 143644
rect 35676 143584 35740 143588
rect 35756 143644 35820 143648
rect 35756 143588 35760 143644
rect 35760 143588 35816 143644
rect 35816 143588 35820 143644
rect 35756 143584 35820 143588
rect 35836 143644 35900 143648
rect 35836 143588 35840 143644
rect 35840 143588 35896 143644
rect 35896 143588 35900 143644
rect 35836 143584 35900 143588
rect 66316 143644 66380 143648
rect 66316 143588 66320 143644
rect 66320 143588 66376 143644
rect 66376 143588 66380 143644
rect 66316 143584 66380 143588
rect 66396 143644 66460 143648
rect 66396 143588 66400 143644
rect 66400 143588 66456 143644
rect 66456 143588 66460 143644
rect 66396 143584 66460 143588
rect 66476 143644 66540 143648
rect 66476 143588 66480 143644
rect 66480 143588 66536 143644
rect 66536 143588 66540 143644
rect 66476 143584 66540 143588
rect 66556 143644 66620 143648
rect 66556 143588 66560 143644
rect 66560 143588 66616 143644
rect 66616 143588 66620 143644
rect 66556 143584 66620 143588
rect 97036 143644 97100 143648
rect 97036 143588 97040 143644
rect 97040 143588 97096 143644
rect 97096 143588 97100 143644
rect 97036 143584 97100 143588
rect 97116 143644 97180 143648
rect 97116 143588 97120 143644
rect 97120 143588 97176 143644
rect 97176 143588 97180 143644
rect 97116 143584 97180 143588
rect 97196 143644 97260 143648
rect 97196 143588 97200 143644
rect 97200 143588 97256 143644
rect 97256 143588 97260 143644
rect 97196 143584 97260 143588
rect 97276 143644 97340 143648
rect 97276 143588 97280 143644
rect 97280 143588 97336 143644
rect 97336 143588 97340 143644
rect 97276 143584 97340 143588
rect 4216 143100 4280 143104
rect 4216 143044 4220 143100
rect 4220 143044 4276 143100
rect 4276 143044 4280 143100
rect 4216 143040 4280 143044
rect 4296 143100 4360 143104
rect 4296 143044 4300 143100
rect 4300 143044 4356 143100
rect 4356 143044 4360 143100
rect 4296 143040 4360 143044
rect 4376 143100 4440 143104
rect 4376 143044 4380 143100
rect 4380 143044 4436 143100
rect 4436 143044 4440 143100
rect 4376 143040 4440 143044
rect 4456 143100 4520 143104
rect 4456 143044 4460 143100
rect 4460 143044 4516 143100
rect 4516 143044 4520 143100
rect 4456 143040 4520 143044
rect 34936 143100 35000 143104
rect 34936 143044 34940 143100
rect 34940 143044 34996 143100
rect 34996 143044 35000 143100
rect 34936 143040 35000 143044
rect 35016 143100 35080 143104
rect 35016 143044 35020 143100
rect 35020 143044 35076 143100
rect 35076 143044 35080 143100
rect 35016 143040 35080 143044
rect 35096 143100 35160 143104
rect 35096 143044 35100 143100
rect 35100 143044 35156 143100
rect 35156 143044 35160 143100
rect 35096 143040 35160 143044
rect 35176 143100 35240 143104
rect 35176 143044 35180 143100
rect 35180 143044 35236 143100
rect 35236 143044 35240 143100
rect 35176 143040 35240 143044
rect 65656 143100 65720 143104
rect 65656 143044 65660 143100
rect 65660 143044 65716 143100
rect 65716 143044 65720 143100
rect 65656 143040 65720 143044
rect 65736 143100 65800 143104
rect 65736 143044 65740 143100
rect 65740 143044 65796 143100
rect 65796 143044 65800 143100
rect 65736 143040 65800 143044
rect 65816 143100 65880 143104
rect 65816 143044 65820 143100
rect 65820 143044 65876 143100
rect 65876 143044 65880 143100
rect 65816 143040 65880 143044
rect 65896 143100 65960 143104
rect 65896 143044 65900 143100
rect 65900 143044 65956 143100
rect 65956 143044 65960 143100
rect 65896 143040 65960 143044
rect 96376 143100 96440 143104
rect 96376 143044 96380 143100
rect 96380 143044 96436 143100
rect 96436 143044 96440 143100
rect 96376 143040 96440 143044
rect 96456 143100 96520 143104
rect 96456 143044 96460 143100
rect 96460 143044 96516 143100
rect 96516 143044 96520 143100
rect 96456 143040 96520 143044
rect 96536 143100 96600 143104
rect 96536 143044 96540 143100
rect 96540 143044 96596 143100
rect 96596 143044 96600 143100
rect 96536 143040 96600 143044
rect 96616 143100 96680 143104
rect 96616 143044 96620 143100
rect 96620 143044 96676 143100
rect 96676 143044 96680 143100
rect 96616 143040 96680 143044
rect 4876 142556 4940 142560
rect 4876 142500 4880 142556
rect 4880 142500 4936 142556
rect 4936 142500 4940 142556
rect 4876 142496 4940 142500
rect 4956 142556 5020 142560
rect 4956 142500 4960 142556
rect 4960 142500 5016 142556
rect 5016 142500 5020 142556
rect 4956 142496 5020 142500
rect 5036 142556 5100 142560
rect 5036 142500 5040 142556
rect 5040 142500 5096 142556
rect 5096 142500 5100 142556
rect 5036 142496 5100 142500
rect 5116 142556 5180 142560
rect 5116 142500 5120 142556
rect 5120 142500 5176 142556
rect 5176 142500 5180 142556
rect 5116 142496 5180 142500
rect 35596 142556 35660 142560
rect 35596 142500 35600 142556
rect 35600 142500 35656 142556
rect 35656 142500 35660 142556
rect 35596 142496 35660 142500
rect 35676 142556 35740 142560
rect 35676 142500 35680 142556
rect 35680 142500 35736 142556
rect 35736 142500 35740 142556
rect 35676 142496 35740 142500
rect 35756 142556 35820 142560
rect 35756 142500 35760 142556
rect 35760 142500 35816 142556
rect 35816 142500 35820 142556
rect 35756 142496 35820 142500
rect 35836 142556 35900 142560
rect 35836 142500 35840 142556
rect 35840 142500 35896 142556
rect 35896 142500 35900 142556
rect 35836 142496 35900 142500
rect 66316 142556 66380 142560
rect 66316 142500 66320 142556
rect 66320 142500 66376 142556
rect 66376 142500 66380 142556
rect 66316 142496 66380 142500
rect 66396 142556 66460 142560
rect 66396 142500 66400 142556
rect 66400 142500 66456 142556
rect 66456 142500 66460 142556
rect 66396 142496 66460 142500
rect 66476 142556 66540 142560
rect 66476 142500 66480 142556
rect 66480 142500 66536 142556
rect 66536 142500 66540 142556
rect 66476 142496 66540 142500
rect 66556 142556 66620 142560
rect 66556 142500 66560 142556
rect 66560 142500 66616 142556
rect 66616 142500 66620 142556
rect 66556 142496 66620 142500
rect 97036 142556 97100 142560
rect 97036 142500 97040 142556
rect 97040 142500 97096 142556
rect 97096 142500 97100 142556
rect 97036 142496 97100 142500
rect 97116 142556 97180 142560
rect 97116 142500 97120 142556
rect 97120 142500 97176 142556
rect 97176 142500 97180 142556
rect 97116 142496 97180 142500
rect 97196 142556 97260 142560
rect 97196 142500 97200 142556
rect 97200 142500 97256 142556
rect 97256 142500 97260 142556
rect 97196 142496 97260 142500
rect 97276 142556 97340 142560
rect 97276 142500 97280 142556
rect 97280 142500 97336 142556
rect 97336 142500 97340 142556
rect 97276 142496 97340 142500
rect 4216 142012 4280 142016
rect 4216 141956 4220 142012
rect 4220 141956 4276 142012
rect 4276 141956 4280 142012
rect 4216 141952 4280 141956
rect 4296 142012 4360 142016
rect 4296 141956 4300 142012
rect 4300 141956 4356 142012
rect 4356 141956 4360 142012
rect 4296 141952 4360 141956
rect 4376 142012 4440 142016
rect 4376 141956 4380 142012
rect 4380 141956 4436 142012
rect 4436 141956 4440 142012
rect 4376 141952 4440 141956
rect 4456 142012 4520 142016
rect 4456 141956 4460 142012
rect 4460 141956 4516 142012
rect 4516 141956 4520 142012
rect 4456 141952 4520 141956
rect 34936 142012 35000 142016
rect 34936 141956 34940 142012
rect 34940 141956 34996 142012
rect 34996 141956 35000 142012
rect 34936 141952 35000 141956
rect 35016 142012 35080 142016
rect 35016 141956 35020 142012
rect 35020 141956 35076 142012
rect 35076 141956 35080 142012
rect 35016 141952 35080 141956
rect 35096 142012 35160 142016
rect 35096 141956 35100 142012
rect 35100 141956 35156 142012
rect 35156 141956 35160 142012
rect 35096 141952 35160 141956
rect 35176 142012 35240 142016
rect 35176 141956 35180 142012
rect 35180 141956 35236 142012
rect 35236 141956 35240 142012
rect 35176 141952 35240 141956
rect 65656 142012 65720 142016
rect 65656 141956 65660 142012
rect 65660 141956 65716 142012
rect 65716 141956 65720 142012
rect 65656 141952 65720 141956
rect 65736 142012 65800 142016
rect 65736 141956 65740 142012
rect 65740 141956 65796 142012
rect 65796 141956 65800 142012
rect 65736 141952 65800 141956
rect 65816 142012 65880 142016
rect 65816 141956 65820 142012
rect 65820 141956 65876 142012
rect 65876 141956 65880 142012
rect 65816 141952 65880 141956
rect 65896 142012 65960 142016
rect 65896 141956 65900 142012
rect 65900 141956 65956 142012
rect 65956 141956 65960 142012
rect 65896 141952 65960 141956
rect 96376 142012 96440 142016
rect 96376 141956 96380 142012
rect 96380 141956 96436 142012
rect 96436 141956 96440 142012
rect 96376 141952 96440 141956
rect 96456 142012 96520 142016
rect 96456 141956 96460 142012
rect 96460 141956 96516 142012
rect 96516 141956 96520 142012
rect 96456 141952 96520 141956
rect 96536 142012 96600 142016
rect 96536 141956 96540 142012
rect 96540 141956 96596 142012
rect 96596 141956 96600 142012
rect 96536 141952 96600 141956
rect 96616 142012 96680 142016
rect 96616 141956 96620 142012
rect 96620 141956 96676 142012
rect 96676 141956 96680 142012
rect 96616 141952 96680 141956
rect 4876 141468 4940 141472
rect 4876 141412 4880 141468
rect 4880 141412 4936 141468
rect 4936 141412 4940 141468
rect 4876 141408 4940 141412
rect 4956 141468 5020 141472
rect 4956 141412 4960 141468
rect 4960 141412 5016 141468
rect 5016 141412 5020 141468
rect 4956 141408 5020 141412
rect 5036 141468 5100 141472
rect 5036 141412 5040 141468
rect 5040 141412 5096 141468
rect 5096 141412 5100 141468
rect 5036 141408 5100 141412
rect 5116 141468 5180 141472
rect 5116 141412 5120 141468
rect 5120 141412 5176 141468
rect 5176 141412 5180 141468
rect 5116 141408 5180 141412
rect 35596 141468 35660 141472
rect 35596 141412 35600 141468
rect 35600 141412 35656 141468
rect 35656 141412 35660 141468
rect 35596 141408 35660 141412
rect 35676 141468 35740 141472
rect 35676 141412 35680 141468
rect 35680 141412 35736 141468
rect 35736 141412 35740 141468
rect 35676 141408 35740 141412
rect 35756 141468 35820 141472
rect 35756 141412 35760 141468
rect 35760 141412 35816 141468
rect 35816 141412 35820 141468
rect 35756 141408 35820 141412
rect 35836 141468 35900 141472
rect 35836 141412 35840 141468
rect 35840 141412 35896 141468
rect 35896 141412 35900 141468
rect 35836 141408 35900 141412
rect 66316 141468 66380 141472
rect 66316 141412 66320 141468
rect 66320 141412 66376 141468
rect 66376 141412 66380 141468
rect 66316 141408 66380 141412
rect 66396 141468 66460 141472
rect 66396 141412 66400 141468
rect 66400 141412 66456 141468
rect 66456 141412 66460 141468
rect 66396 141408 66460 141412
rect 66476 141468 66540 141472
rect 66476 141412 66480 141468
rect 66480 141412 66536 141468
rect 66536 141412 66540 141468
rect 66476 141408 66540 141412
rect 66556 141468 66620 141472
rect 66556 141412 66560 141468
rect 66560 141412 66616 141468
rect 66616 141412 66620 141468
rect 66556 141408 66620 141412
rect 97036 141468 97100 141472
rect 97036 141412 97040 141468
rect 97040 141412 97096 141468
rect 97096 141412 97100 141468
rect 97036 141408 97100 141412
rect 97116 141468 97180 141472
rect 97116 141412 97120 141468
rect 97120 141412 97176 141468
rect 97176 141412 97180 141468
rect 97116 141408 97180 141412
rect 97196 141468 97260 141472
rect 97196 141412 97200 141468
rect 97200 141412 97256 141468
rect 97256 141412 97260 141468
rect 97196 141408 97260 141412
rect 97276 141468 97340 141472
rect 97276 141412 97280 141468
rect 97280 141412 97336 141468
rect 97336 141412 97340 141468
rect 97276 141408 97340 141412
rect 4216 140924 4280 140928
rect 4216 140868 4220 140924
rect 4220 140868 4276 140924
rect 4276 140868 4280 140924
rect 4216 140864 4280 140868
rect 4296 140924 4360 140928
rect 4296 140868 4300 140924
rect 4300 140868 4356 140924
rect 4356 140868 4360 140924
rect 4296 140864 4360 140868
rect 4376 140924 4440 140928
rect 4376 140868 4380 140924
rect 4380 140868 4436 140924
rect 4436 140868 4440 140924
rect 4376 140864 4440 140868
rect 4456 140924 4520 140928
rect 4456 140868 4460 140924
rect 4460 140868 4516 140924
rect 4516 140868 4520 140924
rect 4456 140864 4520 140868
rect 34936 140924 35000 140928
rect 34936 140868 34940 140924
rect 34940 140868 34996 140924
rect 34996 140868 35000 140924
rect 34936 140864 35000 140868
rect 35016 140924 35080 140928
rect 35016 140868 35020 140924
rect 35020 140868 35076 140924
rect 35076 140868 35080 140924
rect 35016 140864 35080 140868
rect 35096 140924 35160 140928
rect 35096 140868 35100 140924
rect 35100 140868 35156 140924
rect 35156 140868 35160 140924
rect 35096 140864 35160 140868
rect 35176 140924 35240 140928
rect 35176 140868 35180 140924
rect 35180 140868 35236 140924
rect 35236 140868 35240 140924
rect 35176 140864 35240 140868
rect 65656 140924 65720 140928
rect 65656 140868 65660 140924
rect 65660 140868 65716 140924
rect 65716 140868 65720 140924
rect 65656 140864 65720 140868
rect 65736 140924 65800 140928
rect 65736 140868 65740 140924
rect 65740 140868 65796 140924
rect 65796 140868 65800 140924
rect 65736 140864 65800 140868
rect 65816 140924 65880 140928
rect 65816 140868 65820 140924
rect 65820 140868 65876 140924
rect 65876 140868 65880 140924
rect 65816 140864 65880 140868
rect 65896 140924 65960 140928
rect 65896 140868 65900 140924
rect 65900 140868 65956 140924
rect 65956 140868 65960 140924
rect 65896 140864 65960 140868
rect 96376 140924 96440 140928
rect 96376 140868 96380 140924
rect 96380 140868 96436 140924
rect 96436 140868 96440 140924
rect 96376 140864 96440 140868
rect 96456 140924 96520 140928
rect 96456 140868 96460 140924
rect 96460 140868 96516 140924
rect 96516 140868 96520 140924
rect 96456 140864 96520 140868
rect 96536 140924 96600 140928
rect 96536 140868 96540 140924
rect 96540 140868 96596 140924
rect 96596 140868 96600 140924
rect 96536 140864 96600 140868
rect 96616 140924 96680 140928
rect 96616 140868 96620 140924
rect 96620 140868 96676 140924
rect 96676 140868 96680 140924
rect 96616 140864 96680 140868
rect 4876 140380 4940 140384
rect 4876 140324 4880 140380
rect 4880 140324 4936 140380
rect 4936 140324 4940 140380
rect 4876 140320 4940 140324
rect 4956 140380 5020 140384
rect 4956 140324 4960 140380
rect 4960 140324 5016 140380
rect 5016 140324 5020 140380
rect 4956 140320 5020 140324
rect 5036 140380 5100 140384
rect 5036 140324 5040 140380
rect 5040 140324 5096 140380
rect 5096 140324 5100 140380
rect 5036 140320 5100 140324
rect 5116 140380 5180 140384
rect 5116 140324 5120 140380
rect 5120 140324 5176 140380
rect 5176 140324 5180 140380
rect 5116 140320 5180 140324
rect 35596 140380 35660 140384
rect 35596 140324 35600 140380
rect 35600 140324 35656 140380
rect 35656 140324 35660 140380
rect 35596 140320 35660 140324
rect 35676 140380 35740 140384
rect 35676 140324 35680 140380
rect 35680 140324 35736 140380
rect 35736 140324 35740 140380
rect 35676 140320 35740 140324
rect 35756 140380 35820 140384
rect 35756 140324 35760 140380
rect 35760 140324 35816 140380
rect 35816 140324 35820 140380
rect 35756 140320 35820 140324
rect 35836 140380 35900 140384
rect 35836 140324 35840 140380
rect 35840 140324 35896 140380
rect 35896 140324 35900 140380
rect 35836 140320 35900 140324
rect 66316 140380 66380 140384
rect 66316 140324 66320 140380
rect 66320 140324 66376 140380
rect 66376 140324 66380 140380
rect 66316 140320 66380 140324
rect 66396 140380 66460 140384
rect 66396 140324 66400 140380
rect 66400 140324 66456 140380
rect 66456 140324 66460 140380
rect 66396 140320 66460 140324
rect 66476 140380 66540 140384
rect 66476 140324 66480 140380
rect 66480 140324 66536 140380
rect 66536 140324 66540 140380
rect 66476 140320 66540 140324
rect 66556 140380 66620 140384
rect 66556 140324 66560 140380
rect 66560 140324 66616 140380
rect 66616 140324 66620 140380
rect 66556 140320 66620 140324
rect 97036 140380 97100 140384
rect 97036 140324 97040 140380
rect 97040 140324 97096 140380
rect 97096 140324 97100 140380
rect 97036 140320 97100 140324
rect 97116 140380 97180 140384
rect 97116 140324 97120 140380
rect 97120 140324 97176 140380
rect 97176 140324 97180 140380
rect 97116 140320 97180 140324
rect 97196 140380 97260 140384
rect 97196 140324 97200 140380
rect 97200 140324 97256 140380
rect 97256 140324 97260 140380
rect 97196 140320 97260 140324
rect 97276 140380 97340 140384
rect 97276 140324 97280 140380
rect 97280 140324 97336 140380
rect 97336 140324 97340 140380
rect 97276 140320 97340 140324
rect 4216 139836 4280 139840
rect 4216 139780 4220 139836
rect 4220 139780 4276 139836
rect 4276 139780 4280 139836
rect 4216 139776 4280 139780
rect 4296 139836 4360 139840
rect 4296 139780 4300 139836
rect 4300 139780 4356 139836
rect 4356 139780 4360 139836
rect 4296 139776 4360 139780
rect 4376 139836 4440 139840
rect 4376 139780 4380 139836
rect 4380 139780 4436 139836
rect 4436 139780 4440 139836
rect 4376 139776 4440 139780
rect 4456 139836 4520 139840
rect 4456 139780 4460 139836
rect 4460 139780 4516 139836
rect 4516 139780 4520 139836
rect 4456 139776 4520 139780
rect 34936 139836 35000 139840
rect 34936 139780 34940 139836
rect 34940 139780 34996 139836
rect 34996 139780 35000 139836
rect 34936 139776 35000 139780
rect 35016 139836 35080 139840
rect 35016 139780 35020 139836
rect 35020 139780 35076 139836
rect 35076 139780 35080 139836
rect 35016 139776 35080 139780
rect 35096 139836 35160 139840
rect 35096 139780 35100 139836
rect 35100 139780 35156 139836
rect 35156 139780 35160 139836
rect 35096 139776 35160 139780
rect 35176 139836 35240 139840
rect 35176 139780 35180 139836
rect 35180 139780 35236 139836
rect 35236 139780 35240 139836
rect 35176 139776 35240 139780
rect 65656 139836 65720 139840
rect 65656 139780 65660 139836
rect 65660 139780 65716 139836
rect 65716 139780 65720 139836
rect 65656 139776 65720 139780
rect 65736 139836 65800 139840
rect 65736 139780 65740 139836
rect 65740 139780 65796 139836
rect 65796 139780 65800 139836
rect 65736 139776 65800 139780
rect 65816 139836 65880 139840
rect 65816 139780 65820 139836
rect 65820 139780 65876 139836
rect 65876 139780 65880 139836
rect 65816 139776 65880 139780
rect 65896 139836 65960 139840
rect 65896 139780 65900 139836
rect 65900 139780 65956 139836
rect 65956 139780 65960 139836
rect 65896 139776 65960 139780
rect 96376 139836 96440 139840
rect 96376 139780 96380 139836
rect 96380 139780 96436 139836
rect 96436 139780 96440 139836
rect 96376 139776 96440 139780
rect 96456 139836 96520 139840
rect 96456 139780 96460 139836
rect 96460 139780 96516 139836
rect 96516 139780 96520 139836
rect 96456 139776 96520 139780
rect 96536 139836 96600 139840
rect 96536 139780 96540 139836
rect 96540 139780 96596 139836
rect 96596 139780 96600 139836
rect 96536 139776 96600 139780
rect 96616 139836 96680 139840
rect 96616 139780 96620 139836
rect 96620 139780 96676 139836
rect 96676 139780 96680 139836
rect 96616 139776 96680 139780
rect 4876 139292 4940 139296
rect 4876 139236 4880 139292
rect 4880 139236 4936 139292
rect 4936 139236 4940 139292
rect 4876 139232 4940 139236
rect 4956 139292 5020 139296
rect 4956 139236 4960 139292
rect 4960 139236 5016 139292
rect 5016 139236 5020 139292
rect 4956 139232 5020 139236
rect 5036 139292 5100 139296
rect 5036 139236 5040 139292
rect 5040 139236 5096 139292
rect 5096 139236 5100 139292
rect 5036 139232 5100 139236
rect 5116 139292 5180 139296
rect 5116 139236 5120 139292
rect 5120 139236 5176 139292
rect 5176 139236 5180 139292
rect 5116 139232 5180 139236
rect 35596 139292 35660 139296
rect 35596 139236 35600 139292
rect 35600 139236 35656 139292
rect 35656 139236 35660 139292
rect 35596 139232 35660 139236
rect 35676 139292 35740 139296
rect 35676 139236 35680 139292
rect 35680 139236 35736 139292
rect 35736 139236 35740 139292
rect 35676 139232 35740 139236
rect 35756 139292 35820 139296
rect 35756 139236 35760 139292
rect 35760 139236 35816 139292
rect 35816 139236 35820 139292
rect 35756 139232 35820 139236
rect 35836 139292 35900 139296
rect 35836 139236 35840 139292
rect 35840 139236 35896 139292
rect 35896 139236 35900 139292
rect 35836 139232 35900 139236
rect 66316 139292 66380 139296
rect 66316 139236 66320 139292
rect 66320 139236 66376 139292
rect 66376 139236 66380 139292
rect 66316 139232 66380 139236
rect 66396 139292 66460 139296
rect 66396 139236 66400 139292
rect 66400 139236 66456 139292
rect 66456 139236 66460 139292
rect 66396 139232 66460 139236
rect 66476 139292 66540 139296
rect 66476 139236 66480 139292
rect 66480 139236 66536 139292
rect 66536 139236 66540 139292
rect 66476 139232 66540 139236
rect 66556 139292 66620 139296
rect 66556 139236 66560 139292
rect 66560 139236 66616 139292
rect 66616 139236 66620 139292
rect 66556 139232 66620 139236
rect 97036 139292 97100 139296
rect 97036 139236 97040 139292
rect 97040 139236 97096 139292
rect 97096 139236 97100 139292
rect 97036 139232 97100 139236
rect 97116 139292 97180 139296
rect 97116 139236 97120 139292
rect 97120 139236 97176 139292
rect 97176 139236 97180 139292
rect 97116 139232 97180 139236
rect 97196 139292 97260 139296
rect 97196 139236 97200 139292
rect 97200 139236 97256 139292
rect 97256 139236 97260 139292
rect 97196 139232 97260 139236
rect 97276 139292 97340 139296
rect 97276 139236 97280 139292
rect 97280 139236 97336 139292
rect 97336 139236 97340 139292
rect 97276 139232 97340 139236
rect 4216 138748 4280 138752
rect 4216 138692 4220 138748
rect 4220 138692 4276 138748
rect 4276 138692 4280 138748
rect 4216 138688 4280 138692
rect 4296 138748 4360 138752
rect 4296 138692 4300 138748
rect 4300 138692 4356 138748
rect 4356 138692 4360 138748
rect 4296 138688 4360 138692
rect 4376 138748 4440 138752
rect 4376 138692 4380 138748
rect 4380 138692 4436 138748
rect 4436 138692 4440 138748
rect 4376 138688 4440 138692
rect 4456 138748 4520 138752
rect 4456 138692 4460 138748
rect 4460 138692 4516 138748
rect 4516 138692 4520 138748
rect 4456 138688 4520 138692
rect 34936 138748 35000 138752
rect 34936 138692 34940 138748
rect 34940 138692 34996 138748
rect 34996 138692 35000 138748
rect 34936 138688 35000 138692
rect 35016 138748 35080 138752
rect 35016 138692 35020 138748
rect 35020 138692 35076 138748
rect 35076 138692 35080 138748
rect 35016 138688 35080 138692
rect 35096 138748 35160 138752
rect 35096 138692 35100 138748
rect 35100 138692 35156 138748
rect 35156 138692 35160 138748
rect 35096 138688 35160 138692
rect 35176 138748 35240 138752
rect 35176 138692 35180 138748
rect 35180 138692 35236 138748
rect 35236 138692 35240 138748
rect 35176 138688 35240 138692
rect 65656 138748 65720 138752
rect 65656 138692 65660 138748
rect 65660 138692 65716 138748
rect 65716 138692 65720 138748
rect 65656 138688 65720 138692
rect 65736 138748 65800 138752
rect 65736 138692 65740 138748
rect 65740 138692 65796 138748
rect 65796 138692 65800 138748
rect 65736 138688 65800 138692
rect 65816 138748 65880 138752
rect 65816 138692 65820 138748
rect 65820 138692 65876 138748
rect 65876 138692 65880 138748
rect 65816 138688 65880 138692
rect 65896 138748 65960 138752
rect 65896 138692 65900 138748
rect 65900 138692 65956 138748
rect 65956 138692 65960 138748
rect 65896 138688 65960 138692
rect 96376 138748 96440 138752
rect 96376 138692 96380 138748
rect 96380 138692 96436 138748
rect 96436 138692 96440 138748
rect 96376 138688 96440 138692
rect 96456 138748 96520 138752
rect 96456 138692 96460 138748
rect 96460 138692 96516 138748
rect 96516 138692 96520 138748
rect 96456 138688 96520 138692
rect 96536 138748 96600 138752
rect 96536 138692 96540 138748
rect 96540 138692 96596 138748
rect 96596 138692 96600 138748
rect 96536 138688 96600 138692
rect 96616 138748 96680 138752
rect 96616 138692 96620 138748
rect 96620 138692 96676 138748
rect 96676 138692 96680 138748
rect 96616 138688 96680 138692
rect 4876 138204 4940 138208
rect 4876 138148 4880 138204
rect 4880 138148 4936 138204
rect 4936 138148 4940 138204
rect 4876 138144 4940 138148
rect 4956 138204 5020 138208
rect 4956 138148 4960 138204
rect 4960 138148 5016 138204
rect 5016 138148 5020 138204
rect 4956 138144 5020 138148
rect 5036 138204 5100 138208
rect 5036 138148 5040 138204
rect 5040 138148 5096 138204
rect 5096 138148 5100 138204
rect 5036 138144 5100 138148
rect 5116 138204 5180 138208
rect 5116 138148 5120 138204
rect 5120 138148 5176 138204
rect 5176 138148 5180 138204
rect 5116 138144 5180 138148
rect 35596 138204 35660 138208
rect 35596 138148 35600 138204
rect 35600 138148 35656 138204
rect 35656 138148 35660 138204
rect 35596 138144 35660 138148
rect 35676 138204 35740 138208
rect 35676 138148 35680 138204
rect 35680 138148 35736 138204
rect 35736 138148 35740 138204
rect 35676 138144 35740 138148
rect 35756 138204 35820 138208
rect 35756 138148 35760 138204
rect 35760 138148 35816 138204
rect 35816 138148 35820 138204
rect 35756 138144 35820 138148
rect 35836 138204 35900 138208
rect 35836 138148 35840 138204
rect 35840 138148 35896 138204
rect 35896 138148 35900 138204
rect 35836 138144 35900 138148
rect 66316 138204 66380 138208
rect 66316 138148 66320 138204
rect 66320 138148 66376 138204
rect 66376 138148 66380 138204
rect 66316 138144 66380 138148
rect 66396 138204 66460 138208
rect 66396 138148 66400 138204
rect 66400 138148 66456 138204
rect 66456 138148 66460 138204
rect 66396 138144 66460 138148
rect 66476 138204 66540 138208
rect 66476 138148 66480 138204
rect 66480 138148 66536 138204
rect 66536 138148 66540 138204
rect 66476 138144 66540 138148
rect 66556 138204 66620 138208
rect 66556 138148 66560 138204
rect 66560 138148 66616 138204
rect 66616 138148 66620 138204
rect 66556 138144 66620 138148
rect 97036 138204 97100 138208
rect 97036 138148 97040 138204
rect 97040 138148 97096 138204
rect 97096 138148 97100 138204
rect 97036 138144 97100 138148
rect 97116 138204 97180 138208
rect 97116 138148 97120 138204
rect 97120 138148 97176 138204
rect 97176 138148 97180 138204
rect 97116 138144 97180 138148
rect 97196 138204 97260 138208
rect 97196 138148 97200 138204
rect 97200 138148 97256 138204
rect 97256 138148 97260 138204
rect 97196 138144 97260 138148
rect 97276 138204 97340 138208
rect 97276 138148 97280 138204
rect 97280 138148 97336 138204
rect 97336 138148 97340 138204
rect 97276 138144 97340 138148
rect 4216 137660 4280 137664
rect 4216 137604 4220 137660
rect 4220 137604 4276 137660
rect 4276 137604 4280 137660
rect 4216 137600 4280 137604
rect 4296 137660 4360 137664
rect 4296 137604 4300 137660
rect 4300 137604 4356 137660
rect 4356 137604 4360 137660
rect 4296 137600 4360 137604
rect 4376 137660 4440 137664
rect 4376 137604 4380 137660
rect 4380 137604 4436 137660
rect 4436 137604 4440 137660
rect 4376 137600 4440 137604
rect 4456 137660 4520 137664
rect 4456 137604 4460 137660
rect 4460 137604 4516 137660
rect 4516 137604 4520 137660
rect 4456 137600 4520 137604
rect 34936 137660 35000 137664
rect 34936 137604 34940 137660
rect 34940 137604 34996 137660
rect 34996 137604 35000 137660
rect 34936 137600 35000 137604
rect 35016 137660 35080 137664
rect 35016 137604 35020 137660
rect 35020 137604 35076 137660
rect 35076 137604 35080 137660
rect 35016 137600 35080 137604
rect 35096 137660 35160 137664
rect 35096 137604 35100 137660
rect 35100 137604 35156 137660
rect 35156 137604 35160 137660
rect 35096 137600 35160 137604
rect 35176 137660 35240 137664
rect 35176 137604 35180 137660
rect 35180 137604 35236 137660
rect 35236 137604 35240 137660
rect 35176 137600 35240 137604
rect 65656 137660 65720 137664
rect 65656 137604 65660 137660
rect 65660 137604 65716 137660
rect 65716 137604 65720 137660
rect 65656 137600 65720 137604
rect 65736 137660 65800 137664
rect 65736 137604 65740 137660
rect 65740 137604 65796 137660
rect 65796 137604 65800 137660
rect 65736 137600 65800 137604
rect 65816 137660 65880 137664
rect 65816 137604 65820 137660
rect 65820 137604 65876 137660
rect 65876 137604 65880 137660
rect 65816 137600 65880 137604
rect 65896 137660 65960 137664
rect 65896 137604 65900 137660
rect 65900 137604 65956 137660
rect 65956 137604 65960 137660
rect 65896 137600 65960 137604
rect 96376 137660 96440 137664
rect 96376 137604 96380 137660
rect 96380 137604 96436 137660
rect 96436 137604 96440 137660
rect 96376 137600 96440 137604
rect 96456 137660 96520 137664
rect 96456 137604 96460 137660
rect 96460 137604 96516 137660
rect 96516 137604 96520 137660
rect 96456 137600 96520 137604
rect 96536 137660 96600 137664
rect 96536 137604 96540 137660
rect 96540 137604 96596 137660
rect 96596 137604 96600 137660
rect 96536 137600 96600 137604
rect 96616 137660 96680 137664
rect 96616 137604 96620 137660
rect 96620 137604 96676 137660
rect 96676 137604 96680 137660
rect 96616 137600 96680 137604
rect 4876 137116 4940 137120
rect 4876 137060 4880 137116
rect 4880 137060 4936 137116
rect 4936 137060 4940 137116
rect 4876 137056 4940 137060
rect 4956 137116 5020 137120
rect 4956 137060 4960 137116
rect 4960 137060 5016 137116
rect 5016 137060 5020 137116
rect 4956 137056 5020 137060
rect 5036 137116 5100 137120
rect 5036 137060 5040 137116
rect 5040 137060 5096 137116
rect 5096 137060 5100 137116
rect 5036 137056 5100 137060
rect 5116 137116 5180 137120
rect 5116 137060 5120 137116
rect 5120 137060 5176 137116
rect 5176 137060 5180 137116
rect 5116 137056 5180 137060
rect 35596 137116 35660 137120
rect 35596 137060 35600 137116
rect 35600 137060 35656 137116
rect 35656 137060 35660 137116
rect 35596 137056 35660 137060
rect 35676 137116 35740 137120
rect 35676 137060 35680 137116
rect 35680 137060 35736 137116
rect 35736 137060 35740 137116
rect 35676 137056 35740 137060
rect 35756 137116 35820 137120
rect 35756 137060 35760 137116
rect 35760 137060 35816 137116
rect 35816 137060 35820 137116
rect 35756 137056 35820 137060
rect 35836 137116 35900 137120
rect 35836 137060 35840 137116
rect 35840 137060 35896 137116
rect 35896 137060 35900 137116
rect 35836 137056 35900 137060
rect 66316 137116 66380 137120
rect 66316 137060 66320 137116
rect 66320 137060 66376 137116
rect 66376 137060 66380 137116
rect 66316 137056 66380 137060
rect 66396 137116 66460 137120
rect 66396 137060 66400 137116
rect 66400 137060 66456 137116
rect 66456 137060 66460 137116
rect 66396 137056 66460 137060
rect 66476 137116 66540 137120
rect 66476 137060 66480 137116
rect 66480 137060 66536 137116
rect 66536 137060 66540 137116
rect 66476 137056 66540 137060
rect 66556 137116 66620 137120
rect 66556 137060 66560 137116
rect 66560 137060 66616 137116
rect 66616 137060 66620 137116
rect 66556 137056 66620 137060
rect 97036 137116 97100 137120
rect 97036 137060 97040 137116
rect 97040 137060 97096 137116
rect 97096 137060 97100 137116
rect 97036 137056 97100 137060
rect 97116 137116 97180 137120
rect 97116 137060 97120 137116
rect 97120 137060 97176 137116
rect 97176 137060 97180 137116
rect 97116 137056 97180 137060
rect 97196 137116 97260 137120
rect 97196 137060 97200 137116
rect 97200 137060 97256 137116
rect 97256 137060 97260 137116
rect 97196 137056 97260 137060
rect 97276 137116 97340 137120
rect 97276 137060 97280 137116
rect 97280 137060 97336 137116
rect 97336 137060 97340 137116
rect 97276 137056 97340 137060
rect 4216 136572 4280 136576
rect 4216 136516 4220 136572
rect 4220 136516 4276 136572
rect 4276 136516 4280 136572
rect 4216 136512 4280 136516
rect 4296 136572 4360 136576
rect 4296 136516 4300 136572
rect 4300 136516 4356 136572
rect 4356 136516 4360 136572
rect 4296 136512 4360 136516
rect 4376 136572 4440 136576
rect 4376 136516 4380 136572
rect 4380 136516 4436 136572
rect 4436 136516 4440 136572
rect 4376 136512 4440 136516
rect 4456 136572 4520 136576
rect 4456 136516 4460 136572
rect 4460 136516 4516 136572
rect 4516 136516 4520 136572
rect 4456 136512 4520 136516
rect 34936 136572 35000 136576
rect 34936 136516 34940 136572
rect 34940 136516 34996 136572
rect 34996 136516 35000 136572
rect 34936 136512 35000 136516
rect 35016 136572 35080 136576
rect 35016 136516 35020 136572
rect 35020 136516 35076 136572
rect 35076 136516 35080 136572
rect 35016 136512 35080 136516
rect 35096 136572 35160 136576
rect 35096 136516 35100 136572
rect 35100 136516 35156 136572
rect 35156 136516 35160 136572
rect 35096 136512 35160 136516
rect 35176 136572 35240 136576
rect 35176 136516 35180 136572
rect 35180 136516 35236 136572
rect 35236 136516 35240 136572
rect 35176 136512 35240 136516
rect 65656 136572 65720 136576
rect 65656 136516 65660 136572
rect 65660 136516 65716 136572
rect 65716 136516 65720 136572
rect 65656 136512 65720 136516
rect 65736 136572 65800 136576
rect 65736 136516 65740 136572
rect 65740 136516 65796 136572
rect 65796 136516 65800 136572
rect 65736 136512 65800 136516
rect 65816 136572 65880 136576
rect 65816 136516 65820 136572
rect 65820 136516 65876 136572
rect 65876 136516 65880 136572
rect 65816 136512 65880 136516
rect 65896 136572 65960 136576
rect 65896 136516 65900 136572
rect 65900 136516 65956 136572
rect 65956 136516 65960 136572
rect 65896 136512 65960 136516
rect 96376 136572 96440 136576
rect 96376 136516 96380 136572
rect 96380 136516 96436 136572
rect 96436 136516 96440 136572
rect 96376 136512 96440 136516
rect 96456 136572 96520 136576
rect 96456 136516 96460 136572
rect 96460 136516 96516 136572
rect 96516 136516 96520 136572
rect 96456 136512 96520 136516
rect 96536 136572 96600 136576
rect 96536 136516 96540 136572
rect 96540 136516 96596 136572
rect 96596 136516 96600 136572
rect 96536 136512 96600 136516
rect 96616 136572 96680 136576
rect 96616 136516 96620 136572
rect 96620 136516 96676 136572
rect 96676 136516 96680 136572
rect 96616 136512 96680 136516
rect 105924 136572 105988 136576
rect 105924 136516 105928 136572
rect 105928 136516 105984 136572
rect 105984 136516 105988 136572
rect 105924 136512 105988 136516
rect 106004 136572 106068 136576
rect 106004 136516 106008 136572
rect 106008 136516 106064 136572
rect 106064 136516 106068 136572
rect 106004 136512 106068 136516
rect 106084 136572 106148 136576
rect 106084 136516 106088 136572
rect 106088 136516 106144 136572
rect 106144 136516 106148 136572
rect 106084 136512 106148 136516
rect 106164 136572 106228 136576
rect 106164 136516 106168 136572
rect 106168 136516 106224 136572
rect 106224 136516 106228 136572
rect 106164 136512 106228 136516
rect 4876 136028 4940 136032
rect 4876 135972 4880 136028
rect 4880 135972 4936 136028
rect 4936 135972 4940 136028
rect 4876 135968 4940 135972
rect 4956 136028 5020 136032
rect 4956 135972 4960 136028
rect 4960 135972 5016 136028
rect 5016 135972 5020 136028
rect 4956 135968 5020 135972
rect 5036 136028 5100 136032
rect 5036 135972 5040 136028
rect 5040 135972 5096 136028
rect 5096 135972 5100 136028
rect 5036 135968 5100 135972
rect 5116 136028 5180 136032
rect 5116 135972 5120 136028
rect 5120 135972 5176 136028
rect 5176 135972 5180 136028
rect 5116 135968 5180 135972
rect 35596 136028 35660 136032
rect 35596 135972 35600 136028
rect 35600 135972 35656 136028
rect 35656 135972 35660 136028
rect 35596 135968 35660 135972
rect 35676 136028 35740 136032
rect 35676 135972 35680 136028
rect 35680 135972 35736 136028
rect 35736 135972 35740 136028
rect 35676 135968 35740 135972
rect 35756 136028 35820 136032
rect 35756 135972 35760 136028
rect 35760 135972 35816 136028
rect 35816 135972 35820 136028
rect 35756 135968 35820 135972
rect 35836 136028 35900 136032
rect 35836 135972 35840 136028
rect 35840 135972 35896 136028
rect 35896 135972 35900 136028
rect 35836 135968 35900 135972
rect 66316 136028 66380 136032
rect 66316 135972 66320 136028
rect 66320 135972 66376 136028
rect 66376 135972 66380 136028
rect 66316 135968 66380 135972
rect 66396 136028 66460 136032
rect 66396 135972 66400 136028
rect 66400 135972 66456 136028
rect 66456 135972 66460 136028
rect 66396 135968 66460 135972
rect 66476 136028 66540 136032
rect 66476 135972 66480 136028
rect 66480 135972 66536 136028
rect 66536 135972 66540 136028
rect 66476 135968 66540 135972
rect 66556 136028 66620 136032
rect 66556 135972 66560 136028
rect 66560 135972 66616 136028
rect 66616 135972 66620 136028
rect 66556 135968 66620 135972
rect 97036 136028 97100 136032
rect 97036 135972 97040 136028
rect 97040 135972 97096 136028
rect 97096 135972 97100 136028
rect 97036 135968 97100 135972
rect 97116 136028 97180 136032
rect 97116 135972 97120 136028
rect 97120 135972 97176 136028
rect 97176 135972 97180 136028
rect 97116 135968 97180 135972
rect 97196 136028 97260 136032
rect 97196 135972 97200 136028
rect 97200 135972 97256 136028
rect 97256 135972 97260 136028
rect 97196 135968 97260 135972
rect 97276 136028 97340 136032
rect 97276 135972 97280 136028
rect 97280 135972 97336 136028
rect 97336 135972 97340 136028
rect 97276 135968 97340 135972
rect 106660 136028 106724 136032
rect 106660 135972 106664 136028
rect 106664 135972 106720 136028
rect 106720 135972 106724 136028
rect 106660 135968 106724 135972
rect 106740 136028 106804 136032
rect 106740 135972 106744 136028
rect 106744 135972 106800 136028
rect 106800 135972 106804 136028
rect 106740 135968 106804 135972
rect 106820 136028 106884 136032
rect 106820 135972 106824 136028
rect 106824 135972 106880 136028
rect 106880 135972 106884 136028
rect 106820 135968 106884 135972
rect 106900 136028 106964 136032
rect 106900 135972 106904 136028
rect 106904 135972 106960 136028
rect 106960 135972 106964 136028
rect 106900 135968 106964 135972
rect 95924 135688 95988 135692
rect 95924 135632 95974 135688
rect 95974 135632 95988 135688
rect 95924 135628 95988 135632
rect 4216 135484 4280 135488
rect 4216 135428 4220 135484
rect 4220 135428 4276 135484
rect 4276 135428 4280 135484
rect 4216 135424 4280 135428
rect 4296 135484 4360 135488
rect 4296 135428 4300 135484
rect 4300 135428 4356 135484
rect 4356 135428 4360 135484
rect 4296 135424 4360 135428
rect 4376 135484 4440 135488
rect 4376 135428 4380 135484
rect 4380 135428 4436 135484
rect 4436 135428 4440 135484
rect 4376 135424 4440 135428
rect 4456 135484 4520 135488
rect 4456 135428 4460 135484
rect 4460 135428 4516 135484
rect 4516 135428 4520 135484
rect 4456 135424 4520 135428
rect 105924 135484 105988 135488
rect 105924 135428 105928 135484
rect 105928 135428 105984 135484
rect 105984 135428 105988 135484
rect 105924 135424 105988 135428
rect 106004 135484 106068 135488
rect 106004 135428 106008 135484
rect 106008 135428 106064 135484
rect 106064 135428 106068 135484
rect 106004 135424 106068 135428
rect 106084 135484 106148 135488
rect 106084 135428 106088 135484
rect 106088 135428 106144 135484
rect 106144 135428 106148 135484
rect 106084 135424 106148 135428
rect 106164 135484 106228 135488
rect 106164 135428 106168 135484
rect 106168 135428 106224 135484
rect 106224 135428 106228 135484
rect 106164 135424 106228 135428
rect 58572 135220 58636 135284
rect 61148 135220 61212 135284
rect 71084 135220 71148 135284
rect 63540 135144 63604 135148
rect 63540 135088 63590 135144
rect 63590 135088 63604 135144
rect 63540 135084 63604 135088
rect 4876 134940 4940 134944
rect 4876 134884 4880 134940
rect 4880 134884 4936 134940
rect 4936 134884 4940 134940
rect 4876 134880 4940 134884
rect 4956 134940 5020 134944
rect 4956 134884 4960 134940
rect 4960 134884 5016 134940
rect 5016 134884 5020 134940
rect 4956 134880 5020 134884
rect 5036 134940 5100 134944
rect 5036 134884 5040 134940
rect 5040 134884 5096 134940
rect 5096 134884 5100 134940
rect 5036 134880 5100 134884
rect 5116 134940 5180 134944
rect 5116 134884 5120 134940
rect 5120 134884 5176 134940
rect 5176 134884 5180 134940
rect 5116 134880 5180 134884
rect 106660 134940 106724 134944
rect 106660 134884 106664 134940
rect 106664 134884 106720 134940
rect 106720 134884 106724 134940
rect 106660 134880 106724 134884
rect 106740 134940 106804 134944
rect 106740 134884 106744 134940
rect 106744 134884 106800 134940
rect 106800 134884 106804 134940
rect 106740 134880 106804 134884
rect 106820 134940 106884 134944
rect 106820 134884 106824 134940
rect 106824 134884 106880 134940
rect 106880 134884 106884 134940
rect 106820 134880 106884 134884
rect 106900 134940 106964 134944
rect 106900 134884 106904 134940
rect 106904 134884 106960 134940
rect 106960 134884 106964 134940
rect 106900 134880 106964 134884
rect 73476 134404 73540 134468
rect 4216 134396 4280 134400
rect 4216 134340 4220 134396
rect 4220 134340 4276 134396
rect 4276 134340 4280 134396
rect 4216 134336 4280 134340
rect 4296 134396 4360 134400
rect 4296 134340 4300 134396
rect 4300 134340 4356 134396
rect 4356 134340 4360 134396
rect 4296 134336 4360 134340
rect 4376 134396 4440 134400
rect 4376 134340 4380 134396
rect 4380 134340 4436 134396
rect 4436 134340 4440 134396
rect 4376 134336 4440 134340
rect 4456 134396 4520 134400
rect 4456 134340 4460 134396
rect 4460 134340 4516 134396
rect 4516 134340 4520 134396
rect 4456 134336 4520 134340
rect 105924 134396 105988 134400
rect 105924 134340 105928 134396
rect 105928 134340 105984 134396
rect 105984 134340 105988 134396
rect 105924 134336 105988 134340
rect 106004 134396 106068 134400
rect 106004 134340 106008 134396
rect 106008 134340 106064 134396
rect 106064 134340 106068 134396
rect 106004 134336 106068 134340
rect 106084 134396 106148 134400
rect 106084 134340 106088 134396
rect 106088 134340 106144 134396
rect 106144 134340 106148 134396
rect 106084 134336 106148 134340
rect 106164 134396 106228 134400
rect 106164 134340 106168 134396
rect 106168 134340 106224 134396
rect 106224 134340 106228 134396
rect 106164 134336 106228 134340
rect 41067 134132 41131 134196
rect 43563 134132 43627 134196
rect 53547 134132 53611 134196
rect 56043 134132 56107 134196
rect 66027 134132 66091 134196
rect 36075 133920 36139 133924
rect 36075 133864 36082 133920
rect 36082 133864 36138 133920
rect 36138 133864 36139 133920
rect 36075 133860 36139 133864
rect 38571 133920 38635 133924
rect 38571 133864 38622 133920
rect 38622 133864 38635 133920
rect 38571 133860 38635 133864
rect 46060 133920 46124 133924
rect 46060 133864 46110 133920
rect 46110 133864 46124 133920
rect 46060 133860 46124 133864
rect 48544 133920 48608 133924
rect 48544 133864 48558 133920
rect 48558 133864 48608 133920
rect 48544 133860 48608 133864
rect 51051 133920 51115 133924
rect 51051 133864 51078 133920
rect 51078 133864 51115 133920
rect 51051 133860 51115 133864
rect 68523 133920 68587 133924
rect 68523 133864 68558 133920
rect 68558 133864 68587 133920
rect 68523 133860 68587 133864
rect 86142 133860 86206 133924
rect 87310 133920 87374 133924
rect 87310 133864 87326 133920
rect 87326 133864 87374 133920
rect 87310 133860 87374 133864
rect 4876 133852 4940 133856
rect 4876 133796 4880 133852
rect 4880 133796 4936 133852
rect 4936 133796 4940 133852
rect 4876 133792 4940 133796
rect 4956 133852 5020 133856
rect 4956 133796 4960 133852
rect 4960 133796 5016 133852
rect 5016 133796 5020 133852
rect 4956 133792 5020 133796
rect 5036 133852 5100 133856
rect 5036 133796 5040 133852
rect 5040 133796 5096 133852
rect 5096 133796 5100 133852
rect 5036 133792 5100 133796
rect 5116 133852 5180 133856
rect 5116 133796 5120 133852
rect 5120 133796 5176 133852
rect 5176 133796 5180 133852
rect 5116 133792 5180 133796
rect 106660 133852 106724 133856
rect 106660 133796 106664 133852
rect 106664 133796 106720 133852
rect 106720 133796 106724 133852
rect 106660 133792 106724 133796
rect 106740 133852 106804 133856
rect 106740 133796 106744 133852
rect 106744 133796 106800 133852
rect 106800 133796 106804 133852
rect 106740 133792 106804 133796
rect 106820 133852 106884 133856
rect 106820 133796 106824 133852
rect 106824 133796 106880 133852
rect 106880 133796 106884 133852
rect 106820 133792 106884 133796
rect 106900 133852 106964 133856
rect 106900 133796 106904 133852
rect 106904 133796 106960 133852
rect 106960 133796 106964 133852
rect 106900 133792 106964 133796
rect 4216 133308 4280 133312
rect 4216 133252 4220 133308
rect 4220 133252 4276 133308
rect 4276 133252 4280 133308
rect 4216 133248 4280 133252
rect 4296 133308 4360 133312
rect 4296 133252 4300 133308
rect 4300 133252 4356 133308
rect 4356 133252 4360 133308
rect 4296 133248 4360 133252
rect 4376 133308 4440 133312
rect 4376 133252 4380 133308
rect 4380 133252 4436 133308
rect 4436 133252 4440 133308
rect 4376 133248 4440 133252
rect 4456 133308 4520 133312
rect 4456 133252 4460 133308
rect 4460 133252 4516 133308
rect 4516 133252 4520 133308
rect 4456 133248 4520 133252
rect 105924 133308 105988 133312
rect 105924 133252 105928 133308
rect 105928 133252 105984 133308
rect 105984 133252 105988 133308
rect 105924 133248 105988 133252
rect 106004 133308 106068 133312
rect 106004 133252 106008 133308
rect 106008 133252 106064 133308
rect 106064 133252 106068 133308
rect 106004 133248 106068 133252
rect 106084 133308 106148 133312
rect 106084 133252 106088 133308
rect 106088 133252 106144 133308
rect 106144 133252 106148 133308
rect 106084 133248 106148 133252
rect 106164 133308 106228 133312
rect 106164 133252 106168 133308
rect 106168 133252 106224 133308
rect 106224 133252 106228 133308
rect 106164 133248 106228 133252
rect 4876 132764 4940 132768
rect 4876 132708 4880 132764
rect 4880 132708 4936 132764
rect 4936 132708 4940 132764
rect 4876 132704 4940 132708
rect 4956 132764 5020 132768
rect 4956 132708 4960 132764
rect 4960 132708 5016 132764
rect 5016 132708 5020 132764
rect 4956 132704 5020 132708
rect 5036 132764 5100 132768
rect 5036 132708 5040 132764
rect 5040 132708 5096 132764
rect 5096 132708 5100 132764
rect 5036 132704 5100 132708
rect 5116 132764 5180 132768
rect 5116 132708 5120 132764
rect 5120 132708 5176 132764
rect 5176 132708 5180 132764
rect 5116 132704 5180 132708
rect 106660 132764 106724 132768
rect 106660 132708 106664 132764
rect 106664 132708 106720 132764
rect 106720 132708 106724 132764
rect 106660 132704 106724 132708
rect 106740 132764 106804 132768
rect 106740 132708 106744 132764
rect 106744 132708 106800 132764
rect 106800 132708 106804 132764
rect 106740 132704 106804 132708
rect 106820 132764 106884 132768
rect 106820 132708 106824 132764
rect 106824 132708 106880 132764
rect 106880 132708 106884 132764
rect 106820 132704 106884 132708
rect 106900 132764 106964 132768
rect 106900 132708 106904 132764
rect 106904 132708 106960 132764
rect 106960 132708 106964 132764
rect 106900 132704 106964 132708
rect 4216 132220 4280 132224
rect 4216 132164 4220 132220
rect 4220 132164 4276 132220
rect 4276 132164 4280 132220
rect 4216 132160 4280 132164
rect 4296 132220 4360 132224
rect 4296 132164 4300 132220
rect 4300 132164 4356 132220
rect 4356 132164 4360 132220
rect 4296 132160 4360 132164
rect 4376 132220 4440 132224
rect 4376 132164 4380 132220
rect 4380 132164 4436 132220
rect 4436 132164 4440 132220
rect 4376 132160 4440 132164
rect 4456 132220 4520 132224
rect 4456 132164 4460 132220
rect 4460 132164 4516 132220
rect 4516 132164 4520 132220
rect 4456 132160 4520 132164
rect 105924 132220 105988 132224
rect 105924 132164 105928 132220
rect 105928 132164 105984 132220
rect 105984 132164 105988 132220
rect 105924 132160 105988 132164
rect 106004 132220 106068 132224
rect 106004 132164 106008 132220
rect 106008 132164 106064 132220
rect 106064 132164 106068 132220
rect 106004 132160 106068 132164
rect 106084 132220 106148 132224
rect 106084 132164 106088 132220
rect 106088 132164 106144 132220
rect 106144 132164 106148 132220
rect 106084 132160 106148 132164
rect 106164 132220 106228 132224
rect 106164 132164 106168 132220
rect 106168 132164 106224 132220
rect 106224 132164 106228 132220
rect 106164 132160 106228 132164
rect 4876 131676 4940 131680
rect 4876 131620 4880 131676
rect 4880 131620 4936 131676
rect 4936 131620 4940 131676
rect 4876 131616 4940 131620
rect 4956 131676 5020 131680
rect 4956 131620 4960 131676
rect 4960 131620 5016 131676
rect 5016 131620 5020 131676
rect 4956 131616 5020 131620
rect 5036 131676 5100 131680
rect 5036 131620 5040 131676
rect 5040 131620 5096 131676
rect 5096 131620 5100 131676
rect 5036 131616 5100 131620
rect 5116 131676 5180 131680
rect 5116 131620 5120 131676
rect 5120 131620 5176 131676
rect 5176 131620 5180 131676
rect 5116 131616 5180 131620
rect 106660 131676 106724 131680
rect 106660 131620 106664 131676
rect 106664 131620 106720 131676
rect 106720 131620 106724 131676
rect 106660 131616 106724 131620
rect 106740 131676 106804 131680
rect 106740 131620 106744 131676
rect 106744 131620 106800 131676
rect 106800 131620 106804 131676
rect 106740 131616 106804 131620
rect 106820 131676 106884 131680
rect 106820 131620 106824 131676
rect 106824 131620 106880 131676
rect 106880 131620 106884 131676
rect 106820 131616 106884 131620
rect 106900 131676 106964 131680
rect 106900 131620 106904 131676
rect 106904 131620 106960 131676
rect 106960 131620 106964 131676
rect 106900 131616 106964 131620
rect 4216 131132 4280 131136
rect 4216 131076 4220 131132
rect 4220 131076 4276 131132
rect 4276 131076 4280 131132
rect 4216 131072 4280 131076
rect 4296 131132 4360 131136
rect 4296 131076 4300 131132
rect 4300 131076 4356 131132
rect 4356 131076 4360 131132
rect 4296 131072 4360 131076
rect 4376 131132 4440 131136
rect 4376 131076 4380 131132
rect 4380 131076 4436 131132
rect 4436 131076 4440 131132
rect 4376 131072 4440 131076
rect 4456 131132 4520 131136
rect 4456 131076 4460 131132
rect 4460 131076 4516 131132
rect 4516 131076 4520 131132
rect 4456 131072 4520 131076
rect 105924 131132 105988 131136
rect 105924 131076 105928 131132
rect 105928 131076 105984 131132
rect 105984 131076 105988 131132
rect 105924 131072 105988 131076
rect 106004 131132 106068 131136
rect 106004 131076 106008 131132
rect 106008 131076 106064 131132
rect 106064 131076 106068 131132
rect 106004 131072 106068 131076
rect 106084 131132 106148 131136
rect 106084 131076 106088 131132
rect 106088 131076 106144 131132
rect 106144 131076 106148 131132
rect 106084 131072 106148 131076
rect 106164 131132 106228 131136
rect 106164 131076 106168 131132
rect 106168 131076 106224 131132
rect 106224 131076 106228 131132
rect 106164 131072 106228 131076
rect 4876 130588 4940 130592
rect 4876 130532 4880 130588
rect 4880 130532 4936 130588
rect 4936 130532 4940 130588
rect 4876 130528 4940 130532
rect 4956 130588 5020 130592
rect 4956 130532 4960 130588
rect 4960 130532 5016 130588
rect 5016 130532 5020 130588
rect 4956 130528 5020 130532
rect 5036 130588 5100 130592
rect 5036 130532 5040 130588
rect 5040 130532 5096 130588
rect 5096 130532 5100 130588
rect 5036 130528 5100 130532
rect 5116 130588 5180 130592
rect 5116 130532 5120 130588
rect 5120 130532 5176 130588
rect 5176 130532 5180 130588
rect 5116 130528 5180 130532
rect 106660 130588 106724 130592
rect 106660 130532 106664 130588
rect 106664 130532 106720 130588
rect 106720 130532 106724 130588
rect 106660 130528 106724 130532
rect 106740 130588 106804 130592
rect 106740 130532 106744 130588
rect 106744 130532 106800 130588
rect 106800 130532 106804 130588
rect 106740 130528 106804 130532
rect 106820 130588 106884 130592
rect 106820 130532 106824 130588
rect 106824 130532 106880 130588
rect 106880 130532 106884 130588
rect 106820 130528 106884 130532
rect 106900 130588 106964 130592
rect 106900 130532 106904 130588
rect 106904 130532 106960 130588
rect 106960 130532 106964 130588
rect 106900 130528 106964 130532
rect 4216 130044 4280 130048
rect 4216 129988 4220 130044
rect 4220 129988 4276 130044
rect 4276 129988 4280 130044
rect 4216 129984 4280 129988
rect 4296 130044 4360 130048
rect 4296 129988 4300 130044
rect 4300 129988 4356 130044
rect 4356 129988 4360 130044
rect 4296 129984 4360 129988
rect 4376 130044 4440 130048
rect 4376 129988 4380 130044
rect 4380 129988 4436 130044
rect 4436 129988 4440 130044
rect 4376 129984 4440 129988
rect 4456 130044 4520 130048
rect 4456 129988 4460 130044
rect 4460 129988 4516 130044
rect 4516 129988 4520 130044
rect 4456 129984 4520 129988
rect 105924 130044 105988 130048
rect 105924 129988 105928 130044
rect 105928 129988 105984 130044
rect 105984 129988 105988 130044
rect 105924 129984 105988 129988
rect 106004 130044 106068 130048
rect 106004 129988 106008 130044
rect 106008 129988 106064 130044
rect 106064 129988 106068 130044
rect 106004 129984 106068 129988
rect 106084 130044 106148 130048
rect 106084 129988 106088 130044
rect 106088 129988 106144 130044
rect 106144 129988 106148 130044
rect 106084 129984 106148 129988
rect 106164 130044 106228 130048
rect 106164 129988 106168 130044
rect 106168 129988 106224 130044
rect 106224 129988 106228 130044
rect 106164 129984 106228 129988
rect 4876 129500 4940 129504
rect 4876 129444 4880 129500
rect 4880 129444 4936 129500
rect 4936 129444 4940 129500
rect 4876 129440 4940 129444
rect 4956 129500 5020 129504
rect 4956 129444 4960 129500
rect 4960 129444 5016 129500
rect 5016 129444 5020 129500
rect 4956 129440 5020 129444
rect 5036 129500 5100 129504
rect 5036 129444 5040 129500
rect 5040 129444 5096 129500
rect 5096 129444 5100 129500
rect 5036 129440 5100 129444
rect 5116 129500 5180 129504
rect 5116 129444 5120 129500
rect 5120 129444 5176 129500
rect 5176 129444 5180 129500
rect 5116 129440 5180 129444
rect 106660 129500 106724 129504
rect 106660 129444 106664 129500
rect 106664 129444 106720 129500
rect 106720 129444 106724 129500
rect 106660 129440 106724 129444
rect 106740 129500 106804 129504
rect 106740 129444 106744 129500
rect 106744 129444 106800 129500
rect 106800 129444 106804 129500
rect 106740 129440 106804 129444
rect 106820 129500 106884 129504
rect 106820 129444 106824 129500
rect 106824 129444 106880 129500
rect 106880 129444 106884 129500
rect 106820 129440 106884 129444
rect 106900 129500 106964 129504
rect 106900 129444 106904 129500
rect 106904 129444 106960 129500
rect 106960 129444 106964 129500
rect 106900 129440 106964 129444
rect 4216 128956 4280 128960
rect 4216 128900 4220 128956
rect 4220 128900 4276 128956
rect 4276 128900 4280 128956
rect 4216 128896 4280 128900
rect 4296 128956 4360 128960
rect 4296 128900 4300 128956
rect 4300 128900 4356 128956
rect 4356 128900 4360 128956
rect 4296 128896 4360 128900
rect 4376 128956 4440 128960
rect 4376 128900 4380 128956
rect 4380 128900 4436 128956
rect 4436 128900 4440 128956
rect 4376 128896 4440 128900
rect 4456 128956 4520 128960
rect 4456 128900 4460 128956
rect 4460 128900 4516 128956
rect 4516 128900 4520 128956
rect 4456 128896 4520 128900
rect 105924 128956 105988 128960
rect 105924 128900 105928 128956
rect 105928 128900 105984 128956
rect 105984 128900 105988 128956
rect 105924 128896 105988 128900
rect 106004 128956 106068 128960
rect 106004 128900 106008 128956
rect 106008 128900 106064 128956
rect 106064 128900 106068 128956
rect 106004 128896 106068 128900
rect 106084 128956 106148 128960
rect 106084 128900 106088 128956
rect 106088 128900 106144 128956
rect 106144 128900 106148 128956
rect 106084 128896 106148 128900
rect 106164 128956 106228 128960
rect 106164 128900 106168 128956
rect 106168 128900 106224 128956
rect 106224 128900 106228 128956
rect 106164 128896 106228 128900
rect 4876 128412 4940 128416
rect 4876 128356 4880 128412
rect 4880 128356 4936 128412
rect 4936 128356 4940 128412
rect 4876 128352 4940 128356
rect 4956 128412 5020 128416
rect 4956 128356 4960 128412
rect 4960 128356 5016 128412
rect 5016 128356 5020 128412
rect 4956 128352 5020 128356
rect 5036 128412 5100 128416
rect 5036 128356 5040 128412
rect 5040 128356 5096 128412
rect 5096 128356 5100 128412
rect 5036 128352 5100 128356
rect 5116 128412 5180 128416
rect 5116 128356 5120 128412
rect 5120 128356 5176 128412
rect 5176 128356 5180 128412
rect 5116 128352 5180 128356
rect 106660 128412 106724 128416
rect 106660 128356 106664 128412
rect 106664 128356 106720 128412
rect 106720 128356 106724 128412
rect 106660 128352 106724 128356
rect 106740 128412 106804 128416
rect 106740 128356 106744 128412
rect 106744 128356 106800 128412
rect 106800 128356 106804 128412
rect 106740 128352 106804 128356
rect 106820 128412 106884 128416
rect 106820 128356 106824 128412
rect 106824 128356 106880 128412
rect 106880 128356 106884 128412
rect 106820 128352 106884 128356
rect 106900 128412 106964 128416
rect 106900 128356 106904 128412
rect 106904 128356 106960 128412
rect 106960 128356 106964 128412
rect 106900 128352 106964 128356
rect 4216 127868 4280 127872
rect 4216 127812 4220 127868
rect 4220 127812 4276 127868
rect 4276 127812 4280 127868
rect 4216 127808 4280 127812
rect 4296 127868 4360 127872
rect 4296 127812 4300 127868
rect 4300 127812 4356 127868
rect 4356 127812 4360 127868
rect 4296 127808 4360 127812
rect 4376 127868 4440 127872
rect 4376 127812 4380 127868
rect 4380 127812 4436 127868
rect 4436 127812 4440 127868
rect 4376 127808 4440 127812
rect 4456 127868 4520 127872
rect 4456 127812 4460 127868
rect 4460 127812 4516 127868
rect 4516 127812 4520 127868
rect 4456 127808 4520 127812
rect 105924 127868 105988 127872
rect 105924 127812 105928 127868
rect 105928 127812 105984 127868
rect 105984 127812 105988 127868
rect 105924 127808 105988 127812
rect 106004 127868 106068 127872
rect 106004 127812 106008 127868
rect 106008 127812 106064 127868
rect 106064 127812 106068 127868
rect 106004 127808 106068 127812
rect 106084 127868 106148 127872
rect 106084 127812 106088 127868
rect 106088 127812 106144 127868
rect 106144 127812 106148 127868
rect 106084 127808 106148 127812
rect 106164 127868 106228 127872
rect 106164 127812 106168 127868
rect 106168 127812 106224 127868
rect 106224 127812 106228 127868
rect 106164 127808 106228 127812
rect 4876 127324 4940 127328
rect 4876 127268 4880 127324
rect 4880 127268 4936 127324
rect 4936 127268 4940 127324
rect 4876 127264 4940 127268
rect 4956 127324 5020 127328
rect 4956 127268 4960 127324
rect 4960 127268 5016 127324
rect 5016 127268 5020 127324
rect 4956 127264 5020 127268
rect 5036 127324 5100 127328
rect 5036 127268 5040 127324
rect 5040 127268 5096 127324
rect 5096 127268 5100 127324
rect 5036 127264 5100 127268
rect 5116 127324 5180 127328
rect 5116 127268 5120 127324
rect 5120 127268 5176 127324
rect 5176 127268 5180 127324
rect 5116 127264 5180 127268
rect 106660 127324 106724 127328
rect 106660 127268 106664 127324
rect 106664 127268 106720 127324
rect 106720 127268 106724 127324
rect 106660 127264 106724 127268
rect 106740 127324 106804 127328
rect 106740 127268 106744 127324
rect 106744 127268 106800 127324
rect 106800 127268 106804 127324
rect 106740 127264 106804 127268
rect 106820 127324 106884 127328
rect 106820 127268 106824 127324
rect 106824 127268 106880 127324
rect 106880 127268 106884 127324
rect 106820 127264 106884 127268
rect 106900 127324 106964 127328
rect 106900 127268 106904 127324
rect 106904 127268 106960 127324
rect 106960 127268 106964 127324
rect 106900 127264 106964 127268
rect 4216 126780 4280 126784
rect 4216 126724 4220 126780
rect 4220 126724 4276 126780
rect 4276 126724 4280 126780
rect 4216 126720 4280 126724
rect 4296 126780 4360 126784
rect 4296 126724 4300 126780
rect 4300 126724 4356 126780
rect 4356 126724 4360 126780
rect 4296 126720 4360 126724
rect 4376 126780 4440 126784
rect 4376 126724 4380 126780
rect 4380 126724 4436 126780
rect 4436 126724 4440 126780
rect 4376 126720 4440 126724
rect 4456 126780 4520 126784
rect 4456 126724 4460 126780
rect 4460 126724 4516 126780
rect 4516 126724 4520 126780
rect 4456 126720 4520 126724
rect 105924 126780 105988 126784
rect 105924 126724 105928 126780
rect 105928 126724 105984 126780
rect 105984 126724 105988 126780
rect 105924 126720 105988 126724
rect 106004 126780 106068 126784
rect 106004 126724 106008 126780
rect 106008 126724 106064 126780
rect 106064 126724 106068 126780
rect 106004 126720 106068 126724
rect 106084 126780 106148 126784
rect 106084 126724 106088 126780
rect 106088 126724 106144 126780
rect 106144 126724 106148 126780
rect 106084 126720 106148 126724
rect 106164 126780 106228 126784
rect 106164 126724 106168 126780
rect 106168 126724 106224 126780
rect 106224 126724 106228 126780
rect 106164 126720 106228 126724
rect 4876 126236 4940 126240
rect 4876 126180 4880 126236
rect 4880 126180 4936 126236
rect 4936 126180 4940 126236
rect 4876 126176 4940 126180
rect 4956 126236 5020 126240
rect 4956 126180 4960 126236
rect 4960 126180 5016 126236
rect 5016 126180 5020 126236
rect 4956 126176 5020 126180
rect 5036 126236 5100 126240
rect 5036 126180 5040 126236
rect 5040 126180 5096 126236
rect 5096 126180 5100 126236
rect 5036 126176 5100 126180
rect 5116 126236 5180 126240
rect 5116 126180 5120 126236
rect 5120 126180 5176 126236
rect 5176 126180 5180 126236
rect 5116 126176 5180 126180
rect 106660 126236 106724 126240
rect 106660 126180 106664 126236
rect 106664 126180 106720 126236
rect 106720 126180 106724 126236
rect 106660 126176 106724 126180
rect 106740 126236 106804 126240
rect 106740 126180 106744 126236
rect 106744 126180 106800 126236
rect 106800 126180 106804 126236
rect 106740 126176 106804 126180
rect 106820 126236 106884 126240
rect 106820 126180 106824 126236
rect 106824 126180 106880 126236
rect 106880 126180 106884 126236
rect 106820 126176 106884 126180
rect 106900 126236 106964 126240
rect 106900 126180 106904 126236
rect 106904 126180 106960 126236
rect 106960 126180 106964 126236
rect 106900 126176 106964 126180
rect 4216 125692 4280 125696
rect 4216 125636 4220 125692
rect 4220 125636 4276 125692
rect 4276 125636 4280 125692
rect 4216 125632 4280 125636
rect 4296 125692 4360 125696
rect 4296 125636 4300 125692
rect 4300 125636 4356 125692
rect 4356 125636 4360 125692
rect 4296 125632 4360 125636
rect 4376 125692 4440 125696
rect 4376 125636 4380 125692
rect 4380 125636 4436 125692
rect 4436 125636 4440 125692
rect 4376 125632 4440 125636
rect 4456 125692 4520 125696
rect 4456 125636 4460 125692
rect 4460 125636 4516 125692
rect 4516 125636 4520 125692
rect 4456 125632 4520 125636
rect 105924 125692 105988 125696
rect 105924 125636 105928 125692
rect 105928 125636 105984 125692
rect 105984 125636 105988 125692
rect 105924 125632 105988 125636
rect 106004 125692 106068 125696
rect 106004 125636 106008 125692
rect 106008 125636 106064 125692
rect 106064 125636 106068 125692
rect 106004 125632 106068 125636
rect 106084 125692 106148 125696
rect 106084 125636 106088 125692
rect 106088 125636 106144 125692
rect 106144 125636 106148 125692
rect 106084 125632 106148 125636
rect 106164 125692 106228 125696
rect 106164 125636 106168 125692
rect 106168 125636 106224 125692
rect 106224 125636 106228 125692
rect 106164 125632 106228 125636
rect 4876 125148 4940 125152
rect 4876 125092 4880 125148
rect 4880 125092 4936 125148
rect 4936 125092 4940 125148
rect 4876 125088 4940 125092
rect 4956 125148 5020 125152
rect 4956 125092 4960 125148
rect 4960 125092 5016 125148
rect 5016 125092 5020 125148
rect 4956 125088 5020 125092
rect 5036 125148 5100 125152
rect 5036 125092 5040 125148
rect 5040 125092 5096 125148
rect 5096 125092 5100 125148
rect 5036 125088 5100 125092
rect 5116 125148 5180 125152
rect 5116 125092 5120 125148
rect 5120 125092 5176 125148
rect 5176 125092 5180 125148
rect 5116 125088 5180 125092
rect 106660 125148 106724 125152
rect 106660 125092 106664 125148
rect 106664 125092 106720 125148
rect 106720 125092 106724 125148
rect 106660 125088 106724 125092
rect 106740 125148 106804 125152
rect 106740 125092 106744 125148
rect 106744 125092 106800 125148
rect 106800 125092 106804 125148
rect 106740 125088 106804 125092
rect 106820 125148 106884 125152
rect 106820 125092 106824 125148
rect 106824 125092 106880 125148
rect 106880 125092 106884 125148
rect 106820 125088 106884 125092
rect 106900 125148 106964 125152
rect 106900 125092 106904 125148
rect 106904 125092 106960 125148
rect 106960 125092 106964 125148
rect 106900 125088 106964 125092
rect 4216 124604 4280 124608
rect 4216 124548 4220 124604
rect 4220 124548 4276 124604
rect 4276 124548 4280 124604
rect 4216 124544 4280 124548
rect 4296 124604 4360 124608
rect 4296 124548 4300 124604
rect 4300 124548 4356 124604
rect 4356 124548 4360 124604
rect 4296 124544 4360 124548
rect 4376 124604 4440 124608
rect 4376 124548 4380 124604
rect 4380 124548 4436 124604
rect 4436 124548 4440 124604
rect 4376 124544 4440 124548
rect 4456 124604 4520 124608
rect 4456 124548 4460 124604
rect 4460 124548 4516 124604
rect 4516 124548 4520 124604
rect 4456 124544 4520 124548
rect 105924 124604 105988 124608
rect 105924 124548 105928 124604
rect 105928 124548 105984 124604
rect 105984 124548 105988 124604
rect 105924 124544 105988 124548
rect 106004 124604 106068 124608
rect 106004 124548 106008 124604
rect 106008 124548 106064 124604
rect 106064 124548 106068 124604
rect 106004 124544 106068 124548
rect 106084 124604 106148 124608
rect 106084 124548 106088 124604
rect 106088 124548 106144 124604
rect 106144 124548 106148 124604
rect 106084 124544 106148 124548
rect 106164 124604 106228 124608
rect 106164 124548 106168 124604
rect 106168 124548 106224 124604
rect 106224 124548 106228 124604
rect 106164 124544 106228 124548
rect 4876 124060 4940 124064
rect 4876 124004 4880 124060
rect 4880 124004 4936 124060
rect 4936 124004 4940 124060
rect 4876 124000 4940 124004
rect 4956 124060 5020 124064
rect 4956 124004 4960 124060
rect 4960 124004 5016 124060
rect 5016 124004 5020 124060
rect 4956 124000 5020 124004
rect 5036 124060 5100 124064
rect 5036 124004 5040 124060
rect 5040 124004 5096 124060
rect 5096 124004 5100 124060
rect 5036 124000 5100 124004
rect 5116 124060 5180 124064
rect 5116 124004 5120 124060
rect 5120 124004 5176 124060
rect 5176 124004 5180 124060
rect 5116 124000 5180 124004
rect 106660 124060 106724 124064
rect 106660 124004 106664 124060
rect 106664 124004 106720 124060
rect 106720 124004 106724 124060
rect 106660 124000 106724 124004
rect 106740 124060 106804 124064
rect 106740 124004 106744 124060
rect 106744 124004 106800 124060
rect 106800 124004 106804 124060
rect 106740 124000 106804 124004
rect 106820 124060 106884 124064
rect 106820 124004 106824 124060
rect 106824 124004 106880 124060
rect 106880 124004 106884 124060
rect 106820 124000 106884 124004
rect 106900 124060 106964 124064
rect 106900 124004 106904 124060
rect 106904 124004 106960 124060
rect 106960 124004 106964 124060
rect 106900 124000 106964 124004
rect 4216 123516 4280 123520
rect 4216 123460 4220 123516
rect 4220 123460 4276 123516
rect 4276 123460 4280 123516
rect 4216 123456 4280 123460
rect 4296 123516 4360 123520
rect 4296 123460 4300 123516
rect 4300 123460 4356 123516
rect 4356 123460 4360 123516
rect 4296 123456 4360 123460
rect 4376 123516 4440 123520
rect 4376 123460 4380 123516
rect 4380 123460 4436 123516
rect 4436 123460 4440 123516
rect 4376 123456 4440 123460
rect 4456 123516 4520 123520
rect 4456 123460 4460 123516
rect 4460 123460 4516 123516
rect 4516 123460 4520 123516
rect 4456 123456 4520 123460
rect 105924 123516 105988 123520
rect 105924 123460 105928 123516
rect 105928 123460 105984 123516
rect 105984 123460 105988 123516
rect 105924 123456 105988 123460
rect 106004 123516 106068 123520
rect 106004 123460 106008 123516
rect 106008 123460 106064 123516
rect 106064 123460 106068 123516
rect 106004 123456 106068 123460
rect 106084 123516 106148 123520
rect 106084 123460 106088 123516
rect 106088 123460 106144 123516
rect 106144 123460 106148 123516
rect 106084 123456 106148 123460
rect 106164 123516 106228 123520
rect 106164 123460 106168 123516
rect 106168 123460 106224 123516
rect 106224 123460 106228 123516
rect 106164 123456 106228 123460
rect 4876 122972 4940 122976
rect 4876 122916 4880 122972
rect 4880 122916 4936 122972
rect 4936 122916 4940 122972
rect 4876 122912 4940 122916
rect 4956 122972 5020 122976
rect 4956 122916 4960 122972
rect 4960 122916 5016 122972
rect 5016 122916 5020 122972
rect 4956 122912 5020 122916
rect 5036 122972 5100 122976
rect 5036 122916 5040 122972
rect 5040 122916 5096 122972
rect 5096 122916 5100 122972
rect 5036 122912 5100 122916
rect 5116 122972 5180 122976
rect 5116 122916 5120 122972
rect 5120 122916 5176 122972
rect 5176 122916 5180 122972
rect 5116 122912 5180 122916
rect 106660 122972 106724 122976
rect 106660 122916 106664 122972
rect 106664 122916 106720 122972
rect 106720 122916 106724 122972
rect 106660 122912 106724 122916
rect 106740 122972 106804 122976
rect 106740 122916 106744 122972
rect 106744 122916 106800 122972
rect 106800 122916 106804 122972
rect 106740 122912 106804 122916
rect 106820 122972 106884 122976
rect 106820 122916 106824 122972
rect 106824 122916 106880 122972
rect 106880 122916 106884 122972
rect 106820 122912 106884 122916
rect 106900 122972 106964 122976
rect 106900 122916 106904 122972
rect 106904 122916 106960 122972
rect 106960 122916 106964 122972
rect 106900 122912 106964 122916
rect 4216 122428 4280 122432
rect 4216 122372 4220 122428
rect 4220 122372 4276 122428
rect 4276 122372 4280 122428
rect 4216 122368 4280 122372
rect 4296 122428 4360 122432
rect 4296 122372 4300 122428
rect 4300 122372 4356 122428
rect 4356 122372 4360 122428
rect 4296 122368 4360 122372
rect 4376 122428 4440 122432
rect 4376 122372 4380 122428
rect 4380 122372 4436 122428
rect 4436 122372 4440 122428
rect 4376 122368 4440 122372
rect 4456 122428 4520 122432
rect 4456 122372 4460 122428
rect 4460 122372 4516 122428
rect 4516 122372 4520 122428
rect 4456 122368 4520 122372
rect 105924 122428 105988 122432
rect 105924 122372 105928 122428
rect 105928 122372 105984 122428
rect 105984 122372 105988 122428
rect 105924 122368 105988 122372
rect 106004 122428 106068 122432
rect 106004 122372 106008 122428
rect 106008 122372 106064 122428
rect 106064 122372 106068 122428
rect 106004 122368 106068 122372
rect 106084 122428 106148 122432
rect 106084 122372 106088 122428
rect 106088 122372 106144 122428
rect 106144 122372 106148 122428
rect 106084 122368 106148 122372
rect 106164 122428 106228 122432
rect 106164 122372 106168 122428
rect 106168 122372 106224 122428
rect 106224 122372 106228 122428
rect 106164 122368 106228 122372
rect 4876 121884 4940 121888
rect 4876 121828 4880 121884
rect 4880 121828 4936 121884
rect 4936 121828 4940 121884
rect 4876 121824 4940 121828
rect 4956 121884 5020 121888
rect 4956 121828 4960 121884
rect 4960 121828 5016 121884
rect 5016 121828 5020 121884
rect 4956 121824 5020 121828
rect 5036 121884 5100 121888
rect 5036 121828 5040 121884
rect 5040 121828 5096 121884
rect 5096 121828 5100 121884
rect 5036 121824 5100 121828
rect 5116 121884 5180 121888
rect 5116 121828 5120 121884
rect 5120 121828 5176 121884
rect 5176 121828 5180 121884
rect 5116 121824 5180 121828
rect 106660 121884 106724 121888
rect 106660 121828 106664 121884
rect 106664 121828 106720 121884
rect 106720 121828 106724 121884
rect 106660 121824 106724 121828
rect 106740 121884 106804 121888
rect 106740 121828 106744 121884
rect 106744 121828 106800 121884
rect 106800 121828 106804 121884
rect 106740 121824 106804 121828
rect 106820 121884 106884 121888
rect 106820 121828 106824 121884
rect 106824 121828 106880 121884
rect 106880 121828 106884 121884
rect 106820 121824 106884 121828
rect 106900 121884 106964 121888
rect 106900 121828 106904 121884
rect 106904 121828 106960 121884
rect 106960 121828 106964 121884
rect 106900 121824 106964 121828
rect 4216 121340 4280 121344
rect 4216 121284 4220 121340
rect 4220 121284 4276 121340
rect 4276 121284 4280 121340
rect 4216 121280 4280 121284
rect 4296 121340 4360 121344
rect 4296 121284 4300 121340
rect 4300 121284 4356 121340
rect 4356 121284 4360 121340
rect 4296 121280 4360 121284
rect 4376 121340 4440 121344
rect 4376 121284 4380 121340
rect 4380 121284 4436 121340
rect 4436 121284 4440 121340
rect 4376 121280 4440 121284
rect 4456 121340 4520 121344
rect 4456 121284 4460 121340
rect 4460 121284 4516 121340
rect 4516 121284 4520 121340
rect 4456 121280 4520 121284
rect 105924 121340 105988 121344
rect 105924 121284 105928 121340
rect 105928 121284 105984 121340
rect 105984 121284 105988 121340
rect 105924 121280 105988 121284
rect 106004 121340 106068 121344
rect 106004 121284 106008 121340
rect 106008 121284 106064 121340
rect 106064 121284 106068 121340
rect 106004 121280 106068 121284
rect 106084 121340 106148 121344
rect 106084 121284 106088 121340
rect 106088 121284 106144 121340
rect 106144 121284 106148 121340
rect 106084 121280 106148 121284
rect 106164 121340 106228 121344
rect 106164 121284 106168 121340
rect 106168 121284 106224 121340
rect 106224 121284 106228 121340
rect 106164 121280 106228 121284
rect 4876 120796 4940 120800
rect 4876 120740 4880 120796
rect 4880 120740 4936 120796
rect 4936 120740 4940 120796
rect 4876 120736 4940 120740
rect 4956 120796 5020 120800
rect 4956 120740 4960 120796
rect 4960 120740 5016 120796
rect 5016 120740 5020 120796
rect 4956 120736 5020 120740
rect 5036 120796 5100 120800
rect 5036 120740 5040 120796
rect 5040 120740 5096 120796
rect 5096 120740 5100 120796
rect 5036 120736 5100 120740
rect 5116 120796 5180 120800
rect 5116 120740 5120 120796
rect 5120 120740 5176 120796
rect 5176 120740 5180 120796
rect 5116 120736 5180 120740
rect 106660 120796 106724 120800
rect 106660 120740 106664 120796
rect 106664 120740 106720 120796
rect 106720 120740 106724 120796
rect 106660 120736 106724 120740
rect 106740 120796 106804 120800
rect 106740 120740 106744 120796
rect 106744 120740 106800 120796
rect 106800 120740 106804 120796
rect 106740 120736 106804 120740
rect 106820 120796 106884 120800
rect 106820 120740 106824 120796
rect 106824 120740 106880 120796
rect 106880 120740 106884 120796
rect 106820 120736 106884 120740
rect 106900 120796 106964 120800
rect 106900 120740 106904 120796
rect 106904 120740 106960 120796
rect 106960 120740 106964 120796
rect 106900 120736 106964 120740
rect 4216 120252 4280 120256
rect 4216 120196 4220 120252
rect 4220 120196 4276 120252
rect 4276 120196 4280 120252
rect 4216 120192 4280 120196
rect 4296 120252 4360 120256
rect 4296 120196 4300 120252
rect 4300 120196 4356 120252
rect 4356 120196 4360 120252
rect 4296 120192 4360 120196
rect 4376 120252 4440 120256
rect 4376 120196 4380 120252
rect 4380 120196 4436 120252
rect 4436 120196 4440 120252
rect 4376 120192 4440 120196
rect 4456 120252 4520 120256
rect 4456 120196 4460 120252
rect 4460 120196 4516 120252
rect 4516 120196 4520 120252
rect 4456 120192 4520 120196
rect 105924 120252 105988 120256
rect 105924 120196 105928 120252
rect 105928 120196 105984 120252
rect 105984 120196 105988 120252
rect 105924 120192 105988 120196
rect 106004 120252 106068 120256
rect 106004 120196 106008 120252
rect 106008 120196 106064 120252
rect 106064 120196 106068 120252
rect 106004 120192 106068 120196
rect 106084 120252 106148 120256
rect 106084 120196 106088 120252
rect 106088 120196 106144 120252
rect 106144 120196 106148 120252
rect 106084 120192 106148 120196
rect 106164 120252 106228 120256
rect 106164 120196 106168 120252
rect 106168 120196 106224 120252
rect 106224 120196 106228 120252
rect 106164 120192 106228 120196
rect 4876 119708 4940 119712
rect 4876 119652 4880 119708
rect 4880 119652 4936 119708
rect 4936 119652 4940 119708
rect 4876 119648 4940 119652
rect 4956 119708 5020 119712
rect 4956 119652 4960 119708
rect 4960 119652 5016 119708
rect 5016 119652 5020 119708
rect 4956 119648 5020 119652
rect 5036 119708 5100 119712
rect 5036 119652 5040 119708
rect 5040 119652 5096 119708
rect 5096 119652 5100 119708
rect 5036 119648 5100 119652
rect 5116 119708 5180 119712
rect 5116 119652 5120 119708
rect 5120 119652 5176 119708
rect 5176 119652 5180 119708
rect 5116 119648 5180 119652
rect 106660 119708 106724 119712
rect 106660 119652 106664 119708
rect 106664 119652 106720 119708
rect 106720 119652 106724 119708
rect 106660 119648 106724 119652
rect 106740 119708 106804 119712
rect 106740 119652 106744 119708
rect 106744 119652 106800 119708
rect 106800 119652 106804 119708
rect 106740 119648 106804 119652
rect 106820 119708 106884 119712
rect 106820 119652 106824 119708
rect 106824 119652 106880 119708
rect 106880 119652 106884 119708
rect 106820 119648 106884 119652
rect 106900 119708 106964 119712
rect 106900 119652 106904 119708
rect 106904 119652 106960 119708
rect 106960 119652 106964 119708
rect 106900 119648 106964 119652
rect 4216 119164 4280 119168
rect 4216 119108 4220 119164
rect 4220 119108 4276 119164
rect 4276 119108 4280 119164
rect 4216 119104 4280 119108
rect 4296 119164 4360 119168
rect 4296 119108 4300 119164
rect 4300 119108 4356 119164
rect 4356 119108 4360 119164
rect 4296 119104 4360 119108
rect 4376 119164 4440 119168
rect 4376 119108 4380 119164
rect 4380 119108 4436 119164
rect 4436 119108 4440 119164
rect 4376 119104 4440 119108
rect 4456 119164 4520 119168
rect 4456 119108 4460 119164
rect 4460 119108 4516 119164
rect 4516 119108 4520 119164
rect 4456 119104 4520 119108
rect 105924 119164 105988 119168
rect 105924 119108 105928 119164
rect 105928 119108 105984 119164
rect 105984 119108 105988 119164
rect 105924 119104 105988 119108
rect 106004 119164 106068 119168
rect 106004 119108 106008 119164
rect 106008 119108 106064 119164
rect 106064 119108 106068 119164
rect 106004 119104 106068 119108
rect 106084 119164 106148 119168
rect 106084 119108 106088 119164
rect 106088 119108 106144 119164
rect 106144 119108 106148 119164
rect 106084 119104 106148 119108
rect 106164 119164 106228 119168
rect 106164 119108 106168 119164
rect 106168 119108 106224 119164
rect 106224 119108 106228 119164
rect 106164 119104 106228 119108
rect 4876 118620 4940 118624
rect 4876 118564 4880 118620
rect 4880 118564 4936 118620
rect 4936 118564 4940 118620
rect 4876 118560 4940 118564
rect 4956 118620 5020 118624
rect 4956 118564 4960 118620
rect 4960 118564 5016 118620
rect 5016 118564 5020 118620
rect 4956 118560 5020 118564
rect 5036 118620 5100 118624
rect 5036 118564 5040 118620
rect 5040 118564 5096 118620
rect 5096 118564 5100 118620
rect 5036 118560 5100 118564
rect 5116 118620 5180 118624
rect 5116 118564 5120 118620
rect 5120 118564 5176 118620
rect 5176 118564 5180 118620
rect 5116 118560 5180 118564
rect 106660 118620 106724 118624
rect 106660 118564 106664 118620
rect 106664 118564 106720 118620
rect 106720 118564 106724 118620
rect 106660 118560 106724 118564
rect 106740 118620 106804 118624
rect 106740 118564 106744 118620
rect 106744 118564 106800 118620
rect 106800 118564 106804 118620
rect 106740 118560 106804 118564
rect 106820 118620 106884 118624
rect 106820 118564 106824 118620
rect 106824 118564 106880 118620
rect 106880 118564 106884 118620
rect 106820 118560 106884 118564
rect 106900 118620 106964 118624
rect 106900 118564 106904 118620
rect 106904 118564 106960 118620
rect 106960 118564 106964 118620
rect 106900 118560 106964 118564
rect 4216 118076 4280 118080
rect 4216 118020 4220 118076
rect 4220 118020 4276 118076
rect 4276 118020 4280 118076
rect 4216 118016 4280 118020
rect 4296 118076 4360 118080
rect 4296 118020 4300 118076
rect 4300 118020 4356 118076
rect 4356 118020 4360 118076
rect 4296 118016 4360 118020
rect 4376 118076 4440 118080
rect 4376 118020 4380 118076
rect 4380 118020 4436 118076
rect 4436 118020 4440 118076
rect 4376 118016 4440 118020
rect 4456 118076 4520 118080
rect 4456 118020 4460 118076
rect 4460 118020 4516 118076
rect 4516 118020 4520 118076
rect 4456 118016 4520 118020
rect 105924 118076 105988 118080
rect 105924 118020 105928 118076
rect 105928 118020 105984 118076
rect 105984 118020 105988 118076
rect 105924 118016 105988 118020
rect 106004 118076 106068 118080
rect 106004 118020 106008 118076
rect 106008 118020 106064 118076
rect 106064 118020 106068 118076
rect 106004 118016 106068 118020
rect 106084 118076 106148 118080
rect 106084 118020 106088 118076
rect 106088 118020 106144 118076
rect 106144 118020 106148 118076
rect 106084 118016 106148 118020
rect 106164 118076 106228 118080
rect 106164 118020 106168 118076
rect 106168 118020 106224 118076
rect 106224 118020 106228 118076
rect 106164 118016 106228 118020
rect 4876 117532 4940 117536
rect 4876 117476 4880 117532
rect 4880 117476 4936 117532
rect 4936 117476 4940 117532
rect 4876 117472 4940 117476
rect 4956 117532 5020 117536
rect 4956 117476 4960 117532
rect 4960 117476 5016 117532
rect 5016 117476 5020 117532
rect 4956 117472 5020 117476
rect 5036 117532 5100 117536
rect 5036 117476 5040 117532
rect 5040 117476 5096 117532
rect 5096 117476 5100 117532
rect 5036 117472 5100 117476
rect 5116 117532 5180 117536
rect 5116 117476 5120 117532
rect 5120 117476 5176 117532
rect 5176 117476 5180 117532
rect 5116 117472 5180 117476
rect 106660 117532 106724 117536
rect 106660 117476 106664 117532
rect 106664 117476 106720 117532
rect 106720 117476 106724 117532
rect 106660 117472 106724 117476
rect 106740 117532 106804 117536
rect 106740 117476 106744 117532
rect 106744 117476 106800 117532
rect 106800 117476 106804 117532
rect 106740 117472 106804 117476
rect 106820 117532 106884 117536
rect 106820 117476 106824 117532
rect 106824 117476 106880 117532
rect 106880 117476 106884 117532
rect 106820 117472 106884 117476
rect 106900 117532 106964 117536
rect 106900 117476 106904 117532
rect 106904 117476 106960 117532
rect 106960 117476 106964 117532
rect 106900 117472 106964 117476
rect 4216 116988 4280 116992
rect 4216 116932 4220 116988
rect 4220 116932 4276 116988
rect 4276 116932 4280 116988
rect 4216 116928 4280 116932
rect 4296 116988 4360 116992
rect 4296 116932 4300 116988
rect 4300 116932 4356 116988
rect 4356 116932 4360 116988
rect 4296 116928 4360 116932
rect 4376 116988 4440 116992
rect 4376 116932 4380 116988
rect 4380 116932 4436 116988
rect 4436 116932 4440 116988
rect 4376 116928 4440 116932
rect 4456 116988 4520 116992
rect 4456 116932 4460 116988
rect 4460 116932 4516 116988
rect 4516 116932 4520 116988
rect 4456 116928 4520 116932
rect 105924 116988 105988 116992
rect 105924 116932 105928 116988
rect 105928 116932 105984 116988
rect 105984 116932 105988 116988
rect 105924 116928 105988 116932
rect 106004 116988 106068 116992
rect 106004 116932 106008 116988
rect 106008 116932 106064 116988
rect 106064 116932 106068 116988
rect 106004 116928 106068 116932
rect 106084 116988 106148 116992
rect 106084 116932 106088 116988
rect 106088 116932 106144 116988
rect 106144 116932 106148 116988
rect 106084 116928 106148 116932
rect 106164 116988 106228 116992
rect 106164 116932 106168 116988
rect 106168 116932 106224 116988
rect 106224 116932 106228 116988
rect 106164 116928 106228 116932
rect 4876 116444 4940 116448
rect 4876 116388 4880 116444
rect 4880 116388 4936 116444
rect 4936 116388 4940 116444
rect 4876 116384 4940 116388
rect 4956 116444 5020 116448
rect 4956 116388 4960 116444
rect 4960 116388 5016 116444
rect 5016 116388 5020 116444
rect 4956 116384 5020 116388
rect 5036 116444 5100 116448
rect 5036 116388 5040 116444
rect 5040 116388 5096 116444
rect 5096 116388 5100 116444
rect 5036 116384 5100 116388
rect 5116 116444 5180 116448
rect 5116 116388 5120 116444
rect 5120 116388 5176 116444
rect 5176 116388 5180 116444
rect 5116 116384 5180 116388
rect 106660 116444 106724 116448
rect 106660 116388 106664 116444
rect 106664 116388 106720 116444
rect 106720 116388 106724 116444
rect 106660 116384 106724 116388
rect 106740 116444 106804 116448
rect 106740 116388 106744 116444
rect 106744 116388 106800 116444
rect 106800 116388 106804 116444
rect 106740 116384 106804 116388
rect 106820 116444 106884 116448
rect 106820 116388 106824 116444
rect 106824 116388 106880 116444
rect 106880 116388 106884 116444
rect 106820 116384 106884 116388
rect 106900 116444 106964 116448
rect 106900 116388 106904 116444
rect 106904 116388 106960 116444
rect 106960 116388 106964 116444
rect 106900 116384 106964 116388
rect 4216 115900 4280 115904
rect 4216 115844 4220 115900
rect 4220 115844 4276 115900
rect 4276 115844 4280 115900
rect 4216 115840 4280 115844
rect 4296 115900 4360 115904
rect 4296 115844 4300 115900
rect 4300 115844 4356 115900
rect 4356 115844 4360 115900
rect 4296 115840 4360 115844
rect 4376 115900 4440 115904
rect 4376 115844 4380 115900
rect 4380 115844 4436 115900
rect 4436 115844 4440 115900
rect 4376 115840 4440 115844
rect 4456 115900 4520 115904
rect 4456 115844 4460 115900
rect 4460 115844 4516 115900
rect 4516 115844 4520 115900
rect 4456 115840 4520 115844
rect 105924 115900 105988 115904
rect 105924 115844 105928 115900
rect 105928 115844 105984 115900
rect 105984 115844 105988 115900
rect 105924 115840 105988 115844
rect 106004 115900 106068 115904
rect 106004 115844 106008 115900
rect 106008 115844 106064 115900
rect 106064 115844 106068 115900
rect 106004 115840 106068 115844
rect 106084 115900 106148 115904
rect 106084 115844 106088 115900
rect 106088 115844 106144 115900
rect 106144 115844 106148 115900
rect 106084 115840 106148 115844
rect 106164 115900 106228 115904
rect 106164 115844 106168 115900
rect 106168 115844 106224 115900
rect 106224 115844 106228 115900
rect 106164 115840 106228 115844
rect 4876 115356 4940 115360
rect 4876 115300 4880 115356
rect 4880 115300 4936 115356
rect 4936 115300 4940 115356
rect 4876 115296 4940 115300
rect 4956 115356 5020 115360
rect 4956 115300 4960 115356
rect 4960 115300 5016 115356
rect 5016 115300 5020 115356
rect 4956 115296 5020 115300
rect 5036 115356 5100 115360
rect 5036 115300 5040 115356
rect 5040 115300 5096 115356
rect 5096 115300 5100 115356
rect 5036 115296 5100 115300
rect 5116 115356 5180 115360
rect 5116 115300 5120 115356
rect 5120 115300 5176 115356
rect 5176 115300 5180 115356
rect 5116 115296 5180 115300
rect 106660 115356 106724 115360
rect 106660 115300 106664 115356
rect 106664 115300 106720 115356
rect 106720 115300 106724 115356
rect 106660 115296 106724 115300
rect 106740 115356 106804 115360
rect 106740 115300 106744 115356
rect 106744 115300 106800 115356
rect 106800 115300 106804 115356
rect 106740 115296 106804 115300
rect 106820 115356 106884 115360
rect 106820 115300 106824 115356
rect 106824 115300 106880 115356
rect 106880 115300 106884 115356
rect 106820 115296 106884 115300
rect 106900 115356 106964 115360
rect 106900 115300 106904 115356
rect 106904 115300 106960 115356
rect 106960 115300 106964 115356
rect 106900 115296 106964 115300
rect 4216 114812 4280 114816
rect 4216 114756 4220 114812
rect 4220 114756 4276 114812
rect 4276 114756 4280 114812
rect 4216 114752 4280 114756
rect 4296 114812 4360 114816
rect 4296 114756 4300 114812
rect 4300 114756 4356 114812
rect 4356 114756 4360 114812
rect 4296 114752 4360 114756
rect 4376 114812 4440 114816
rect 4376 114756 4380 114812
rect 4380 114756 4436 114812
rect 4436 114756 4440 114812
rect 4376 114752 4440 114756
rect 4456 114812 4520 114816
rect 4456 114756 4460 114812
rect 4460 114756 4516 114812
rect 4516 114756 4520 114812
rect 4456 114752 4520 114756
rect 105924 114812 105988 114816
rect 105924 114756 105928 114812
rect 105928 114756 105984 114812
rect 105984 114756 105988 114812
rect 105924 114752 105988 114756
rect 106004 114812 106068 114816
rect 106004 114756 106008 114812
rect 106008 114756 106064 114812
rect 106064 114756 106068 114812
rect 106004 114752 106068 114756
rect 106084 114812 106148 114816
rect 106084 114756 106088 114812
rect 106088 114756 106144 114812
rect 106144 114756 106148 114812
rect 106084 114752 106148 114756
rect 106164 114812 106228 114816
rect 106164 114756 106168 114812
rect 106168 114756 106224 114812
rect 106224 114756 106228 114812
rect 106164 114752 106228 114756
rect 4876 114268 4940 114272
rect 4876 114212 4880 114268
rect 4880 114212 4936 114268
rect 4936 114212 4940 114268
rect 4876 114208 4940 114212
rect 4956 114268 5020 114272
rect 4956 114212 4960 114268
rect 4960 114212 5016 114268
rect 5016 114212 5020 114268
rect 4956 114208 5020 114212
rect 5036 114268 5100 114272
rect 5036 114212 5040 114268
rect 5040 114212 5096 114268
rect 5096 114212 5100 114268
rect 5036 114208 5100 114212
rect 5116 114268 5180 114272
rect 5116 114212 5120 114268
rect 5120 114212 5176 114268
rect 5176 114212 5180 114268
rect 5116 114208 5180 114212
rect 106660 114268 106724 114272
rect 106660 114212 106664 114268
rect 106664 114212 106720 114268
rect 106720 114212 106724 114268
rect 106660 114208 106724 114212
rect 106740 114268 106804 114272
rect 106740 114212 106744 114268
rect 106744 114212 106800 114268
rect 106800 114212 106804 114268
rect 106740 114208 106804 114212
rect 106820 114268 106884 114272
rect 106820 114212 106824 114268
rect 106824 114212 106880 114268
rect 106880 114212 106884 114268
rect 106820 114208 106884 114212
rect 106900 114268 106964 114272
rect 106900 114212 106904 114268
rect 106904 114212 106960 114268
rect 106960 114212 106964 114268
rect 106900 114208 106964 114212
rect 4216 113724 4280 113728
rect 4216 113668 4220 113724
rect 4220 113668 4276 113724
rect 4276 113668 4280 113724
rect 4216 113664 4280 113668
rect 4296 113724 4360 113728
rect 4296 113668 4300 113724
rect 4300 113668 4356 113724
rect 4356 113668 4360 113724
rect 4296 113664 4360 113668
rect 4376 113724 4440 113728
rect 4376 113668 4380 113724
rect 4380 113668 4436 113724
rect 4436 113668 4440 113724
rect 4376 113664 4440 113668
rect 4456 113724 4520 113728
rect 4456 113668 4460 113724
rect 4460 113668 4516 113724
rect 4516 113668 4520 113724
rect 4456 113664 4520 113668
rect 105924 113724 105988 113728
rect 105924 113668 105928 113724
rect 105928 113668 105984 113724
rect 105984 113668 105988 113724
rect 105924 113664 105988 113668
rect 106004 113724 106068 113728
rect 106004 113668 106008 113724
rect 106008 113668 106064 113724
rect 106064 113668 106068 113724
rect 106004 113664 106068 113668
rect 106084 113724 106148 113728
rect 106084 113668 106088 113724
rect 106088 113668 106144 113724
rect 106144 113668 106148 113724
rect 106084 113664 106148 113668
rect 106164 113724 106228 113728
rect 106164 113668 106168 113724
rect 106168 113668 106224 113724
rect 106224 113668 106228 113724
rect 106164 113664 106228 113668
rect 4876 113180 4940 113184
rect 4876 113124 4880 113180
rect 4880 113124 4936 113180
rect 4936 113124 4940 113180
rect 4876 113120 4940 113124
rect 4956 113180 5020 113184
rect 4956 113124 4960 113180
rect 4960 113124 5016 113180
rect 5016 113124 5020 113180
rect 4956 113120 5020 113124
rect 5036 113180 5100 113184
rect 5036 113124 5040 113180
rect 5040 113124 5096 113180
rect 5096 113124 5100 113180
rect 5036 113120 5100 113124
rect 5116 113180 5180 113184
rect 5116 113124 5120 113180
rect 5120 113124 5176 113180
rect 5176 113124 5180 113180
rect 5116 113120 5180 113124
rect 106660 113180 106724 113184
rect 106660 113124 106664 113180
rect 106664 113124 106720 113180
rect 106720 113124 106724 113180
rect 106660 113120 106724 113124
rect 106740 113180 106804 113184
rect 106740 113124 106744 113180
rect 106744 113124 106800 113180
rect 106800 113124 106804 113180
rect 106740 113120 106804 113124
rect 106820 113180 106884 113184
rect 106820 113124 106824 113180
rect 106824 113124 106880 113180
rect 106880 113124 106884 113180
rect 106820 113120 106884 113124
rect 106900 113180 106964 113184
rect 106900 113124 106904 113180
rect 106904 113124 106960 113180
rect 106960 113124 106964 113180
rect 106900 113120 106964 113124
rect 4216 112636 4280 112640
rect 4216 112580 4220 112636
rect 4220 112580 4276 112636
rect 4276 112580 4280 112636
rect 4216 112576 4280 112580
rect 4296 112636 4360 112640
rect 4296 112580 4300 112636
rect 4300 112580 4356 112636
rect 4356 112580 4360 112636
rect 4296 112576 4360 112580
rect 4376 112636 4440 112640
rect 4376 112580 4380 112636
rect 4380 112580 4436 112636
rect 4436 112580 4440 112636
rect 4376 112576 4440 112580
rect 4456 112636 4520 112640
rect 4456 112580 4460 112636
rect 4460 112580 4516 112636
rect 4516 112580 4520 112636
rect 4456 112576 4520 112580
rect 105924 112636 105988 112640
rect 105924 112580 105928 112636
rect 105928 112580 105984 112636
rect 105984 112580 105988 112636
rect 105924 112576 105988 112580
rect 106004 112636 106068 112640
rect 106004 112580 106008 112636
rect 106008 112580 106064 112636
rect 106064 112580 106068 112636
rect 106004 112576 106068 112580
rect 106084 112636 106148 112640
rect 106084 112580 106088 112636
rect 106088 112580 106144 112636
rect 106144 112580 106148 112636
rect 106084 112576 106148 112580
rect 106164 112636 106228 112640
rect 106164 112580 106168 112636
rect 106168 112580 106224 112636
rect 106224 112580 106228 112636
rect 106164 112576 106228 112580
rect 4876 112092 4940 112096
rect 4876 112036 4880 112092
rect 4880 112036 4936 112092
rect 4936 112036 4940 112092
rect 4876 112032 4940 112036
rect 4956 112092 5020 112096
rect 4956 112036 4960 112092
rect 4960 112036 5016 112092
rect 5016 112036 5020 112092
rect 4956 112032 5020 112036
rect 5036 112092 5100 112096
rect 5036 112036 5040 112092
rect 5040 112036 5096 112092
rect 5096 112036 5100 112092
rect 5036 112032 5100 112036
rect 5116 112092 5180 112096
rect 5116 112036 5120 112092
rect 5120 112036 5176 112092
rect 5176 112036 5180 112092
rect 5116 112032 5180 112036
rect 106660 112092 106724 112096
rect 106660 112036 106664 112092
rect 106664 112036 106720 112092
rect 106720 112036 106724 112092
rect 106660 112032 106724 112036
rect 106740 112092 106804 112096
rect 106740 112036 106744 112092
rect 106744 112036 106800 112092
rect 106800 112036 106804 112092
rect 106740 112032 106804 112036
rect 106820 112092 106884 112096
rect 106820 112036 106824 112092
rect 106824 112036 106880 112092
rect 106880 112036 106884 112092
rect 106820 112032 106884 112036
rect 106900 112092 106964 112096
rect 106900 112036 106904 112092
rect 106904 112036 106960 112092
rect 106960 112036 106964 112092
rect 106900 112032 106964 112036
rect 4216 111548 4280 111552
rect 4216 111492 4220 111548
rect 4220 111492 4276 111548
rect 4276 111492 4280 111548
rect 4216 111488 4280 111492
rect 4296 111548 4360 111552
rect 4296 111492 4300 111548
rect 4300 111492 4356 111548
rect 4356 111492 4360 111548
rect 4296 111488 4360 111492
rect 4376 111548 4440 111552
rect 4376 111492 4380 111548
rect 4380 111492 4436 111548
rect 4436 111492 4440 111548
rect 4376 111488 4440 111492
rect 4456 111548 4520 111552
rect 4456 111492 4460 111548
rect 4460 111492 4516 111548
rect 4516 111492 4520 111548
rect 4456 111488 4520 111492
rect 105924 111548 105988 111552
rect 105924 111492 105928 111548
rect 105928 111492 105984 111548
rect 105984 111492 105988 111548
rect 105924 111488 105988 111492
rect 106004 111548 106068 111552
rect 106004 111492 106008 111548
rect 106008 111492 106064 111548
rect 106064 111492 106068 111548
rect 106004 111488 106068 111492
rect 106084 111548 106148 111552
rect 106084 111492 106088 111548
rect 106088 111492 106144 111548
rect 106144 111492 106148 111548
rect 106084 111488 106148 111492
rect 106164 111548 106228 111552
rect 106164 111492 106168 111548
rect 106168 111492 106224 111548
rect 106224 111492 106228 111548
rect 106164 111488 106228 111492
rect 4876 111004 4940 111008
rect 4876 110948 4880 111004
rect 4880 110948 4936 111004
rect 4936 110948 4940 111004
rect 4876 110944 4940 110948
rect 4956 111004 5020 111008
rect 4956 110948 4960 111004
rect 4960 110948 5016 111004
rect 5016 110948 5020 111004
rect 4956 110944 5020 110948
rect 5036 111004 5100 111008
rect 5036 110948 5040 111004
rect 5040 110948 5096 111004
rect 5096 110948 5100 111004
rect 5036 110944 5100 110948
rect 5116 111004 5180 111008
rect 5116 110948 5120 111004
rect 5120 110948 5176 111004
rect 5176 110948 5180 111004
rect 5116 110944 5180 110948
rect 106660 111004 106724 111008
rect 106660 110948 106664 111004
rect 106664 110948 106720 111004
rect 106720 110948 106724 111004
rect 106660 110944 106724 110948
rect 106740 111004 106804 111008
rect 106740 110948 106744 111004
rect 106744 110948 106800 111004
rect 106800 110948 106804 111004
rect 106740 110944 106804 110948
rect 106820 111004 106884 111008
rect 106820 110948 106824 111004
rect 106824 110948 106880 111004
rect 106880 110948 106884 111004
rect 106820 110944 106884 110948
rect 106900 111004 106964 111008
rect 106900 110948 106904 111004
rect 106904 110948 106960 111004
rect 106960 110948 106964 111004
rect 106900 110944 106964 110948
rect 4216 110460 4280 110464
rect 4216 110404 4220 110460
rect 4220 110404 4276 110460
rect 4276 110404 4280 110460
rect 4216 110400 4280 110404
rect 4296 110460 4360 110464
rect 4296 110404 4300 110460
rect 4300 110404 4356 110460
rect 4356 110404 4360 110460
rect 4296 110400 4360 110404
rect 4376 110460 4440 110464
rect 4376 110404 4380 110460
rect 4380 110404 4436 110460
rect 4436 110404 4440 110460
rect 4376 110400 4440 110404
rect 4456 110460 4520 110464
rect 4456 110404 4460 110460
rect 4460 110404 4516 110460
rect 4516 110404 4520 110460
rect 4456 110400 4520 110404
rect 105924 110460 105988 110464
rect 105924 110404 105928 110460
rect 105928 110404 105984 110460
rect 105984 110404 105988 110460
rect 105924 110400 105988 110404
rect 106004 110460 106068 110464
rect 106004 110404 106008 110460
rect 106008 110404 106064 110460
rect 106064 110404 106068 110460
rect 106004 110400 106068 110404
rect 106084 110460 106148 110464
rect 106084 110404 106088 110460
rect 106088 110404 106144 110460
rect 106144 110404 106148 110460
rect 106084 110400 106148 110404
rect 106164 110460 106228 110464
rect 106164 110404 106168 110460
rect 106168 110404 106224 110460
rect 106224 110404 106228 110460
rect 106164 110400 106228 110404
rect 4876 109916 4940 109920
rect 4876 109860 4880 109916
rect 4880 109860 4936 109916
rect 4936 109860 4940 109916
rect 4876 109856 4940 109860
rect 4956 109916 5020 109920
rect 4956 109860 4960 109916
rect 4960 109860 5016 109916
rect 5016 109860 5020 109916
rect 4956 109856 5020 109860
rect 5036 109916 5100 109920
rect 5036 109860 5040 109916
rect 5040 109860 5096 109916
rect 5096 109860 5100 109916
rect 5036 109856 5100 109860
rect 5116 109916 5180 109920
rect 5116 109860 5120 109916
rect 5120 109860 5176 109916
rect 5176 109860 5180 109916
rect 5116 109856 5180 109860
rect 106660 109916 106724 109920
rect 106660 109860 106664 109916
rect 106664 109860 106720 109916
rect 106720 109860 106724 109916
rect 106660 109856 106724 109860
rect 106740 109916 106804 109920
rect 106740 109860 106744 109916
rect 106744 109860 106800 109916
rect 106800 109860 106804 109916
rect 106740 109856 106804 109860
rect 106820 109916 106884 109920
rect 106820 109860 106824 109916
rect 106824 109860 106880 109916
rect 106880 109860 106884 109916
rect 106820 109856 106884 109860
rect 106900 109916 106964 109920
rect 106900 109860 106904 109916
rect 106904 109860 106960 109916
rect 106960 109860 106964 109916
rect 106900 109856 106964 109860
rect 4216 109372 4280 109376
rect 4216 109316 4220 109372
rect 4220 109316 4276 109372
rect 4276 109316 4280 109372
rect 4216 109312 4280 109316
rect 4296 109372 4360 109376
rect 4296 109316 4300 109372
rect 4300 109316 4356 109372
rect 4356 109316 4360 109372
rect 4296 109312 4360 109316
rect 4376 109372 4440 109376
rect 4376 109316 4380 109372
rect 4380 109316 4436 109372
rect 4436 109316 4440 109372
rect 4376 109312 4440 109316
rect 4456 109372 4520 109376
rect 4456 109316 4460 109372
rect 4460 109316 4516 109372
rect 4516 109316 4520 109372
rect 4456 109312 4520 109316
rect 105924 109372 105988 109376
rect 105924 109316 105928 109372
rect 105928 109316 105984 109372
rect 105984 109316 105988 109372
rect 105924 109312 105988 109316
rect 106004 109372 106068 109376
rect 106004 109316 106008 109372
rect 106008 109316 106064 109372
rect 106064 109316 106068 109372
rect 106004 109312 106068 109316
rect 106084 109372 106148 109376
rect 106084 109316 106088 109372
rect 106088 109316 106144 109372
rect 106144 109316 106148 109372
rect 106084 109312 106148 109316
rect 106164 109372 106228 109376
rect 106164 109316 106168 109372
rect 106168 109316 106224 109372
rect 106224 109316 106228 109372
rect 106164 109312 106228 109316
rect 4876 108828 4940 108832
rect 4876 108772 4880 108828
rect 4880 108772 4936 108828
rect 4936 108772 4940 108828
rect 4876 108768 4940 108772
rect 4956 108828 5020 108832
rect 4956 108772 4960 108828
rect 4960 108772 5016 108828
rect 5016 108772 5020 108828
rect 4956 108768 5020 108772
rect 5036 108828 5100 108832
rect 5036 108772 5040 108828
rect 5040 108772 5096 108828
rect 5096 108772 5100 108828
rect 5036 108768 5100 108772
rect 5116 108828 5180 108832
rect 5116 108772 5120 108828
rect 5120 108772 5176 108828
rect 5176 108772 5180 108828
rect 5116 108768 5180 108772
rect 106660 108828 106724 108832
rect 106660 108772 106664 108828
rect 106664 108772 106720 108828
rect 106720 108772 106724 108828
rect 106660 108768 106724 108772
rect 106740 108828 106804 108832
rect 106740 108772 106744 108828
rect 106744 108772 106800 108828
rect 106800 108772 106804 108828
rect 106740 108768 106804 108772
rect 106820 108828 106884 108832
rect 106820 108772 106824 108828
rect 106824 108772 106880 108828
rect 106880 108772 106884 108828
rect 106820 108768 106884 108772
rect 106900 108828 106964 108832
rect 106900 108772 106904 108828
rect 106904 108772 106960 108828
rect 106960 108772 106964 108828
rect 106900 108768 106964 108772
rect 4216 108284 4280 108288
rect 4216 108228 4220 108284
rect 4220 108228 4276 108284
rect 4276 108228 4280 108284
rect 4216 108224 4280 108228
rect 4296 108284 4360 108288
rect 4296 108228 4300 108284
rect 4300 108228 4356 108284
rect 4356 108228 4360 108284
rect 4296 108224 4360 108228
rect 4376 108284 4440 108288
rect 4376 108228 4380 108284
rect 4380 108228 4436 108284
rect 4436 108228 4440 108284
rect 4376 108224 4440 108228
rect 4456 108284 4520 108288
rect 4456 108228 4460 108284
rect 4460 108228 4516 108284
rect 4516 108228 4520 108284
rect 4456 108224 4520 108228
rect 105924 108284 105988 108288
rect 105924 108228 105928 108284
rect 105928 108228 105984 108284
rect 105984 108228 105988 108284
rect 105924 108224 105988 108228
rect 106004 108284 106068 108288
rect 106004 108228 106008 108284
rect 106008 108228 106064 108284
rect 106064 108228 106068 108284
rect 106004 108224 106068 108228
rect 106084 108284 106148 108288
rect 106084 108228 106088 108284
rect 106088 108228 106144 108284
rect 106144 108228 106148 108284
rect 106084 108224 106148 108228
rect 106164 108284 106228 108288
rect 106164 108228 106168 108284
rect 106168 108228 106224 108284
rect 106224 108228 106228 108284
rect 106164 108224 106228 108228
rect 4876 107740 4940 107744
rect 4876 107684 4880 107740
rect 4880 107684 4936 107740
rect 4936 107684 4940 107740
rect 4876 107680 4940 107684
rect 4956 107740 5020 107744
rect 4956 107684 4960 107740
rect 4960 107684 5016 107740
rect 5016 107684 5020 107740
rect 4956 107680 5020 107684
rect 5036 107740 5100 107744
rect 5036 107684 5040 107740
rect 5040 107684 5096 107740
rect 5096 107684 5100 107740
rect 5036 107680 5100 107684
rect 5116 107740 5180 107744
rect 5116 107684 5120 107740
rect 5120 107684 5176 107740
rect 5176 107684 5180 107740
rect 5116 107680 5180 107684
rect 106660 107740 106724 107744
rect 106660 107684 106664 107740
rect 106664 107684 106720 107740
rect 106720 107684 106724 107740
rect 106660 107680 106724 107684
rect 106740 107740 106804 107744
rect 106740 107684 106744 107740
rect 106744 107684 106800 107740
rect 106800 107684 106804 107740
rect 106740 107680 106804 107684
rect 106820 107740 106884 107744
rect 106820 107684 106824 107740
rect 106824 107684 106880 107740
rect 106880 107684 106884 107740
rect 106820 107680 106884 107684
rect 106900 107740 106964 107744
rect 106900 107684 106904 107740
rect 106904 107684 106960 107740
rect 106960 107684 106964 107740
rect 106900 107680 106964 107684
rect 4216 107196 4280 107200
rect 4216 107140 4220 107196
rect 4220 107140 4276 107196
rect 4276 107140 4280 107196
rect 4216 107136 4280 107140
rect 4296 107196 4360 107200
rect 4296 107140 4300 107196
rect 4300 107140 4356 107196
rect 4356 107140 4360 107196
rect 4296 107136 4360 107140
rect 4376 107196 4440 107200
rect 4376 107140 4380 107196
rect 4380 107140 4436 107196
rect 4436 107140 4440 107196
rect 4376 107136 4440 107140
rect 4456 107196 4520 107200
rect 4456 107140 4460 107196
rect 4460 107140 4516 107196
rect 4516 107140 4520 107196
rect 4456 107136 4520 107140
rect 105924 107196 105988 107200
rect 105924 107140 105928 107196
rect 105928 107140 105984 107196
rect 105984 107140 105988 107196
rect 105924 107136 105988 107140
rect 106004 107196 106068 107200
rect 106004 107140 106008 107196
rect 106008 107140 106064 107196
rect 106064 107140 106068 107196
rect 106004 107136 106068 107140
rect 106084 107196 106148 107200
rect 106084 107140 106088 107196
rect 106088 107140 106144 107196
rect 106144 107140 106148 107196
rect 106084 107136 106148 107140
rect 106164 107196 106228 107200
rect 106164 107140 106168 107196
rect 106168 107140 106224 107196
rect 106224 107140 106228 107196
rect 106164 107136 106228 107140
rect 4876 106652 4940 106656
rect 4876 106596 4880 106652
rect 4880 106596 4936 106652
rect 4936 106596 4940 106652
rect 4876 106592 4940 106596
rect 4956 106652 5020 106656
rect 4956 106596 4960 106652
rect 4960 106596 5016 106652
rect 5016 106596 5020 106652
rect 4956 106592 5020 106596
rect 5036 106652 5100 106656
rect 5036 106596 5040 106652
rect 5040 106596 5096 106652
rect 5096 106596 5100 106652
rect 5036 106592 5100 106596
rect 5116 106652 5180 106656
rect 5116 106596 5120 106652
rect 5120 106596 5176 106652
rect 5176 106596 5180 106652
rect 5116 106592 5180 106596
rect 106660 106652 106724 106656
rect 106660 106596 106664 106652
rect 106664 106596 106720 106652
rect 106720 106596 106724 106652
rect 106660 106592 106724 106596
rect 106740 106652 106804 106656
rect 106740 106596 106744 106652
rect 106744 106596 106800 106652
rect 106800 106596 106804 106652
rect 106740 106592 106804 106596
rect 106820 106652 106884 106656
rect 106820 106596 106824 106652
rect 106824 106596 106880 106652
rect 106880 106596 106884 106652
rect 106820 106592 106884 106596
rect 106900 106652 106964 106656
rect 106900 106596 106904 106652
rect 106904 106596 106960 106652
rect 106960 106596 106964 106652
rect 106900 106592 106964 106596
rect 4216 106108 4280 106112
rect 4216 106052 4220 106108
rect 4220 106052 4276 106108
rect 4276 106052 4280 106108
rect 4216 106048 4280 106052
rect 4296 106108 4360 106112
rect 4296 106052 4300 106108
rect 4300 106052 4356 106108
rect 4356 106052 4360 106108
rect 4296 106048 4360 106052
rect 4376 106108 4440 106112
rect 4376 106052 4380 106108
rect 4380 106052 4436 106108
rect 4436 106052 4440 106108
rect 4376 106048 4440 106052
rect 4456 106108 4520 106112
rect 4456 106052 4460 106108
rect 4460 106052 4516 106108
rect 4516 106052 4520 106108
rect 4456 106048 4520 106052
rect 105924 106108 105988 106112
rect 105924 106052 105928 106108
rect 105928 106052 105984 106108
rect 105984 106052 105988 106108
rect 105924 106048 105988 106052
rect 106004 106108 106068 106112
rect 106004 106052 106008 106108
rect 106008 106052 106064 106108
rect 106064 106052 106068 106108
rect 106004 106048 106068 106052
rect 106084 106108 106148 106112
rect 106084 106052 106088 106108
rect 106088 106052 106144 106108
rect 106144 106052 106148 106108
rect 106084 106048 106148 106052
rect 106164 106108 106228 106112
rect 106164 106052 106168 106108
rect 106168 106052 106224 106108
rect 106224 106052 106228 106108
rect 106164 106048 106228 106052
rect 4876 105564 4940 105568
rect 4876 105508 4880 105564
rect 4880 105508 4936 105564
rect 4936 105508 4940 105564
rect 4876 105504 4940 105508
rect 4956 105564 5020 105568
rect 4956 105508 4960 105564
rect 4960 105508 5016 105564
rect 5016 105508 5020 105564
rect 4956 105504 5020 105508
rect 5036 105564 5100 105568
rect 5036 105508 5040 105564
rect 5040 105508 5096 105564
rect 5096 105508 5100 105564
rect 5036 105504 5100 105508
rect 5116 105564 5180 105568
rect 5116 105508 5120 105564
rect 5120 105508 5176 105564
rect 5176 105508 5180 105564
rect 5116 105504 5180 105508
rect 106660 105564 106724 105568
rect 106660 105508 106664 105564
rect 106664 105508 106720 105564
rect 106720 105508 106724 105564
rect 106660 105504 106724 105508
rect 106740 105564 106804 105568
rect 106740 105508 106744 105564
rect 106744 105508 106800 105564
rect 106800 105508 106804 105564
rect 106740 105504 106804 105508
rect 106820 105564 106884 105568
rect 106820 105508 106824 105564
rect 106824 105508 106880 105564
rect 106880 105508 106884 105564
rect 106820 105504 106884 105508
rect 106900 105564 106964 105568
rect 106900 105508 106904 105564
rect 106904 105508 106960 105564
rect 106960 105508 106964 105564
rect 106900 105504 106964 105508
rect 4216 105020 4280 105024
rect 4216 104964 4220 105020
rect 4220 104964 4276 105020
rect 4276 104964 4280 105020
rect 4216 104960 4280 104964
rect 4296 105020 4360 105024
rect 4296 104964 4300 105020
rect 4300 104964 4356 105020
rect 4356 104964 4360 105020
rect 4296 104960 4360 104964
rect 4376 105020 4440 105024
rect 4376 104964 4380 105020
rect 4380 104964 4436 105020
rect 4436 104964 4440 105020
rect 4376 104960 4440 104964
rect 4456 105020 4520 105024
rect 4456 104964 4460 105020
rect 4460 104964 4516 105020
rect 4516 104964 4520 105020
rect 4456 104960 4520 104964
rect 105924 105020 105988 105024
rect 105924 104964 105928 105020
rect 105928 104964 105984 105020
rect 105984 104964 105988 105020
rect 105924 104960 105988 104964
rect 106004 105020 106068 105024
rect 106004 104964 106008 105020
rect 106008 104964 106064 105020
rect 106064 104964 106068 105020
rect 106004 104960 106068 104964
rect 106084 105020 106148 105024
rect 106084 104964 106088 105020
rect 106088 104964 106144 105020
rect 106144 104964 106148 105020
rect 106084 104960 106148 104964
rect 106164 105020 106228 105024
rect 106164 104964 106168 105020
rect 106168 104964 106224 105020
rect 106224 104964 106228 105020
rect 106164 104960 106228 104964
rect 4876 104476 4940 104480
rect 4876 104420 4880 104476
rect 4880 104420 4936 104476
rect 4936 104420 4940 104476
rect 4876 104416 4940 104420
rect 4956 104476 5020 104480
rect 4956 104420 4960 104476
rect 4960 104420 5016 104476
rect 5016 104420 5020 104476
rect 4956 104416 5020 104420
rect 5036 104476 5100 104480
rect 5036 104420 5040 104476
rect 5040 104420 5096 104476
rect 5096 104420 5100 104476
rect 5036 104416 5100 104420
rect 5116 104476 5180 104480
rect 5116 104420 5120 104476
rect 5120 104420 5176 104476
rect 5176 104420 5180 104476
rect 5116 104416 5180 104420
rect 106660 104476 106724 104480
rect 106660 104420 106664 104476
rect 106664 104420 106720 104476
rect 106720 104420 106724 104476
rect 106660 104416 106724 104420
rect 106740 104476 106804 104480
rect 106740 104420 106744 104476
rect 106744 104420 106800 104476
rect 106800 104420 106804 104476
rect 106740 104416 106804 104420
rect 106820 104476 106884 104480
rect 106820 104420 106824 104476
rect 106824 104420 106880 104476
rect 106880 104420 106884 104476
rect 106820 104416 106884 104420
rect 106900 104476 106964 104480
rect 106900 104420 106904 104476
rect 106904 104420 106960 104476
rect 106960 104420 106964 104476
rect 106900 104416 106964 104420
rect 4216 103932 4280 103936
rect 4216 103876 4220 103932
rect 4220 103876 4276 103932
rect 4276 103876 4280 103932
rect 4216 103872 4280 103876
rect 4296 103932 4360 103936
rect 4296 103876 4300 103932
rect 4300 103876 4356 103932
rect 4356 103876 4360 103932
rect 4296 103872 4360 103876
rect 4376 103932 4440 103936
rect 4376 103876 4380 103932
rect 4380 103876 4436 103932
rect 4436 103876 4440 103932
rect 4376 103872 4440 103876
rect 4456 103932 4520 103936
rect 4456 103876 4460 103932
rect 4460 103876 4516 103932
rect 4516 103876 4520 103932
rect 4456 103872 4520 103876
rect 105924 103932 105988 103936
rect 105924 103876 105928 103932
rect 105928 103876 105984 103932
rect 105984 103876 105988 103932
rect 105924 103872 105988 103876
rect 106004 103932 106068 103936
rect 106004 103876 106008 103932
rect 106008 103876 106064 103932
rect 106064 103876 106068 103932
rect 106004 103872 106068 103876
rect 106084 103932 106148 103936
rect 106084 103876 106088 103932
rect 106088 103876 106144 103932
rect 106144 103876 106148 103932
rect 106084 103872 106148 103876
rect 106164 103932 106228 103936
rect 106164 103876 106168 103932
rect 106168 103876 106224 103932
rect 106224 103876 106228 103932
rect 106164 103872 106228 103876
rect 4876 103388 4940 103392
rect 4876 103332 4880 103388
rect 4880 103332 4936 103388
rect 4936 103332 4940 103388
rect 4876 103328 4940 103332
rect 4956 103388 5020 103392
rect 4956 103332 4960 103388
rect 4960 103332 5016 103388
rect 5016 103332 5020 103388
rect 4956 103328 5020 103332
rect 5036 103388 5100 103392
rect 5036 103332 5040 103388
rect 5040 103332 5096 103388
rect 5096 103332 5100 103388
rect 5036 103328 5100 103332
rect 5116 103388 5180 103392
rect 5116 103332 5120 103388
rect 5120 103332 5176 103388
rect 5176 103332 5180 103388
rect 5116 103328 5180 103332
rect 106660 103388 106724 103392
rect 106660 103332 106664 103388
rect 106664 103332 106720 103388
rect 106720 103332 106724 103388
rect 106660 103328 106724 103332
rect 106740 103388 106804 103392
rect 106740 103332 106744 103388
rect 106744 103332 106800 103388
rect 106800 103332 106804 103388
rect 106740 103328 106804 103332
rect 106820 103388 106884 103392
rect 106820 103332 106824 103388
rect 106824 103332 106880 103388
rect 106880 103332 106884 103388
rect 106820 103328 106884 103332
rect 106900 103388 106964 103392
rect 106900 103332 106904 103388
rect 106904 103332 106960 103388
rect 106960 103332 106964 103388
rect 106900 103328 106964 103332
rect 4216 102844 4280 102848
rect 4216 102788 4220 102844
rect 4220 102788 4276 102844
rect 4276 102788 4280 102844
rect 4216 102784 4280 102788
rect 4296 102844 4360 102848
rect 4296 102788 4300 102844
rect 4300 102788 4356 102844
rect 4356 102788 4360 102844
rect 4296 102784 4360 102788
rect 4376 102844 4440 102848
rect 4376 102788 4380 102844
rect 4380 102788 4436 102844
rect 4436 102788 4440 102844
rect 4376 102784 4440 102788
rect 4456 102844 4520 102848
rect 4456 102788 4460 102844
rect 4460 102788 4516 102844
rect 4516 102788 4520 102844
rect 4456 102784 4520 102788
rect 105924 102844 105988 102848
rect 105924 102788 105928 102844
rect 105928 102788 105984 102844
rect 105984 102788 105988 102844
rect 105924 102784 105988 102788
rect 106004 102844 106068 102848
rect 106004 102788 106008 102844
rect 106008 102788 106064 102844
rect 106064 102788 106068 102844
rect 106004 102784 106068 102788
rect 106084 102844 106148 102848
rect 106084 102788 106088 102844
rect 106088 102788 106144 102844
rect 106144 102788 106148 102844
rect 106084 102784 106148 102788
rect 106164 102844 106228 102848
rect 106164 102788 106168 102844
rect 106168 102788 106224 102844
rect 106224 102788 106228 102844
rect 106164 102784 106228 102788
rect 4876 102300 4940 102304
rect 4876 102244 4880 102300
rect 4880 102244 4936 102300
rect 4936 102244 4940 102300
rect 4876 102240 4940 102244
rect 4956 102300 5020 102304
rect 4956 102244 4960 102300
rect 4960 102244 5016 102300
rect 5016 102244 5020 102300
rect 4956 102240 5020 102244
rect 5036 102300 5100 102304
rect 5036 102244 5040 102300
rect 5040 102244 5096 102300
rect 5096 102244 5100 102300
rect 5036 102240 5100 102244
rect 5116 102300 5180 102304
rect 5116 102244 5120 102300
rect 5120 102244 5176 102300
rect 5176 102244 5180 102300
rect 5116 102240 5180 102244
rect 106660 102300 106724 102304
rect 106660 102244 106664 102300
rect 106664 102244 106720 102300
rect 106720 102244 106724 102300
rect 106660 102240 106724 102244
rect 106740 102300 106804 102304
rect 106740 102244 106744 102300
rect 106744 102244 106800 102300
rect 106800 102244 106804 102300
rect 106740 102240 106804 102244
rect 106820 102300 106884 102304
rect 106820 102244 106824 102300
rect 106824 102244 106880 102300
rect 106880 102244 106884 102300
rect 106820 102240 106884 102244
rect 106900 102300 106964 102304
rect 106900 102244 106904 102300
rect 106904 102244 106960 102300
rect 106960 102244 106964 102300
rect 106900 102240 106964 102244
rect 4216 101756 4280 101760
rect 4216 101700 4220 101756
rect 4220 101700 4276 101756
rect 4276 101700 4280 101756
rect 4216 101696 4280 101700
rect 4296 101756 4360 101760
rect 4296 101700 4300 101756
rect 4300 101700 4356 101756
rect 4356 101700 4360 101756
rect 4296 101696 4360 101700
rect 4376 101756 4440 101760
rect 4376 101700 4380 101756
rect 4380 101700 4436 101756
rect 4436 101700 4440 101756
rect 4376 101696 4440 101700
rect 4456 101756 4520 101760
rect 4456 101700 4460 101756
rect 4460 101700 4516 101756
rect 4516 101700 4520 101756
rect 4456 101696 4520 101700
rect 105924 101756 105988 101760
rect 105924 101700 105928 101756
rect 105928 101700 105984 101756
rect 105984 101700 105988 101756
rect 105924 101696 105988 101700
rect 106004 101756 106068 101760
rect 106004 101700 106008 101756
rect 106008 101700 106064 101756
rect 106064 101700 106068 101756
rect 106004 101696 106068 101700
rect 106084 101756 106148 101760
rect 106084 101700 106088 101756
rect 106088 101700 106144 101756
rect 106144 101700 106148 101756
rect 106084 101696 106148 101700
rect 106164 101756 106228 101760
rect 106164 101700 106168 101756
rect 106168 101700 106224 101756
rect 106224 101700 106228 101756
rect 106164 101696 106228 101700
rect 4876 101212 4940 101216
rect 4876 101156 4880 101212
rect 4880 101156 4936 101212
rect 4936 101156 4940 101212
rect 4876 101152 4940 101156
rect 4956 101212 5020 101216
rect 4956 101156 4960 101212
rect 4960 101156 5016 101212
rect 5016 101156 5020 101212
rect 4956 101152 5020 101156
rect 5036 101212 5100 101216
rect 5036 101156 5040 101212
rect 5040 101156 5096 101212
rect 5096 101156 5100 101212
rect 5036 101152 5100 101156
rect 5116 101212 5180 101216
rect 5116 101156 5120 101212
rect 5120 101156 5176 101212
rect 5176 101156 5180 101212
rect 5116 101152 5180 101156
rect 106660 101212 106724 101216
rect 106660 101156 106664 101212
rect 106664 101156 106720 101212
rect 106720 101156 106724 101212
rect 106660 101152 106724 101156
rect 106740 101212 106804 101216
rect 106740 101156 106744 101212
rect 106744 101156 106800 101212
rect 106800 101156 106804 101212
rect 106740 101152 106804 101156
rect 106820 101212 106884 101216
rect 106820 101156 106824 101212
rect 106824 101156 106880 101212
rect 106880 101156 106884 101212
rect 106820 101152 106884 101156
rect 106900 101212 106964 101216
rect 106900 101156 106904 101212
rect 106904 101156 106960 101212
rect 106960 101156 106964 101212
rect 106900 101152 106964 101156
rect 4216 100668 4280 100672
rect 4216 100612 4220 100668
rect 4220 100612 4276 100668
rect 4276 100612 4280 100668
rect 4216 100608 4280 100612
rect 4296 100668 4360 100672
rect 4296 100612 4300 100668
rect 4300 100612 4356 100668
rect 4356 100612 4360 100668
rect 4296 100608 4360 100612
rect 4376 100668 4440 100672
rect 4376 100612 4380 100668
rect 4380 100612 4436 100668
rect 4436 100612 4440 100668
rect 4376 100608 4440 100612
rect 4456 100668 4520 100672
rect 4456 100612 4460 100668
rect 4460 100612 4516 100668
rect 4516 100612 4520 100668
rect 4456 100608 4520 100612
rect 105924 100668 105988 100672
rect 105924 100612 105928 100668
rect 105928 100612 105984 100668
rect 105984 100612 105988 100668
rect 105924 100608 105988 100612
rect 106004 100668 106068 100672
rect 106004 100612 106008 100668
rect 106008 100612 106064 100668
rect 106064 100612 106068 100668
rect 106004 100608 106068 100612
rect 106084 100668 106148 100672
rect 106084 100612 106088 100668
rect 106088 100612 106144 100668
rect 106144 100612 106148 100668
rect 106084 100608 106148 100612
rect 106164 100668 106228 100672
rect 106164 100612 106168 100668
rect 106168 100612 106224 100668
rect 106224 100612 106228 100668
rect 106164 100608 106228 100612
rect 4876 100124 4940 100128
rect 4876 100068 4880 100124
rect 4880 100068 4936 100124
rect 4936 100068 4940 100124
rect 4876 100064 4940 100068
rect 4956 100124 5020 100128
rect 4956 100068 4960 100124
rect 4960 100068 5016 100124
rect 5016 100068 5020 100124
rect 4956 100064 5020 100068
rect 5036 100124 5100 100128
rect 5036 100068 5040 100124
rect 5040 100068 5096 100124
rect 5096 100068 5100 100124
rect 5036 100064 5100 100068
rect 5116 100124 5180 100128
rect 5116 100068 5120 100124
rect 5120 100068 5176 100124
rect 5176 100068 5180 100124
rect 5116 100064 5180 100068
rect 106660 100124 106724 100128
rect 106660 100068 106664 100124
rect 106664 100068 106720 100124
rect 106720 100068 106724 100124
rect 106660 100064 106724 100068
rect 106740 100124 106804 100128
rect 106740 100068 106744 100124
rect 106744 100068 106800 100124
rect 106800 100068 106804 100124
rect 106740 100064 106804 100068
rect 106820 100124 106884 100128
rect 106820 100068 106824 100124
rect 106824 100068 106880 100124
rect 106880 100068 106884 100124
rect 106820 100064 106884 100068
rect 106900 100124 106964 100128
rect 106900 100068 106904 100124
rect 106904 100068 106960 100124
rect 106960 100068 106964 100124
rect 106900 100064 106964 100068
rect 4216 99580 4280 99584
rect 4216 99524 4220 99580
rect 4220 99524 4276 99580
rect 4276 99524 4280 99580
rect 4216 99520 4280 99524
rect 4296 99580 4360 99584
rect 4296 99524 4300 99580
rect 4300 99524 4356 99580
rect 4356 99524 4360 99580
rect 4296 99520 4360 99524
rect 4376 99580 4440 99584
rect 4376 99524 4380 99580
rect 4380 99524 4436 99580
rect 4436 99524 4440 99580
rect 4376 99520 4440 99524
rect 4456 99580 4520 99584
rect 4456 99524 4460 99580
rect 4460 99524 4516 99580
rect 4516 99524 4520 99580
rect 4456 99520 4520 99524
rect 105924 99580 105988 99584
rect 105924 99524 105928 99580
rect 105928 99524 105984 99580
rect 105984 99524 105988 99580
rect 105924 99520 105988 99524
rect 106004 99580 106068 99584
rect 106004 99524 106008 99580
rect 106008 99524 106064 99580
rect 106064 99524 106068 99580
rect 106004 99520 106068 99524
rect 106084 99580 106148 99584
rect 106084 99524 106088 99580
rect 106088 99524 106144 99580
rect 106144 99524 106148 99580
rect 106084 99520 106148 99524
rect 106164 99580 106228 99584
rect 106164 99524 106168 99580
rect 106168 99524 106224 99580
rect 106224 99524 106228 99580
rect 106164 99520 106228 99524
rect 4876 99036 4940 99040
rect 4876 98980 4880 99036
rect 4880 98980 4936 99036
rect 4936 98980 4940 99036
rect 4876 98976 4940 98980
rect 4956 99036 5020 99040
rect 4956 98980 4960 99036
rect 4960 98980 5016 99036
rect 5016 98980 5020 99036
rect 4956 98976 5020 98980
rect 5036 99036 5100 99040
rect 5036 98980 5040 99036
rect 5040 98980 5096 99036
rect 5096 98980 5100 99036
rect 5036 98976 5100 98980
rect 5116 99036 5180 99040
rect 5116 98980 5120 99036
rect 5120 98980 5176 99036
rect 5176 98980 5180 99036
rect 5116 98976 5180 98980
rect 106660 99036 106724 99040
rect 106660 98980 106664 99036
rect 106664 98980 106720 99036
rect 106720 98980 106724 99036
rect 106660 98976 106724 98980
rect 106740 99036 106804 99040
rect 106740 98980 106744 99036
rect 106744 98980 106800 99036
rect 106800 98980 106804 99036
rect 106740 98976 106804 98980
rect 106820 99036 106884 99040
rect 106820 98980 106824 99036
rect 106824 98980 106880 99036
rect 106880 98980 106884 99036
rect 106820 98976 106884 98980
rect 106900 99036 106964 99040
rect 106900 98980 106904 99036
rect 106904 98980 106960 99036
rect 106960 98980 106964 99036
rect 106900 98976 106964 98980
rect 4216 98492 4280 98496
rect 4216 98436 4220 98492
rect 4220 98436 4276 98492
rect 4276 98436 4280 98492
rect 4216 98432 4280 98436
rect 4296 98492 4360 98496
rect 4296 98436 4300 98492
rect 4300 98436 4356 98492
rect 4356 98436 4360 98492
rect 4296 98432 4360 98436
rect 4376 98492 4440 98496
rect 4376 98436 4380 98492
rect 4380 98436 4436 98492
rect 4436 98436 4440 98492
rect 4376 98432 4440 98436
rect 4456 98492 4520 98496
rect 4456 98436 4460 98492
rect 4460 98436 4516 98492
rect 4516 98436 4520 98492
rect 4456 98432 4520 98436
rect 105924 98492 105988 98496
rect 105924 98436 105928 98492
rect 105928 98436 105984 98492
rect 105984 98436 105988 98492
rect 105924 98432 105988 98436
rect 106004 98492 106068 98496
rect 106004 98436 106008 98492
rect 106008 98436 106064 98492
rect 106064 98436 106068 98492
rect 106004 98432 106068 98436
rect 106084 98492 106148 98496
rect 106084 98436 106088 98492
rect 106088 98436 106144 98492
rect 106144 98436 106148 98492
rect 106084 98432 106148 98436
rect 106164 98492 106228 98496
rect 106164 98436 106168 98492
rect 106168 98436 106224 98492
rect 106224 98436 106228 98492
rect 106164 98432 106228 98436
rect 4876 97948 4940 97952
rect 4876 97892 4880 97948
rect 4880 97892 4936 97948
rect 4936 97892 4940 97948
rect 4876 97888 4940 97892
rect 4956 97948 5020 97952
rect 4956 97892 4960 97948
rect 4960 97892 5016 97948
rect 5016 97892 5020 97948
rect 4956 97888 5020 97892
rect 5036 97948 5100 97952
rect 5036 97892 5040 97948
rect 5040 97892 5096 97948
rect 5096 97892 5100 97948
rect 5036 97888 5100 97892
rect 5116 97948 5180 97952
rect 5116 97892 5120 97948
rect 5120 97892 5176 97948
rect 5176 97892 5180 97948
rect 5116 97888 5180 97892
rect 106660 97948 106724 97952
rect 106660 97892 106664 97948
rect 106664 97892 106720 97948
rect 106720 97892 106724 97948
rect 106660 97888 106724 97892
rect 106740 97948 106804 97952
rect 106740 97892 106744 97948
rect 106744 97892 106800 97948
rect 106800 97892 106804 97948
rect 106740 97888 106804 97892
rect 106820 97948 106884 97952
rect 106820 97892 106824 97948
rect 106824 97892 106880 97948
rect 106880 97892 106884 97948
rect 106820 97888 106884 97892
rect 106900 97948 106964 97952
rect 106900 97892 106904 97948
rect 106904 97892 106960 97948
rect 106960 97892 106964 97948
rect 106900 97888 106964 97892
rect 4216 97404 4280 97408
rect 4216 97348 4220 97404
rect 4220 97348 4276 97404
rect 4276 97348 4280 97404
rect 4216 97344 4280 97348
rect 4296 97404 4360 97408
rect 4296 97348 4300 97404
rect 4300 97348 4356 97404
rect 4356 97348 4360 97404
rect 4296 97344 4360 97348
rect 4376 97404 4440 97408
rect 4376 97348 4380 97404
rect 4380 97348 4436 97404
rect 4436 97348 4440 97404
rect 4376 97344 4440 97348
rect 4456 97404 4520 97408
rect 4456 97348 4460 97404
rect 4460 97348 4516 97404
rect 4516 97348 4520 97404
rect 4456 97344 4520 97348
rect 105924 97404 105988 97408
rect 105924 97348 105928 97404
rect 105928 97348 105984 97404
rect 105984 97348 105988 97404
rect 105924 97344 105988 97348
rect 106004 97404 106068 97408
rect 106004 97348 106008 97404
rect 106008 97348 106064 97404
rect 106064 97348 106068 97404
rect 106004 97344 106068 97348
rect 106084 97404 106148 97408
rect 106084 97348 106088 97404
rect 106088 97348 106144 97404
rect 106144 97348 106148 97404
rect 106084 97344 106148 97348
rect 106164 97404 106228 97408
rect 106164 97348 106168 97404
rect 106168 97348 106224 97404
rect 106224 97348 106228 97404
rect 106164 97344 106228 97348
rect 4876 96860 4940 96864
rect 4876 96804 4880 96860
rect 4880 96804 4936 96860
rect 4936 96804 4940 96860
rect 4876 96800 4940 96804
rect 4956 96860 5020 96864
rect 4956 96804 4960 96860
rect 4960 96804 5016 96860
rect 5016 96804 5020 96860
rect 4956 96800 5020 96804
rect 5036 96860 5100 96864
rect 5036 96804 5040 96860
rect 5040 96804 5096 96860
rect 5096 96804 5100 96860
rect 5036 96800 5100 96804
rect 5116 96860 5180 96864
rect 5116 96804 5120 96860
rect 5120 96804 5176 96860
rect 5176 96804 5180 96860
rect 5116 96800 5180 96804
rect 106660 96860 106724 96864
rect 106660 96804 106664 96860
rect 106664 96804 106720 96860
rect 106720 96804 106724 96860
rect 106660 96800 106724 96804
rect 106740 96860 106804 96864
rect 106740 96804 106744 96860
rect 106744 96804 106800 96860
rect 106800 96804 106804 96860
rect 106740 96800 106804 96804
rect 106820 96860 106884 96864
rect 106820 96804 106824 96860
rect 106824 96804 106880 96860
rect 106880 96804 106884 96860
rect 106820 96800 106884 96804
rect 106900 96860 106964 96864
rect 106900 96804 106904 96860
rect 106904 96804 106960 96860
rect 106960 96804 106964 96860
rect 106900 96800 106964 96804
rect 4216 96316 4280 96320
rect 4216 96260 4220 96316
rect 4220 96260 4276 96316
rect 4276 96260 4280 96316
rect 4216 96256 4280 96260
rect 4296 96316 4360 96320
rect 4296 96260 4300 96316
rect 4300 96260 4356 96316
rect 4356 96260 4360 96316
rect 4296 96256 4360 96260
rect 4376 96316 4440 96320
rect 4376 96260 4380 96316
rect 4380 96260 4436 96316
rect 4436 96260 4440 96316
rect 4376 96256 4440 96260
rect 4456 96316 4520 96320
rect 4456 96260 4460 96316
rect 4460 96260 4516 96316
rect 4516 96260 4520 96316
rect 4456 96256 4520 96260
rect 105924 96316 105988 96320
rect 105924 96260 105928 96316
rect 105928 96260 105984 96316
rect 105984 96260 105988 96316
rect 105924 96256 105988 96260
rect 106004 96316 106068 96320
rect 106004 96260 106008 96316
rect 106008 96260 106064 96316
rect 106064 96260 106068 96316
rect 106004 96256 106068 96260
rect 106084 96316 106148 96320
rect 106084 96260 106088 96316
rect 106088 96260 106144 96316
rect 106144 96260 106148 96316
rect 106084 96256 106148 96260
rect 106164 96316 106228 96320
rect 106164 96260 106168 96316
rect 106168 96260 106224 96316
rect 106224 96260 106228 96316
rect 106164 96256 106228 96260
rect 4876 95772 4940 95776
rect 4876 95716 4880 95772
rect 4880 95716 4936 95772
rect 4936 95716 4940 95772
rect 4876 95712 4940 95716
rect 4956 95772 5020 95776
rect 4956 95716 4960 95772
rect 4960 95716 5016 95772
rect 5016 95716 5020 95772
rect 4956 95712 5020 95716
rect 5036 95772 5100 95776
rect 5036 95716 5040 95772
rect 5040 95716 5096 95772
rect 5096 95716 5100 95772
rect 5036 95712 5100 95716
rect 5116 95772 5180 95776
rect 5116 95716 5120 95772
rect 5120 95716 5176 95772
rect 5176 95716 5180 95772
rect 5116 95712 5180 95716
rect 106660 95772 106724 95776
rect 106660 95716 106664 95772
rect 106664 95716 106720 95772
rect 106720 95716 106724 95772
rect 106660 95712 106724 95716
rect 106740 95772 106804 95776
rect 106740 95716 106744 95772
rect 106744 95716 106800 95772
rect 106800 95716 106804 95772
rect 106740 95712 106804 95716
rect 106820 95772 106884 95776
rect 106820 95716 106824 95772
rect 106824 95716 106880 95772
rect 106880 95716 106884 95772
rect 106820 95712 106884 95716
rect 106900 95772 106964 95776
rect 106900 95716 106904 95772
rect 106904 95716 106960 95772
rect 106960 95716 106964 95772
rect 106900 95712 106964 95716
rect 4216 95228 4280 95232
rect 4216 95172 4220 95228
rect 4220 95172 4276 95228
rect 4276 95172 4280 95228
rect 4216 95168 4280 95172
rect 4296 95228 4360 95232
rect 4296 95172 4300 95228
rect 4300 95172 4356 95228
rect 4356 95172 4360 95228
rect 4296 95168 4360 95172
rect 4376 95228 4440 95232
rect 4376 95172 4380 95228
rect 4380 95172 4436 95228
rect 4436 95172 4440 95228
rect 4376 95168 4440 95172
rect 4456 95228 4520 95232
rect 4456 95172 4460 95228
rect 4460 95172 4516 95228
rect 4516 95172 4520 95228
rect 4456 95168 4520 95172
rect 105924 95228 105988 95232
rect 105924 95172 105928 95228
rect 105928 95172 105984 95228
rect 105984 95172 105988 95228
rect 105924 95168 105988 95172
rect 106004 95228 106068 95232
rect 106004 95172 106008 95228
rect 106008 95172 106064 95228
rect 106064 95172 106068 95228
rect 106004 95168 106068 95172
rect 106084 95228 106148 95232
rect 106084 95172 106088 95228
rect 106088 95172 106144 95228
rect 106144 95172 106148 95228
rect 106084 95168 106148 95172
rect 106164 95228 106228 95232
rect 106164 95172 106168 95228
rect 106168 95172 106224 95228
rect 106224 95172 106228 95228
rect 106164 95168 106228 95172
rect 4876 94684 4940 94688
rect 4876 94628 4880 94684
rect 4880 94628 4936 94684
rect 4936 94628 4940 94684
rect 4876 94624 4940 94628
rect 4956 94684 5020 94688
rect 4956 94628 4960 94684
rect 4960 94628 5016 94684
rect 5016 94628 5020 94684
rect 4956 94624 5020 94628
rect 5036 94684 5100 94688
rect 5036 94628 5040 94684
rect 5040 94628 5096 94684
rect 5096 94628 5100 94684
rect 5036 94624 5100 94628
rect 5116 94684 5180 94688
rect 5116 94628 5120 94684
rect 5120 94628 5176 94684
rect 5176 94628 5180 94684
rect 5116 94624 5180 94628
rect 106660 94684 106724 94688
rect 106660 94628 106664 94684
rect 106664 94628 106720 94684
rect 106720 94628 106724 94684
rect 106660 94624 106724 94628
rect 106740 94684 106804 94688
rect 106740 94628 106744 94684
rect 106744 94628 106800 94684
rect 106800 94628 106804 94684
rect 106740 94624 106804 94628
rect 106820 94684 106884 94688
rect 106820 94628 106824 94684
rect 106824 94628 106880 94684
rect 106880 94628 106884 94684
rect 106820 94624 106884 94628
rect 106900 94684 106964 94688
rect 106900 94628 106904 94684
rect 106904 94628 106960 94684
rect 106960 94628 106964 94684
rect 106900 94624 106964 94628
rect 4216 94140 4280 94144
rect 4216 94084 4220 94140
rect 4220 94084 4276 94140
rect 4276 94084 4280 94140
rect 4216 94080 4280 94084
rect 4296 94140 4360 94144
rect 4296 94084 4300 94140
rect 4300 94084 4356 94140
rect 4356 94084 4360 94140
rect 4296 94080 4360 94084
rect 4376 94140 4440 94144
rect 4376 94084 4380 94140
rect 4380 94084 4436 94140
rect 4436 94084 4440 94140
rect 4376 94080 4440 94084
rect 4456 94140 4520 94144
rect 4456 94084 4460 94140
rect 4460 94084 4516 94140
rect 4516 94084 4520 94140
rect 4456 94080 4520 94084
rect 105924 94140 105988 94144
rect 105924 94084 105928 94140
rect 105928 94084 105984 94140
rect 105984 94084 105988 94140
rect 105924 94080 105988 94084
rect 106004 94140 106068 94144
rect 106004 94084 106008 94140
rect 106008 94084 106064 94140
rect 106064 94084 106068 94140
rect 106004 94080 106068 94084
rect 106084 94140 106148 94144
rect 106084 94084 106088 94140
rect 106088 94084 106144 94140
rect 106144 94084 106148 94140
rect 106084 94080 106148 94084
rect 106164 94140 106228 94144
rect 106164 94084 106168 94140
rect 106168 94084 106224 94140
rect 106224 94084 106228 94140
rect 106164 94080 106228 94084
rect 4876 93596 4940 93600
rect 4876 93540 4880 93596
rect 4880 93540 4936 93596
rect 4936 93540 4940 93596
rect 4876 93536 4940 93540
rect 4956 93596 5020 93600
rect 4956 93540 4960 93596
rect 4960 93540 5016 93596
rect 5016 93540 5020 93596
rect 4956 93536 5020 93540
rect 5036 93596 5100 93600
rect 5036 93540 5040 93596
rect 5040 93540 5096 93596
rect 5096 93540 5100 93596
rect 5036 93536 5100 93540
rect 5116 93596 5180 93600
rect 5116 93540 5120 93596
rect 5120 93540 5176 93596
rect 5176 93540 5180 93596
rect 5116 93536 5180 93540
rect 106660 93596 106724 93600
rect 106660 93540 106664 93596
rect 106664 93540 106720 93596
rect 106720 93540 106724 93596
rect 106660 93536 106724 93540
rect 106740 93596 106804 93600
rect 106740 93540 106744 93596
rect 106744 93540 106800 93596
rect 106800 93540 106804 93596
rect 106740 93536 106804 93540
rect 106820 93596 106884 93600
rect 106820 93540 106824 93596
rect 106824 93540 106880 93596
rect 106880 93540 106884 93596
rect 106820 93536 106884 93540
rect 106900 93596 106964 93600
rect 106900 93540 106904 93596
rect 106904 93540 106960 93596
rect 106960 93540 106964 93596
rect 106900 93536 106964 93540
rect 102180 93328 102244 93392
rect 4216 93052 4280 93056
rect 4216 92996 4220 93052
rect 4220 92996 4276 93052
rect 4276 92996 4280 93052
rect 4216 92992 4280 92996
rect 4296 93052 4360 93056
rect 4296 92996 4300 93052
rect 4300 92996 4356 93052
rect 4356 92996 4360 93052
rect 4296 92992 4360 92996
rect 4376 93052 4440 93056
rect 4376 92996 4380 93052
rect 4380 92996 4436 93052
rect 4436 92996 4440 93052
rect 4376 92992 4440 92996
rect 4456 93052 4520 93056
rect 4456 92996 4460 93052
rect 4460 92996 4516 93052
rect 4516 92996 4520 93052
rect 4456 92992 4520 92996
rect 105924 93052 105988 93056
rect 105924 92996 105928 93052
rect 105928 92996 105984 93052
rect 105984 92996 105988 93052
rect 105924 92992 105988 92996
rect 106004 93052 106068 93056
rect 106004 92996 106008 93052
rect 106008 92996 106064 93052
rect 106064 92996 106068 93052
rect 106004 92992 106068 92996
rect 106084 93052 106148 93056
rect 106084 92996 106088 93052
rect 106088 92996 106144 93052
rect 106144 92996 106148 93052
rect 106084 92992 106148 92996
rect 106164 93052 106228 93056
rect 106164 92996 106168 93052
rect 106168 92996 106224 93052
rect 106224 92996 106228 93052
rect 106164 92992 106228 92996
rect 4876 92508 4940 92512
rect 4876 92452 4880 92508
rect 4880 92452 4936 92508
rect 4936 92452 4940 92508
rect 4876 92448 4940 92452
rect 4956 92508 5020 92512
rect 4956 92452 4960 92508
rect 4960 92452 5016 92508
rect 5016 92452 5020 92508
rect 4956 92448 5020 92452
rect 5036 92508 5100 92512
rect 5036 92452 5040 92508
rect 5040 92452 5096 92508
rect 5096 92452 5100 92508
rect 5036 92448 5100 92452
rect 5116 92508 5180 92512
rect 5116 92452 5120 92508
rect 5120 92452 5176 92508
rect 5176 92452 5180 92508
rect 5116 92448 5180 92452
rect 106660 92508 106724 92512
rect 106660 92452 106664 92508
rect 106664 92452 106720 92508
rect 106720 92452 106724 92508
rect 106660 92448 106724 92452
rect 106740 92508 106804 92512
rect 106740 92452 106744 92508
rect 106744 92452 106800 92508
rect 106800 92452 106804 92508
rect 106740 92448 106804 92452
rect 106820 92508 106884 92512
rect 106820 92452 106824 92508
rect 106824 92452 106880 92508
rect 106880 92452 106884 92508
rect 106820 92448 106884 92452
rect 106900 92508 106964 92512
rect 106900 92452 106904 92508
rect 106904 92452 106960 92508
rect 106960 92452 106964 92508
rect 106900 92448 106964 92452
rect 4216 91964 4280 91968
rect 4216 91908 4220 91964
rect 4220 91908 4276 91964
rect 4276 91908 4280 91964
rect 4216 91904 4280 91908
rect 4296 91964 4360 91968
rect 4296 91908 4300 91964
rect 4300 91908 4356 91964
rect 4356 91908 4360 91964
rect 4296 91904 4360 91908
rect 4376 91964 4440 91968
rect 4376 91908 4380 91964
rect 4380 91908 4436 91964
rect 4436 91908 4440 91964
rect 4376 91904 4440 91908
rect 4456 91964 4520 91968
rect 4456 91908 4460 91964
rect 4460 91908 4516 91964
rect 4516 91908 4520 91964
rect 4456 91904 4520 91908
rect 105924 91964 105988 91968
rect 105924 91908 105928 91964
rect 105928 91908 105984 91964
rect 105984 91908 105988 91964
rect 105924 91904 105988 91908
rect 106004 91964 106068 91968
rect 106004 91908 106008 91964
rect 106008 91908 106064 91964
rect 106064 91908 106068 91964
rect 106004 91904 106068 91908
rect 106084 91964 106148 91968
rect 106084 91908 106088 91964
rect 106088 91908 106144 91964
rect 106144 91908 106148 91964
rect 106084 91904 106148 91908
rect 106164 91964 106228 91968
rect 106164 91908 106168 91964
rect 106168 91908 106224 91964
rect 106224 91908 106228 91964
rect 106164 91904 106228 91908
rect 4876 91420 4940 91424
rect 4876 91364 4880 91420
rect 4880 91364 4936 91420
rect 4936 91364 4940 91420
rect 4876 91360 4940 91364
rect 4956 91420 5020 91424
rect 4956 91364 4960 91420
rect 4960 91364 5016 91420
rect 5016 91364 5020 91420
rect 4956 91360 5020 91364
rect 5036 91420 5100 91424
rect 5036 91364 5040 91420
rect 5040 91364 5096 91420
rect 5096 91364 5100 91420
rect 5036 91360 5100 91364
rect 5116 91420 5180 91424
rect 5116 91364 5120 91420
rect 5120 91364 5176 91420
rect 5176 91364 5180 91420
rect 5116 91360 5180 91364
rect 106660 91420 106724 91424
rect 106660 91364 106664 91420
rect 106664 91364 106720 91420
rect 106720 91364 106724 91420
rect 106660 91360 106724 91364
rect 106740 91420 106804 91424
rect 106740 91364 106744 91420
rect 106744 91364 106800 91420
rect 106800 91364 106804 91420
rect 106740 91360 106804 91364
rect 106820 91420 106884 91424
rect 106820 91364 106824 91420
rect 106824 91364 106880 91420
rect 106880 91364 106884 91420
rect 106820 91360 106884 91364
rect 106900 91420 106964 91424
rect 106900 91364 106904 91420
rect 106904 91364 106960 91420
rect 106960 91364 106964 91420
rect 106900 91360 106964 91364
rect 4216 90876 4280 90880
rect 4216 90820 4220 90876
rect 4220 90820 4276 90876
rect 4276 90820 4280 90876
rect 4216 90816 4280 90820
rect 4296 90876 4360 90880
rect 4296 90820 4300 90876
rect 4300 90820 4356 90876
rect 4356 90820 4360 90876
rect 4296 90816 4360 90820
rect 4376 90876 4440 90880
rect 4376 90820 4380 90876
rect 4380 90820 4436 90876
rect 4436 90820 4440 90876
rect 4376 90816 4440 90820
rect 4456 90876 4520 90880
rect 4456 90820 4460 90876
rect 4460 90820 4516 90876
rect 4516 90820 4520 90876
rect 4456 90816 4520 90820
rect 105924 90876 105988 90880
rect 105924 90820 105928 90876
rect 105928 90820 105984 90876
rect 105984 90820 105988 90876
rect 105924 90816 105988 90820
rect 106004 90876 106068 90880
rect 106004 90820 106008 90876
rect 106008 90820 106064 90876
rect 106064 90820 106068 90876
rect 106004 90816 106068 90820
rect 106084 90876 106148 90880
rect 106084 90820 106088 90876
rect 106088 90820 106144 90876
rect 106144 90820 106148 90876
rect 106084 90816 106148 90820
rect 106164 90876 106228 90880
rect 106164 90820 106168 90876
rect 106168 90820 106224 90876
rect 106224 90820 106228 90876
rect 106164 90816 106228 90820
rect 4876 90332 4940 90336
rect 4876 90276 4880 90332
rect 4880 90276 4936 90332
rect 4936 90276 4940 90332
rect 4876 90272 4940 90276
rect 4956 90332 5020 90336
rect 4956 90276 4960 90332
rect 4960 90276 5016 90332
rect 5016 90276 5020 90332
rect 4956 90272 5020 90276
rect 5036 90332 5100 90336
rect 5036 90276 5040 90332
rect 5040 90276 5096 90332
rect 5096 90276 5100 90332
rect 5036 90272 5100 90276
rect 5116 90332 5180 90336
rect 5116 90276 5120 90332
rect 5120 90276 5176 90332
rect 5176 90276 5180 90332
rect 5116 90272 5180 90276
rect 106660 90332 106724 90336
rect 106660 90276 106664 90332
rect 106664 90276 106720 90332
rect 106720 90276 106724 90332
rect 106660 90272 106724 90276
rect 106740 90332 106804 90336
rect 106740 90276 106744 90332
rect 106744 90276 106800 90332
rect 106800 90276 106804 90332
rect 106740 90272 106804 90276
rect 106820 90332 106884 90336
rect 106820 90276 106824 90332
rect 106824 90276 106880 90332
rect 106880 90276 106884 90332
rect 106820 90272 106884 90276
rect 106900 90332 106964 90336
rect 106900 90276 106904 90332
rect 106904 90276 106960 90332
rect 106960 90276 106964 90332
rect 106900 90272 106964 90276
rect 4216 89788 4280 89792
rect 4216 89732 4220 89788
rect 4220 89732 4276 89788
rect 4276 89732 4280 89788
rect 4216 89728 4280 89732
rect 4296 89788 4360 89792
rect 4296 89732 4300 89788
rect 4300 89732 4356 89788
rect 4356 89732 4360 89788
rect 4296 89728 4360 89732
rect 4376 89788 4440 89792
rect 4376 89732 4380 89788
rect 4380 89732 4436 89788
rect 4436 89732 4440 89788
rect 4376 89728 4440 89732
rect 4456 89788 4520 89792
rect 4456 89732 4460 89788
rect 4460 89732 4516 89788
rect 4516 89732 4520 89788
rect 4456 89728 4520 89732
rect 105924 89788 105988 89792
rect 105924 89732 105928 89788
rect 105928 89732 105984 89788
rect 105984 89732 105988 89788
rect 105924 89728 105988 89732
rect 106004 89788 106068 89792
rect 106004 89732 106008 89788
rect 106008 89732 106064 89788
rect 106064 89732 106068 89788
rect 106004 89728 106068 89732
rect 106084 89788 106148 89792
rect 106084 89732 106088 89788
rect 106088 89732 106144 89788
rect 106144 89732 106148 89788
rect 106084 89728 106148 89732
rect 106164 89788 106228 89792
rect 106164 89732 106168 89788
rect 106168 89732 106224 89788
rect 106224 89732 106228 89788
rect 106164 89728 106228 89732
rect 4876 89244 4940 89248
rect 4876 89188 4880 89244
rect 4880 89188 4936 89244
rect 4936 89188 4940 89244
rect 4876 89184 4940 89188
rect 4956 89244 5020 89248
rect 4956 89188 4960 89244
rect 4960 89188 5016 89244
rect 5016 89188 5020 89244
rect 4956 89184 5020 89188
rect 5036 89244 5100 89248
rect 5036 89188 5040 89244
rect 5040 89188 5096 89244
rect 5096 89188 5100 89244
rect 5036 89184 5100 89188
rect 5116 89244 5180 89248
rect 5116 89188 5120 89244
rect 5120 89188 5176 89244
rect 5176 89188 5180 89244
rect 5116 89184 5180 89188
rect 106660 89244 106724 89248
rect 106660 89188 106664 89244
rect 106664 89188 106720 89244
rect 106720 89188 106724 89244
rect 106660 89184 106724 89188
rect 106740 89244 106804 89248
rect 106740 89188 106744 89244
rect 106744 89188 106800 89244
rect 106800 89188 106804 89244
rect 106740 89184 106804 89188
rect 106820 89244 106884 89248
rect 106820 89188 106824 89244
rect 106824 89188 106880 89244
rect 106880 89188 106884 89244
rect 106820 89184 106884 89188
rect 106900 89244 106964 89248
rect 106900 89188 106904 89244
rect 106904 89188 106960 89244
rect 106960 89188 106964 89244
rect 106900 89184 106964 89188
rect 4216 88700 4280 88704
rect 4216 88644 4220 88700
rect 4220 88644 4276 88700
rect 4276 88644 4280 88700
rect 4216 88640 4280 88644
rect 4296 88700 4360 88704
rect 4296 88644 4300 88700
rect 4300 88644 4356 88700
rect 4356 88644 4360 88700
rect 4296 88640 4360 88644
rect 4376 88700 4440 88704
rect 4376 88644 4380 88700
rect 4380 88644 4436 88700
rect 4436 88644 4440 88700
rect 4376 88640 4440 88644
rect 4456 88700 4520 88704
rect 4456 88644 4460 88700
rect 4460 88644 4516 88700
rect 4516 88644 4520 88700
rect 4456 88640 4520 88644
rect 105924 88700 105988 88704
rect 105924 88644 105928 88700
rect 105928 88644 105984 88700
rect 105984 88644 105988 88700
rect 105924 88640 105988 88644
rect 106004 88700 106068 88704
rect 106004 88644 106008 88700
rect 106008 88644 106064 88700
rect 106064 88644 106068 88700
rect 106004 88640 106068 88644
rect 106084 88700 106148 88704
rect 106084 88644 106088 88700
rect 106088 88644 106144 88700
rect 106144 88644 106148 88700
rect 106084 88640 106148 88644
rect 106164 88700 106228 88704
rect 106164 88644 106168 88700
rect 106168 88644 106224 88700
rect 106224 88644 106228 88700
rect 106164 88640 106228 88644
rect 4876 88156 4940 88160
rect 4876 88100 4880 88156
rect 4880 88100 4936 88156
rect 4936 88100 4940 88156
rect 4876 88096 4940 88100
rect 4956 88156 5020 88160
rect 4956 88100 4960 88156
rect 4960 88100 5016 88156
rect 5016 88100 5020 88156
rect 4956 88096 5020 88100
rect 5036 88156 5100 88160
rect 5036 88100 5040 88156
rect 5040 88100 5096 88156
rect 5096 88100 5100 88156
rect 5036 88096 5100 88100
rect 5116 88156 5180 88160
rect 5116 88100 5120 88156
rect 5120 88100 5176 88156
rect 5176 88100 5180 88156
rect 5116 88096 5180 88100
rect 106660 88156 106724 88160
rect 106660 88100 106664 88156
rect 106664 88100 106720 88156
rect 106720 88100 106724 88156
rect 106660 88096 106724 88100
rect 106740 88156 106804 88160
rect 106740 88100 106744 88156
rect 106744 88100 106800 88156
rect 106800 88100 106804 88156
rect 106740 88096 106804 88100
rect 106820 88156 106884 88160
rect 106820 88100 106824 88156
rect 106824 88100 106880 88156
rect 106880 88100 106884 88156
rect 106820 88096 106884 88100
rect 106900 88156 106964 88160
rect 106900 88100 106904 88156
rect 106904 88100 106960 88156
rect 106960 88100 106964 88156
rect 106900 88096 106964 88100
rect 4216 87612 4280 87616
rect 4216 87556 4220 87612
rect 4220 87556 4276 87612
rect 4276 87556 4280 87612
rect 4216 87552 4280 87556
rect 4296 87612 4360 87616
rect 4296 87556 4300 87612
rect 4300 87556 4356 87612
rect 4356 87556 4360 87612
rect 4296 87552 4360 87556
rect 4376 87612 4440 87616
rect 4376 87556 4380 87612
rect 4380 87556 4436 87612
rect 4436 87556 4440 87612
rect 4376 87552 4440 87556
rect 4456 87612 4520 87616
rect 4456 87556 4460 87612
rect 4460 87556 4516 87612
rect 4516 87556 4520 87612
rect 4456 87552 4520 87556
rect 105924 87612 105988 87616
rect 105924 87556 105928 87612
rect 105928 87556 105984 87612
rect 105984 87556 105988 87612
rect 105924 87552 105988 87556
rect 106004 87612 106068 87616
rect 106004 87556 106008 87612
rect 106008 87556 106064 87612
rect 106064 87556 106068 87612
rect 106004 87552 106068 87556
rect 106084 87612 106148 87616
rect 106084 87556 106088 87612
rect 106088 87556 106144 87612
rect 106144 87556 106148 87612
rect 106084 87552 106148 87556
rect 106164 87612 106228 87616
rect 106164 87556 106168 87612
rect 106168 87556 106224 87612
rect 106224 87556 106228 87612
rect 106164 87552 106228 87556
rect 4876 87068 4940 87072
rect 4876 87012 4880 87068
rect 4880 87012 4936 87068
rect 4936 87012 4940 87068
rect 4876 87008 4940 87012
rect 4956 87068 5020 87072
rect 4956 87012 4960 87068
rect 4960 87012 5016 87068
rect 5016 87012 5020 87068
rect 4956 87008 5020 87012
rect 5036 87068 5100 87072
rect 5036 87012 5040 87068
rect 5040 87012 5096 87068
rect 5096 87012 5100 87068
rect 5036 87008 5100 87012
rect 5116 87068 5180 87072
rect 5116 87012 5120 87068
rect 5120 87012 5176 87068
rect 5176 87012 5180 87068
rect 5116 87008 5180 87012
rect 106660 87068 106724 87072
rect 106660 87012 106664 87068
rect 106664 87012 106720 87068
rect 106720 87012 106724 87068
rect 106660 87008 106724 87012
rect 106740 87068 106804 87072
rect 106740 87012 106744 87068
rect 106744 87012 106800 87068
rect 106800 87012 106804 87068
rect 106740 87008 106804 87012
rect 106820 87068 106884 87072
rect 106820 87012 106824 87068
rect 106824 87012 106880 87068
rect 106880 87012 106884 87068
rect 106820 87008 106884 87012
rect 106900 87068 106964 87072
rect 106900 87012 106904 87068
rect 106904 87012 106960 87068
rect 106960 87012 106964 87068
rect 106900 87008 106964 87012
rect 4216 86524 4280 86528
rect 4216 86468 4220 86524
rect 4220 86468 4276 86524
rect 4276 86468 4280 86524
rect 4216 86464 4280 86468
rect 4296 86524 4360 86528
rect 4296 86468 4300 86524
rect 4300 86468 4356 86524
rect 4356 86468 4360 86524
rect 4296 86464 4360 86468
rect 4376 86524 4440 86528
rect 4376 86468 4380 86524
rect 4380 86468 4436 86524
rect 4436 86468 4440 86524
rect 4376 86464 4440 86468
rect 4456 86524 4520 86528
rect 4456 86468 4460 86524
rect 4460 86468 4516 86524
rect 4516 86468 4520 86524
rect 4456 86464 4520 86468
rect 105924 86524 105988 86528
rect 105924 86468 105928 86524
rect 105928 86468 105984 86524
rect 105984 86468 105988 86524
rect 105924 86464 105988 86468
rect 106004 86524 106068 86528
rect 106004 86468 106008 86524
rect 106008 86468 106064 86524
rect 106064 86468 106068 86524
rect 106004 86464 106068 86468
rect 106084 86524 106148 86528
rect 106084 86468 106088 86524
rect 106088 86468 106144 86524
rect 106144 86468 106148 86524
rect 106084 86464 106148 86468
rect 106164 86524 106228 86528
rect 106164 86468 106168 86524
rect 106168 86468 106224 86524
rect 106224 86468 106228 86524
rect 106164 86464 106228 86468
rect 4876 85980 4940 85984
rect 4876 85924 4880 85980
rect 4880 85924 4936 85980
rect 4936 85924 4940 85980
rect 4876 85920 4940 85924
rect 4956 85980 5020 85984
rect 4956 85924 4960 85980
rect 4960 85924 5016 85980
rect 5016 85924 5020 85980
rect 4956 85920 5020 85924
rect 5036 85980 5100 85984
rect 5036 85924 5040 85980
rect 5040 85924 5096 85980
rect 5096 85924 5100 85980
rect 5036 85920 5100 85924
rect 5116 85980 5180 85984
rect 5116 85924 5120 85980
rect 5120 85924 5176 85980
rect 5176 85924 5180 85980
rect 5116 85920 5180 85924
rect 106660 85980 106724 85984
rect 106660 85924 106664 85980
rect 106664 85924 106720 85980
rect 106720 85924 106724 85980
rect 106660 85920 106724 85924
rect 106740 85980 106804 85984
rect 106740 85924 106744 85980
rect 106744 85924 106800 85980
rect 106800 85924 106804 85980
rect 106740 85920 106804 85924
rect 106820 85980 106884 85984
rect 106820 85924 106824 85980
rect 106824 85924 106880 85980
rect 106880 85924 106884 85980
rect 106820 85920 106884 85924
rect 106900 85980 106964 85984
rect 106900 85924 106904 85980
rect 106904 85924 106960 85980
rect 106960 85924 106964 85980
rect 106900 85920 106964 85924
rect 4216 85436 4280 85440
rect 4216 85380 4220 85436
rect 4220 85380 4276 85436
rect 4276 85380 4280 85436
rect 4216 85376 4280 85380
rect 4296 85436 4360 85440
rect 4296 85380 4300 85436
rect 4300 85380 4356 85436
rect 4356 85380 4360 85436
rect 4296 85376 4360 85380
rect 4376 85436 4440 85440
rect 4376 85380 4380 85436
rect 4380 85380 4436 85436
rect 4436 85380 4440 85436
rect 4376 85376 4440 85380
rect 4456 85436 4520 85440
rect 4456 85380 4460 85436
rect 4460 85380 4516 85436
rect 4516 85380 4520 85436
rect 4456 85376 4520 85380
rect 105924 85436 105988 85440
rect 105924 85380 105928 85436
rect 105928 85380 105984 85436
rect 105984 85380 105988 85436
rect 105924 85376 105988 85380
rect 106004 85436 106068 85440
rect 106004 85380 106008 85436
rect 106008 85380 106064 85436
rect 106064 85380 106068 85436
rect 106004 85376 106068 85380
rect 106084 85436 106148 85440
rect 106084 85380 106088 85436
rect 106088 85380 106144 85436
rect 106144 85380 106148 85436
rect 106084 85376 106148 85380
rect 106164 85436 106228 85440
rect 106164 85380 106168 85436
rect 106168 85380 106224 85436
rect 106224 85380 106228 85436
rect 106164 85376 106228 85380
rect 4876 84892 4940 84896
rect 4876 84836 4880 84892
rect 4880 84836 4936 84892
rect 4936 84836 4940 84892
rect 4876 84832 4940 84836
rect 4956 84892 5020 84896
rect 4956 84836 4960 84892
rect 4960 84836 5016 84892
rect 5016 84836 5020 84892
rect 4956 84832 5020 84836
rect 5036 84892 5100 84896
rect 5036 84836 5040 84892
rect 5040 84836 5096 84892
rect 5096 84836 5100 84892
rect 5036 84832 5100 84836
rect 5116 84892 5180 84896
rect 5116 84836 5120 84892
rect 5120 84836 5176 84892
rect 5176 84836 5180 84892
rect 5116 84832 5180 84836
rect 106660 84892 106724 84896
rect 106660 84836 106664 84892
rect 106664 84836 106720 84892
rect 106720 84836 106724 84892
rect 106660 84832 106724 84836
rect 106740 84892 106804 84896
rect 106740 84836 106744 84892
rect 106744 84836 106800 84892
rect 106800 84836 106804 84892
rect 106740 84832 106804 84836
rect 106820 84892 106884 84896
rect 106820 84836 106824 84892
rect 106824 84836 106880 84892
rect 106880 84836 106884 84892
rect 106820 84832 106884 84836
rect 106900 84892 106964 84896
rect 106900 84836 106904 84892
rect 106904 84836 106960 84892
rect 106960 84836 106964 84892
rect 106900 84832 106964 84836
rect 4216 84348 4280 84352
rect 4216 84292 4220 84348
rect 4220 84292 4276 84348
rect 4276 84292 4280 84348
rect 4216 84288 4280 84292
rect 4296 84348 4360 84352
rect 4296 84292 4300 84348
rect 4300 84292 4356 84348
rect 4356 84292 4360 84348
rect 4296 84288 4360 84292
rect 4376 84348 4440 84352
rect 4376 84292 4380 84348
rect 4380 84292 4436 84348
rect 4436 84292 4440 84348
rect 4376 84288 4440 84292
rect 4456 84348 4520 84352
rect 4456 84292 4460 84348
rect 4460 84292 4516 84348
rect 4516 84292 4520 84348
rect 4456 84288 4520 84292
rect 105924 84348 105988 84352
rect 105924 84292 105928 84348
rect 105928 84292 105984 84348
rect 105984 84292 105988 84348
rect 105924 84288 105988 84292
rect 106004 84348 106068 84352
rect 106004 84292 106008 84348
rect 106008 84292 106064 84348
rect 106064 84292 106068 84348
rect 106004 84288 106068 84292
rect 106084 84348 106148 84352
rect 106084 84292 106088 84348
rect 106088 84292 106144 84348
rect 106144 84292 106148 84348
rect 106084 84288 106148 84292
rect 106164 84348 106228 84352
rect 106164 84292 106168 84348
rect 106168 84292 106224 84348
rect 106224 84292 106228 84348
rect 106164 84288 106228 84292
rect 4876 83804 4940 83808
rect 4876 83748 4880 83804
rect 4880 83748 4936 83804
rect 4936 83748 4940 83804
rect 4876 83744 4940 83748
rect 4956 83804 5020 83808
rect 4956 83748 4960 83804
rect 4960 83748 5016 83804
rect 5016 83748 5020 83804
rect 4956 83744 5020 83748
rect 5036 83804 5100 83808
rect 5036 83748 5040 83804
rect 5040 83748 5096 83804
rect 5096 83748 5100 83804
rect 5036 83744 5100 83748
rect 5116 83804 5180 83808
rect 5116 83748 5120 83804
rect 5120 83748 5176 83804
rect 5176 83748 5180 83804
rect 5116 83744 5180 83748
rect 106660 83804 106724 83808
rect 106660 83748 106664 83804
rect 106664 83748 106720 83804
rect 106720 83748 106724 83804
rect 106660 83744 106724 83748
rect 106740 83804 106804 83808
rect 106740 83748 106744 83804
rect 106744 83748 106800 83804
rect 106800 83748 106804 83804
rect 106740 83744 106804 83748
rect 106820 83804 106884 83808
rect 106820 83748 106824 83804
rect 106824 83748 106880 83804
rect 106880 83748 106884 83804
rect 106820 83744 106884 83748
rect 106900 83804 106964 83808
rect 106900 83748 106904 83804
rect 106904 83748 106960 83804
rect 106960 83748 106964 83804
rect 106900 83744 106964 83748
rect 4216 83260 4280 83264
rect 4216 83204 4220 83260
rect 4220 83204 4276 83260
rect 4276 83204 4280 83260
rect 4216 83200 4280 83204
rect 4296 83260 4360 83264
rect 4296 83204 4300 83260
rect 4300 83204 4356 83260
rect 4356 83204 4360 83260
rect 4296 83200 4360 83204
rect 4376 83260 4440 83264
rect 4376 83204 4380 83260
rect 4380 83204 4436 83260
rect 4436 83204 4440 83260
rect 4376 83200 4440 83204
rect 4456 83260 4520 83264
rect 4456 83204 4460 83260
rect 4460 83204 4516 83260
rect 4516 83204 4520 83260
rect 4456 83200 4520 83204
rect 105924 83260 105988 83264
rect 105924 83204 105928 83260
rect 105928 83204 105984 83260
rect 105984 83204 105988 83260
rect 105924 83200 105988 83204
rect 106004 83260 106068 83264
rect 106004 83204 106008 83260
rect 106008 83204 106064 83260
rect 106064 83204 106068 83260
rect 106004 83200 106068 83204
rect 106084 83260 106148 83264
rect 106084 83204 106088 83260
rect 106088 83204 106144 83260
rect 106144 83204 106148 83260
rect 106084 83200 106148 83204
rect 106164 83260 106228 83264
rect 106164 83204 106168 83260
rect 106168 83204 106224 83260
rect 106224 83204 106228 83260
rect 106164 83200 106228 83204
rect 4876 82716 4940 82720
rect 4876 82660 4880 82716
rect 4880 82660 4936 82716
rect 4936 82660 4940 82716
rect 4876 82656 4940 82660
rect 4956 82716 5020 82720
rect 4956 82660 4960 82716
rect 4960 82660 5016 82716
rect 5016 82660 5020 82716
rect 4956 82656 5020 82660
rect 5036 82716 5100 82720
rect 5036 82660 5040 82716
rect 5040 82660 5096 82716
rect 5096 82660 5100 82716
rect 5036 82656 5100 82660
rect 5116 82716 5180 82720
rect 5116 82660 5120 82716
rect 5120 82660 5176 82716
rect 5176 82660 5180 82716
rect 5116 82656 5180 82660
rect 106660 82716 106724 82720
rect 106660 82660 106664 82716
rect 106664 82660 106720 82716
rect 106720 82660 106724 82716
rect 106660 82656 106724 82660
rect 106740 82716 106804 82720
rect 106740 82660 106744 82716
rect 106744 82660 106800 82716
rect 106800 82660 106804 82716
rect 106740 82656 106804 82660
rect 106820 82716 106884 82720
rect 106820 82660 106824 82716
rect 106824 82660 106880 82716
rect 106880 82660 106884 82716
rect 106820 82656 106884 82660
rect 106900 82716 106964 82720
rect 106900 82660 106904 82716
rect 106904 82660 106960 82716
rect 106960 82660 106964 82716
rect 106900 82656 106964 82660
rect 4216 82172 4280 82176
rect 4216 82116 4220 82172
rect 4220 82116 4276 82172
rect 4276 82116 4280 82172
rect 4216 82112 4280 82116
rect 4296 82172 4360 82176
rect 4296 82116 4300 82172
rect 4300 82116 4356 82172
rect 4356 82116 4360 82172
rect 4296 82112 4360 82116
rect 4376 82172 4440 82176
rect 4376 82116 4380 82172
rect 4380 82116 4436 82172
rect 4436 82116 4440 82172
rect 4376 82112 4440 82116
rect 4456 82172 4520 82176
rect 4456 82116 4460 82172
rect 4460 82116 4516 82172
rect 4516 82116 4520 82172
rect 4456 82112 4520 82116
rect 105924 82172 105988 82176
rect 105924 82116 105928 82172
rect 105928 82116 105984 82172
rect 105984 82116 105988 82172
rect 105924 82112 105988 82116
rect 106004 82172 106068 82176
rect 106004 82116 106008 82172
rect 106008 82116 106064 82172
rect 106064 82116 106068 82172
rect 106004 82112 106068 82116
rect 106084 82172 106148 82176
rect 106084 82116 106088 82172
rect 106088 82116 106144 82172
rect 106144 82116 106148 82172
rect 106084 82112 106148 82116
rect 106164 82172 106228 82176
rect 106164 82116 106168 82172
rect 106168 82116 106224 82172
rect 106224 82116 106228 82172
rect 106164 82112 106228 82116
rect 4876 81628 4940 81632
rect 4876 81572 4880 81628
rect 4880 81572 4936 81628
rect 4936 81572 4940 81628
rect 4876 81568 4940 81572
rect 4956 81628 5020 81632
rect 4956 81572 4960 81628
rect 4960 81572 5016 81628
rect 5016 81572 5020 81628
rect 4956 81568 5020 81572
rect 5036 81628 5100 81632
rect 5036 81572 5040 81628
rect 5040 81572 5096 81628
rect 5096 81572 5100 81628
rect 5036 81568 5100 81572
rect 5116 81628 5180 81632
rect 5116 81572 5120 81628
rect 5120 81572 5176 81628
rect 5176 81572 5180 81628
rect 5116 81568 5180 81572
rect 106660 81628 106724 81632
rect 106660 81572 106664 81628
rect 106664 81572 106720 81628
rect 106720 81572 106724 81628
rect 106660 81568 106724 81572
rect 106740 81628 106804 81632
rect 106740 81572 106744 81628
rect 106744 81572 106800 81628
rect 106800 81572 106804 81628
rect 106740 81568 106804 81572
rect 106820 81628 106884 81632
rect 106820 81572 106824 81628
rect 106824 81572 106880 81628
rect 106880 81572 106884 81628
rect 106820 81568 106884 81572
rect 106900 81628 106964 81632
rect 106900 81572 106904 81628
rect 106904 81572 106960 81628
rect 106960 81572 106964 81628
rect 106900 81568 106964 81572
rect 4216 81084 4280 81088
rect 4216 81028 4220 81084
rect 4220 81028 4276 81084
rect 4276 81028 4280 81084
rect 4216 81024 4280 81028
rect 4296 81084 4360 81088
rect 4296 81028 4300 81084
rect 4300 81028 4356 81084
rect 4356 81028 4360 81084
rect 4296 81024 4360 81028
rect 4376 81084 4440 81088
rect 4376 81028 4380 81084
rect 4380 81028 4436 81084
rect 4436 81028 4440 81084
rect 4376 81024 4440 81028
rect 4456 81084 4520 81088
rect 4456 81028 4460 81084
rect 4460 81028 4516 81084
rect 4516 81028 4520 81084
rect 4456 81024 4520 81028
rect 105924 81084 105988 81088
rect 105924 81028 105928 81084
rect 105928 81028 105984 81084
rect 105984 81028 105988 81084
rect 105924 81024 105988 81028
rect 106004 81084 106068 81088
rect 106004 81028 106008 81084
rect 106008 81028 106064 81084
rect 106064 81028 106068 81084
rect 106004 81024 106068 81028
rect 106084 81084 106148 81088
rect 106084 81028 106088 81084
rect 106088 81028 106144 81084
rect 106144 81028 106148 81084
rect 106084 81024 106148 81028
rect 106164 81084 106228 81088
rect 106164 81028 106168 81084
rect 106168 81028 106224 81084
rect 106224 81028 106228 81084
rect 106164 81024 106228 81028
rect 4876 80540 4940 80544
rect 4876 80484 4880 80540
rect 4880 80484 4936 80540
rect 4936 80484 4940 80540
rect 4876 80480 4940 80484
rect 4956 80540 5020 80544
rect 4956 80484 4960 80540
rect 4960 80484 5016 80540
rect 5016 80484 5020 80540
rect 4956 80480 5020 80484
rect 5036 80540 5100 80544
rect 5036 80484 5040 80540
rect 5040 80484 5096 80540
rect 5096 80484 5100 80540
rect 5036 80480 5100 80484
rect 5116 80540 5180 80544
rect 5116 80484 5120 80540
rect 5120 80484 5176 80540
rect 5176 80484 5180 80540
rect 5116 80480 5180 80484
rect 106660 80540 106724 80544
rect 106660 80484 106664 80540
rect 106664 80484 106720 80540
rect 106720 80484 106724 80540
rect 106660 80480 106724 80484
rect 106740 80540 106804 80544
rect 106740 80484 106744 80540
rect 106744 80484 106800 80540
rect 106800 80484 106804 80540
rect 106740 80480 106804 80484
rect 106820 80540 106884 80544
rect 106820 80484 106824 80540
rect 106824 80484 106880 80540
rect 106880 80484 106884 80540
rect 106820 80480 106884 80484
rect 106900 80540 106964 80544
rect 106900 80484 106904 80540
rect 106904 80484 106960 80540
rect 106960 80484 106964 80540
rect 106900 80480 106964 80484
rect 4216 79996 4280 80000
rect 4216 79940 4220 79996
rect 4220 79940 4276 79996
rect 4276 79940 4280 79996
rect 4216 79936 4280 79940
rect 4296 79996 4360 80000
rect 4296 79940 4300 79996
rect 4300 79940 4356 79996
rect 4356 79940 4360 79996
rect 4296 79936 4360 79940
rect 4376 79996 4440 80000
rect 4376 79940 4380 79996
rect 4380 79940 4436 79996
rect 4436 79940 4440 79996
rect 4376 79936 4440 79940
rect 4456 79996 4520 80000
rect 4456 79940 4460 79996
rect 4460 79940 4516 79996
rect 4516 79940 4520 79996
rect 4456 79936 4520 79940
rect 105924 79996 105988 80000
rect 105924 79940 105928 79996
rect 105928 79940 105984 79996
rect 105984 79940 105988 79996
rect 105924 79936 105988 79940
rect 106004 79996 106068 80000
rect 106004 79940 106008 79996
rect 106008 79940 106064 79996
rect 106064 79940 106068 79996
rect 106004 79936 106068 79940
rect 106084 79996 106148 80000
rect 106084 79940 106088 79996
rect 106088 79940 106144 79996
rect 106144 79940 106148 79996
rect 106084 79936 106148 79940
rect 106164 79996 106228 80000
rect 106164 79940 106168 79996
rect 106168 79940 106224 79996
rect 106224 79940 106228 79996
rect 106164 79936 106228 79940
rect 16068 79928 16132 79932
rect 16068 79872 16118 79928
rect 16118 79872 16132 79928
rect 16068 79868 16132 79872
rect 23438 79928 23502 79932
rect 23438 79872 23478 79928
rect 23478 79872 23502 79928
rect 23438 79868 23502 79872
rect 36286 79928 36350 79932
rect 36286 79872 36322 79928
rect 36322 79872 36350 79928
rect 36286 79868 36350 79872
rect 39790 79928 39854 79932
rect 39790 79872 39818 79928
rect 39818 79872 39854 79928
rect 39790 79868 39854 79872
rect 40958 79928 41022 79932
rect 40958 79872 41014 79928
rect 41014 79872 41022 79928
rect 40958 79868 41022 79872
rect 43294 79928 43358 79932
rect 43294 79872 43314 79928
rect 43314 79872 43358 79928
rect 43294 79868 43358 79872
rect 32782 79732 32846 79796
rect 38622 79792 38686 79796
rect 38622 79736 38658 79792
rect 38658 79736 38686 79792
rect 38622 79732 38686 79736
rect 30446 79656 30510 79660
rect 30446 79600 30470 79656
rect 30470 79600 30510 79656
rect 30446 79596 30510 79600
rect 31616 79656 31680 79660
rect 31616 79600 31666 79656
rect 31666 79600 31680 79656
rect 31616 79596 31680 79600
rect 37454 79656 37518 79660
rect 37454 79600 37462 79656
rect 37462 79600 37518 79656
rect 37454 79596 37518 79600
rect 24624 79520 24688 79524
rect 24624 79464 24674 79520
rect 24674 79464 24688 79520
rect 24624 79460 24688 79464
rect 25774 79460 25838 79524
rect 26942 79520 27006 79524
rect 26942 79464 26974 79520
rect 26974 79464 27006 79520
rect 26942 79460 27006 79464
rect 28120 79520 28184 79524
rect 28120 79464 28170 79520
rect 28170 79464 28184 79520
rect 28120 79460 28184 79464
rect 29278 79460 29342 79524
rect 33950 79520 34014 79524
rect 33950 79464 33966 79520
rect 33966 79464 34014 79520
rect 33950 79460 34014 79464
rect 35118 79460 35182 79524
rect 42126 79520 42190 79524
rect 42126 79464 42154 79520
rect 42154 79464 42190 79520
rect 42126 79460 42190 79464
rect 4876 79452 4940 79456
rect 4876 79396 4880 79452
rect 4880 79396 4936 79452
rect 4936 79396 4940 79452
rect 4876 79392 4940 79396
rect 4956 79452 5020 79456
rect 4956 79396 4960 79452
rect 4960 79396 5016 79452
rect 5016 79396 5020 79452
rect 4956 79392 5020 79396
rect 5036 79452 5100 79456
rect 5036 79396 5040 79452
rect 5040 79396 5096 79452
rect 5096 79396 5100 79452
rect 5036 79392 5100 79396
rect 5116 79452 5180 79456
rect 5116 79396 5120 79452
rect 5120 79396 5176 79452
rect 5176 79396 5180 79452
rect 5116 79392 5180 79396
rect 106660 79452 106724 79456
rect 106660 79396 106664 79452
rect 106664 79396 106720 79452
rect 106720 79396 106724 79452
rect 106660 79392 106724 79396
rect 106740 79452 106804 79456
rect 106740 79396 106744 79452
rect 106744 79396 106800 79452
rect 106800 79396 106804 79452
rect 106740 79392 106804 79396
rect 106820 79452 106884 79456
rect 106820 79396 106824 79452
rect 106824 79396 106880 79452
rect 106880 79396 106884 79452
rect 106820 79392 106884 79396
rect 106900 79452 106964 79456
rect 106900 79396 106904 79452
rect 106904 79396 106960 79452
rect 106960 79396 106964 79452
rect 106900 79392 106964 79396
rect 32812 79112 32876 79116
rect 32812 79056 32862 79112
rect 32862 79056 32876 79112
rect 32812 79052 32876 79056
rect 4216 78908 4280 78912
rect 4216 78852 4220 78908
rect 4220 78852 4276 78908
rect 4276 78852 4280 78908
rect 4216 78848 4280 78852
rect 4296 78908 4360 78912
rect 4296 78852 4300 78908
rect 4300 78852 4356 78908
rect 4356 78852 4360 78908
rect 4296 78848 4360 78852
rect 4376 78908 4440 78912
rect 4376 78852 4380 78908
rect 4380 78852 4436 78908
rect 4436 78852 4440 78908
rect 4376 78848 4440 78852
rect 4456 78908 4520 78912
rect 4456 78852 4460 78908
rect 4460 78852 4516 78908
rect 4516 78852 4520 78908
rect 4456 78848 4520 78852
rect 105924 78908 105988 78912
rect 105924 78852 105928 78908
rect 105928 78852 105984 78908
rect 105984 78852 105988 78908
rect 105924 78848 105988 78852
rect 106004 78908 106068 78912
rect 106004 78852 106008 78908
rect 106008 78852 106064 78908
rect 106064 78852 106068 78908
rect 106004 78848 106068 78852
rect 106084 78908 106148 78912
rect 106084 78852 106088 78908
rect 106088 78852 106144 78908
rect 106144 78852 106148 78908
rect 106084 78848 106148 78852
rect 106164 78908 106228 78912
rect 106164 78852 106168 78908
rect 106168 78852 106224 78908
rect 106224 78852 106228 78908
rect 106164 78848 106228 78852
rect 4876 78364 4940 78368
rect 4876 78308 4880 78364
rect 4880 78308 4936 78364
rect 4936 78308 4940 78364
rect 4876 78304 4940 78308
rect 4956 78364 5020 78368
rect 4956 78308 4960 78364
rect 4960 78308 5016 78364
rect 5016 78308 5020 78364
rect 4956 78304 5020 78308
rect 5036 78364 5100 78368
rect 5036 78308 5040 78364
rect 5040 78308 5096 78364
rect 5096 78308 5100 78364
rect 5036 78304 5100 78308
rect 5116 78364 5180 78368
rect 5116 78308 5120 78364
rect 5120 78308 5176 78364
rect 5176 78308 5180 78364
rect 5116 78304 5180 78308
rect 106660 78364 106724 78368
rect 106660 78308 106664 78364
rect 106664 78308 106720 78364
rect 106720 78308 106724 78364
rect 106660 78304 106724 78308
rect 106740 78364 106804 78368
rect 106740 78308 106744 78364
rect 106744 78308 106800 78364
rect 106800 78308 106804 78364
rect 106740 78304 106804 78308
rect 106820 78364 106884 78368
rect 106820 78308 106824 78364
rect 106824 78308 106880 78364
rect 106880 78308 106884 78364
rect 106820 78304 106884 78308
rect 106900 78364 106964 78368
rect 106900 78308 106904 78364
rect 106904 78308 106960 78364
rect 106960 78308 106964 78364
rect 106900 78304 106964 78308
rect 4216 77820 4280 77824
rect 4216 77764 4220 77820
rect 4220 77764 4276 77820
rect 4276 77764 4280 77820
rect 4216 77760 4280 77764
rect 4296 77820 4360 77824
rect 4296 77764 4300 77820
rect 4300 77764 4356 77820
rect 4356 77764 4360 77820
rect 4296 77760 4360 77764
rect 4376 77820 4440 77824
rect 4376 77764 4380 77820
rect 4380 77764 4436 77820
rect 4436 77764 4440 77820
rect 4376 77760 4440 77764
rect 4456 77820 4520 77824
rect 4456 77764 4460 77820
rect 4460 77764 4516 77820
rect 4516 77764 4520 77820
rect 4456 77760 4520 77764
rect 34936 77820 35000 77824
rect 34936 77764 34940 77820
rect 34940 77764 34996 77820
rect 34996 77764 35000 77820
rect 34936 77760 35000 77764
rect 35016 77820 35080 77824
rect 35016 77764 35020 77820
rect 35020 77764 35076 77820
rect 35076 77764 35080 77820
rect 35016 77760 35080 77764
rect 35096 77820 35160 77824
rect 35096 77764 35100 77820
rect 35100 77764 35156 77820
rect 35156 77764 35160 77820
rect 35096 77760 35160 77764
rect 35176 77820 35240 77824
rect 35176 77764 35180 77820
rect 35180 77764 35236 77820
rect 35236 77764 35240 77820
rect 35176 77760 35240 77764
rect 65656 77820 65720 77824
rect 65656 77764 65660 77820
rect 65660 77764 65716 77820
rect 65716 77764 65720 77820
rect 65656 77760 65720 77764
rect 65736 77820 65800 77824
rect 65736 77764 65740 77820
rect 65740 77764 65796 77820
rect 65796 77764 65800 77820
rect 65736 77760 65800 77764
rect 65816 77820 65880 77824
rect 65816 77764 65820 77820
rect 65820 77764 65876 77820
rect 65876 77764 65880 77820
rect 65816 77760 65880 77764
rect 65896 77820 65960 77824
rect 65896 77764 65900 77820
rect 65900 77764 65956 77820
rect 65956 77764 65960 77820
rect 65896 77760 65960 77764
rect 96376 77820 96440 77824
rect 96376 77764 96380 77820
rect 96380 77764 96436 77820
rect 96436 77764 96440 77820
rect 96376 77760 96440 77764
rect 96456 77820 96520 77824
rect 96456 77764 96460 77820
rect 96460 77764 96516 77820
rect 96516 77764 96520 77820
rect 96456 77760 96520 77764
rect 96536 77820 96600 77824
rect 96536 77764 96540 77820
rect 96540 77764 96596 77820
rect 96596 77764 96600 77820
rect 96536 77760 96600 77764
rect 96616 77820 96680 77824
rect 96616 77764 96620 77820
rect 96620 77764 96676 77820
rect 96676 77764 96680 77820
rect 96616 77760 96680 77764
rect 105924 77820 105988 77824
rect 105924 77764 105928 77820
rect 105928 77764 105984 77820
rect 105984 77764 105988 77820
rect 105924 77760 105988 77764
rect 106004 77820 106068 77824
rect 106004 77764 106008 77820
rect 106008 77764 106064 77820
rect 106064 77764 106068 77820
rect 106004 77760 106068 77764
rect 106084 77820 106148 77824
rect 106084 77764 106088 77820
rect 106088 77764 106144 77820
rect 106144 77764 106148 77820
rect 106084 77760 106148 77764
rect 106164 77820 106228 77824
rect 106164 77764 106168 77820
rect 106168 77764 106224 77820
rect 106224 77764 106228 77820
rect 106164 77760 106228 77764
rect 90404 77692 90468 77756
rect 90956 77556 91020 77620
rect 90772 77420 90836 77484
rect 4876 77276 4940 77280
rect 4876 77220 4880 77276
rect 4880 77220 4936 77276
rect 4936 77220 4940 77276
rect 4876 77216 4940 77220
rect 4956 77276 5020 77280
rect 4956 77220 4960 77276
rect 4960 77220 5016 77276
rect 5016 77220 5020 77276
rect 4956 77216 5020 77220
rect 5036 77276 5100 77280
rect 5036 77220 5040 77276
rect 5040 77220 5096 77276
rect 5096 77220 5100 77276
rect 5036 77216 5100 77220
rect 5116 77276 5180 77280
rect 5116 77220 5120 77276
rect 5120 77220 5176 77276
rect 5176 77220 5180 77276
rect 5116 77216 5180 77220
rect 35596 77276 35660 77280
rect 35596 77220 35600 77276
rect 35600 77220 35656 77276
rect 35656 77220 35660 77276
rect 35596 77216 35660 77220
rect 35676 77276 35740 77280
rect 35676 77220 35680 77276
rect 35680 77220 35736 77276
rect 35736 77220 35740 77276
rect 35676 77216 35740 77220
rect 35756 77276 35820 77280
rect 35756 77220 35760 77276
rect 35760 77220 35816 77276
rect 35816 77220 35820 77276
rect 35756 77216 35820 77220
rect 35836 77276 35900 77280
rect 35836 77220 35840 77276
rect 35840 77220 35896 77276
rect 35896 77220 35900 77276
rect 35836 77216 35900 77220
rect 66316 77276 66380 77280
rect 66316 77220 66320 77276
rect 66320 77220 66376 77276
rect 66376 77220 66380 77276
rect 66316 77216 66380 77220
rect 66396 77276 66460 77280
rect 66396 77220 66400 77276
rect 66400 77220 66456 77276
rect 66456 77220 66460 77276
rect 66396 77216 66460 77220
rect 66476 77276 66540 77280
rect 66476 77220 66480 77276
rect 66480 77220 66536 77276
rect 66536 77220 66540 77276
rect 66476 77216 66540 77220
rect 66556 77276 66620 77280
rect 66556 77220 66560 77276
rect 66560 77220 66616 77276
rect 66616 77220 66620 77276
rect 66556 77216 66620 77220
rect 97036 77276 97100 77280
rect 97036 77220 97040 77276
rect 97040 77220 97096 77276
rect 97096 77220 97100 77276
rect 97036 77216 97100 77220
rect 97116 77276 97180 77280
rect 97116 77220 97120 77276
rect 97120 77220 97176 77276
rect 97176 77220 97180 77276
rect 97116 77216 97180 77220
rect 97196 77276 97260 77280
rect 97196 77220 97200 77276
rect 97200 77220 97256 77276
rect 97256 77220 97260 77276
rect 97196 77216 97260 77220
rect 97276 77276 97340 77280
rect 97276 77220 97280 77276
rect 97280 77220 97336 77276
rect 97336 77220 97340 77276
rect 97276 77216 97340 77220
rect 106660 77276 106724 77280
rect 106660 77220 106664 77276
rect 106664 77220 106720 77276
rect 106720 77220 106724 77276
rect 106660 77216 106724 77220
rect 106740 77276 106804 77280
rect 106740 77220 106744 77276
rect 106744 77220 106800 77276
rect 106800 77220 106804 77276
rect 106740 77216 106804 77220
rect 106820 77276 106884 77280
rect 106820 77220 106824 77276
rect 106824 77220 106880 77276
rect 106880 77220 106884 77276
rect 106820 77216 106884 77220
rect 106900 77276 106964 77280
rect 106900 77220 106904 77276
rect 106904 77220 106960 77276
rect 106960 77220 106964 77276
rect 106900 77216 106964 77220
rect 4216 76732 4280 76736
rect 4216 76676 4220 76732
rect 4220 76676 4276 76732
rect 4276 76676 4280 76732
rect 4216 76672 4280 76676
rect 4296 76732 4360 76736
rect 4296 76676 4300 76732
rect 4300 76676 4356 76732
rect 4356 76676 4360 76732
rect 4296 76672 4360 76676
rect 4376 76732 4440 76736
rect 4376 76676 4380 76732
rect 4380 76676 4436 76732
rect 4436 76676 4440 76732
rect 4376 76672 4440 76676
rect 4456 76732 4520 76736
rect 4456 76676 4460 76732
rect 4460 76676 4516 76732
rect 4516 76676 4520 76732
rect 4456 76672 4520 76676
rect 34936 76732 35000 76736
rect 34936 76676 34940 76732
rect 34940 76676 34996 76732
rect 34996 76676 35000 76732
rect 34936 76672 35000 76676
rect 35016 76732 35080 76736
rect 35016 76676 35020 76732
rect 35020 76676 35076 76732
rect 35076 76676 35080 76732
rect 35016 76672 35080 76676
rect 35096 76732 35160 76736
rect 35096 76676 35100 76732
rect 35100 76676 35156 76732
rect 35156 76676 35160 76732
rect 35096 76672 35160 76676
rect 35176 76732 35240 76736
rect 35176 76676 35180 76732
rect 35180 76676 35236 76732
rect 35236 76676 35240 76732
rect 35176 76672 35240 76676
rect 65656 76732 65720 76736
rect 65656 76676 65660 76732
rect 65660 76676 65716 76732
rect 65716 76676 65720 76732
rect 65656 76672 65720 76676
rect 65736 76732 65800 76736
rect 65736 76676 65740 76732
rect 65740 76676 65796 76732
rect 65796 76676 65800 76732
rect 65736 76672 65800 76676
rect 65816 76732 65880 76736
rect 65816 76676 65820 76732
rect 65820 76676 65876 76732
rect 65876 76676 65880 76732
rect 65816 76672 65880 76676
rect 65896 76732 65960 76736
rect 65896 76676 65900 76732
rect 65900 76676 65956 76732
rect 65956 76676 65960 76732
rect 65896 76672 65960 76676
rect 96376 76732 96440 76736
rect 96376 76676 96380 76732
rect 96380 76676 96436 76732
rect 96436 76676 96440 76732
rect 96376 76672 96440 76676
rect 96456 76732 96520 76736
rect 96456 76676 96460 76732
rect 96460 76676 96516 76732
rect 96516 76676 96520 76732
rect 96456 76672 96520 76676
rect 96536 76732 96600 76736
rect 96536 76676 96540 76732
rect 96540 76676 96596 76732
rect 96596 76676 96600 76732
rect 96536 76672 96600 76676
rect 96616 76732 96680 76736
rect 96616 76676 96620 76732
rect 96620 76676 96676 76732
rect 96676 76676 96680 76732
rect 96616 76672 96680 76676
rect 4876 76188 4940 76192
rect 4876 76132 4880 76188
rect 4880 76132 4936 76188
rect 4936 76132 4940 76188
rect 4876 76128 4940 76132
rect 4956 76188 5020 76192
rect 4956 76132 4960 76188
rect 4960 76132 5016 76188
rect 5016 76132 5020 76188
rect 4956 76128 5020 76132
rect 5036 76188 5100 76192
rect 5036 76132 5040 76188
rect 5040 76132 5096 76188
rect 5096 76132 5100 76188
rect 5036 76128 5100 76132
rect 5116 76188 5180 76192
rect 5116 76132 5120 76188
rect 5120 76132 5176 76188
rect 5176 76132 5180 76188
rect 5116 76128 5180 76132
rect 35596 76188 35660 76192
rect 35596 76132 35600 76188
rect 35600 76132 35656 76188
rect 35656 76132 35660 76188
rect 35596 76128 35660 76132
rect 35676 76188 35740 76192
rect 35676 76132 35680 76188
rect 35680 76132 35736 76188
rect 35736 76132 35740 76188
rect 35676 76128 35740 76132
rect 35756 76188 35820 76192
rect 35756 76132 35760 76188
rect 35760 76132 35816 76188
rect 35816 76132 35820 76188
rect 35756 76128 35820 76132
rect 35836 76188 35900 76192
rect 35836 76132 35840 76188
rect 35840 76132 35896 76188
rect 35896 76132 35900 76188
rect 35836 76128 35900 76132
rect 66316 76188 66380 76192
rect 66316 76132 66320 76188
rect 66320 76132 66376 76188
rect 66376 76132 66380 76188
rect 66316 76128 66380 76132
rect 66396 76188 66460 76192
rect 66396 76132 66400 76188
rect 66400 76132 66456 76188
rect 66456 76132 66460 76188
rect 66396 76128 66460 76132
rect 66476 76188 66540 76192
rect 66476 76132 66480 76188
rect 66480 76132 66536 76188
rect 66536 76132 66540 76188
rect 66476 76128 66540 76132
rect 66556 76188 66620 76192
rect 66556 76132 66560 76188
rect 66560 76132 66616 76188
rect 66616 76132 66620 76188
rect 66556 76128 66620 76132
rect 97036 76188 97100 76192
rect 97036 76132 97040 76188
rect 97040 76132 97096 76188
rect 97096 76132 97100 76188
rect 97036 76128 97100 76132
rect 97116 76188 97180 76192
rect 97116 76132 97120 76188
rect 97120 76132 97176 76188
rect 97176 76132 97180 76188
rect 97116 76128 97180 76132
rect 97196 76188 97260 76192
rect 97196 76132 97200 76188
rect 97200 76132 97256 76188
rect 97256 76132 97260 76188
rect 97196 76128 97260 76132
rect 97276 76188 97340 76192
rect 97276 76132 97280 76188
rect 97280 76132 97336 76188
rect 97336 76132 97340 76188
rect 97276 76128 97340 76132
rect 4216 75644 4280 75648
rect 4216 75588 4220 75644
rect 4220 75588 4276 75644
rect 4276 75588 4280 75644
rect 4216 75584 4280 75588
rect 4296 75644 4360 75648
rect 4296 75588 4300 75644
rect 4300 75588 4356 75644
rect 4356 75588 4360 75644
rect 4296 75584 4360 75588
rect 4376 75644 4440 75648
rect 4376 75588 4380 75644
rect 4380 75588 4436 75644
rect 4436 75588 4440 75644
rect 4376 75584 4440 75588
rect 4456 75644 4520 75648
rect 4456 75588 4460 75644
rect 4460 75588 4516 75644
rect 4516 75588 4520 75644
rect 4456 75584 4520 75588
rect 34936 75644 35000 75648
rect 34936 75588 34940 75644
rect 34940 75588 34996 75644
rect 34996 75588 35000 75644
rect 34936 75584 35000 75588
rect 35016 75644 35080 75648
rect 35016 75588 35020 75644
rect 35020 75588 35076 75644
rect 35076 75588 35080 75644
rect 35016 75584 35080 75588
rect 35096 75644 35160 75648
rect 35096 75588 35100 75644
rect 35100 75588 35156 75644
rect 35156 75588 35160 75644
rect 35096 75584 35160 75588
rect 35176 75644 35240 75648
rect 35176 75588 35180 75644
rect 35180 75588 35236 75644
rect 35236 75588 35240 75644
rect 35176 75584 35240 75588
rect 65656 75644 65720 75648
rect 65656 75588 65660 75644
rect 65660 75588 65716 75644
rect 65716 75588 65720 75644
rect 65656 75584 65720 75588
rect 65736 75644 65800 75648
rect 65736 75588 65740 75644
rect 65740 75588 65796 75644
rect 65796 75588 65800 75644
rect 65736 75584 65800 75588
rect 65816 75644 65880 75648
rect 65816 75588 65820 75644
rect 65820 75588 65876 75644
rect 65876 75588 65880 75644
rect 65816 75584 65880 75588
rect 65896 75644 65960 75648
rect 65896 75588 65900 75644
rect 65900 75588 65956 75644
rect 65956 75588 65960 75644
rect 65896 75584 65960 75588
rect 96376 75644 96440 75648
rect 96376 75588 96380 75644
rect 96380 75588 96436 75644
rect 96436 75588 96440 75644
rect 96376 75584 96440 75588
rect 96456 75644 96520 75648
rect 96456 75588 96460 75644
rect 96460 75588 96516 75644
rect 96516 75588 96520 75644
rect 96456 75584 96520 75588
rect 96536 75644 96600 75648
rect 96536 75588 96540 75644
rect 96540 75588 96596 75644
rect 96596 75588 96600 75644
rect 96536 75584 96600 75588
rect 96616 75644 96680 75648
rect 96616 75588 96620 75644
rect 96620 75588 96676 75644
rect 96676 75588 96680 75644
rect 96616 75584 96680 75588
rect 4876 75100 4940 75104
rect 4876 75044 4880 75100
rect 4880 75044 4936 75100
rect 4936 75044 4940 75100
rect 4876 75040 4940 75044
rect 4956 75100 5020 75104
rect 4956 75044 4960 75100
rect 4960 75044 5016 75100
rect 5016 75044 5020 75100
rect 4956 75040 5020 75044
rect 5036 75100 5100 75104
rect 5036 75044 5040 75100
rect 5040 75044 5096 75100
rect 5096 75044 5100 75100
rect 5036 75040 5100 75044
rect 5116 75100 5180 75104
rect 5116 75044 5120 75100
rect 5120 75044 5176 75100
rect 5176 75044 5180 75100
rect 5116 75040 5180 75044
rect 35596 75100 35660 75104
rect 35596 75044 35600 75100
rect 35600 75044 35656 75100
rect 35656 75044 35660 75100
rect 35596 75040 35660 75044
rect 35676 75100 35740 75104
rect 35676 75044 35680 75100
rect 35680 75044 35736 75100
rect 35736 75044 35740 75100
rect 35676 75040 35740 75044
rect 35756 75100 35820 75104
rect 35756 75044 35760 75100
rect 35760 75044 35816 75100
rect 35816 75044 35820 75100
rect 35756 75040 35820 75044
rect 35836 75100 35900 75104
rect 35836 75044 35840 75100
rect 35840 75044 35896 75100
rect 35896 75044 35900 75100
rect 35836 75040 35900 75044
rect 66316 75100 66380 75104
rect 66316 75044 66320 75100
rect 66320 75044 66376 75100
rect 66376 75044 66380 75100
rect 66316 75040 66380 75044
rect 66396 75100 66460 75104
rect 66396 75044 66400 75100
rect 66400 75044 66456 75100
rect 66456 75044 66460 75100
rect 66396 75040 66460 75044
rect 66476 75100 66540 75104
rect 66476 75044 66480 75100
rect 66480 75044 66536 75100
rect 66536 75044 66540 75100
rect 66476 75040 66540 75044
rect 66556 75100 66620 75104
rect 66556 75044 66560 75100
rect 66560 75044 66616 75100
rect 66616 75044 66620 75100
rect 66556 75040 66620 75044
rect 97036 75100 97100 75104
rect 97036 75044 97040 75100
rect 97040 75044 97096 75100
rect 97096 75044 97100 75100
rect 97036 75040 97100 75044
rect 97116 75100 97180 75104
rect 97116 75044 97120 75100
rect 97120 75044 97176 75100
rect 97176 75044 97180 75100
rect 97116 75040 97180 75044
rect 97196 75100 97260 75104
rect 97196 75044 97200 75100
rect 97200 75044 97256 75100
rect 97256 75044 97260 75100
rect 97196 75040 97260 75044
rect 97276 75100 97340 75104
rect 97276 75044 97280 75100
rect 97280 75044 97336 75100
rect 97336 75044 97340 75100
rect 97276 75040 97340 75044
rect 4216 74556 4280 74560
rect 4216 74500 4220 74556
rect 4220 74500 4276 74556
rect 4276 74500 4280 74556
rect 4216 74496 4280 74500
rect 4296 74556 4360 74560
rect 4296 74500 4300 74556
rect 4300 74500 4356 74556
rect 4356 74500 4360 74556
rect 4296 74496 4360 74500
rect 4376 74556 4440 74560
rect 4376 74500 4380 74556
rect 4380 74500 4436 74556
rect 4436 74500 4440 74556
rect 4376 74496 4440 74500
rect 4456 74556 4520 74560
rect 4456 74500 4460 74556
rect 4460 74500 4516 74556
rect 4516 74500 4520 74556
rect 4456 74496 4520 74500
rect 34936 74556 35000 74560
rect 34936 74500 34940 74556
rect 34940 74500 34996 74556
rect 34996 74500 35000 74556
rect 34936 74496 35000 74500
rect 35016 74556 35080 74560
rect 35016 74500 35020 74556
rect 35020 74500 35076 74556
rect 35076 74500 35080 74556
rect 35016 74496 35080 74500
rect 35096 74556 35160 74560
rect 35096 74500 35100 74556
rect 35100 74500 35156 74556
rect 35156 74500 35160 74556
rect 35096 74496 35160 74500
rect 35176 74556 35240 74560
rect 35176 74500 35180 74556
rect 35180 74500 35236 74556
rect 35236 74500 35240 74556
rect 35176 74496 35240 74500
rect 65656 74556 65720 74560
rect 65656 74500 65660 74556
rect 65660 74500 65716 74556
rect 65716 74500 65720 74556
rect 65656 74496 65720 74500
rect 65736 74556 65800 74560
rect 65736 74500 65740 74556
rect 65740 74500 65796 74556
rect 65796 74500 65800 74556
rect 65736 74496 65800 74500
rect 65816 74556 65880 74560
rect 65816 74500 65820 74556
rect 65820 74500 65876 74556
rect 65876 74500 65880 74556
rect 65816 74496 65880 74500
rect 65896 74556 65960 74560
rect 65896 74500 65900 74556
rect 65900 74500 65956 74556
rect 65956 74500 65960 74556
rect 65896 74496 65960 74500
rect 96376 74556 96440 74560
rect 96376 74500 96380 74556
rect 96380 74500 96436 74556
rect 96436 74500 96440 74556
rect 96376 74496 96440 74500
rect 96456 74556 96520 74560
rect 96456 74500 96460 74556
rect 96460 74500 96516 74556
rect 96516 74500 96520 74556
rect 96456 74496 96520 74500
rect 96536 74556 96600 74560
rect 96536 74500 96540 74556
rect 96540 74500 96596 74556
rect 96596 74500 96600 74556
rect 96536 74496 96600 74500
rect 96616 74556 96680 74560
rect 96616 74500 96620 74556
rect 96620 74500 96676 74556
rect 96676 74500 96680 74556
rect 96616 74496 96680 74500
rect 4876 74012 4940 74016
rect 4876 73956 4880 74012
rect 4880 73956 4936 74012
rect 4936 73956 4940 74012
rect 4876 73952 4940 73956
rect 4956 74012 5020 74016
rect 4956 73956 4960 74012
rect 4960 73956 5016 74012
rect 5016 73956 5020 74012
rect 4956 73952 5020 73956
rect 5036 74012 5100 74016
rect 5036 73956 5040 74012
rect 5040 73956 5096 74012
rect 5096 73956 5100 74012
rect 5036 73952 5100 73956
rect 5116 74012 5180 74016
rect 5116 73956 5120 74012
rect 5120 73956 5176 74012
rect 5176 73956 5180 74012
rect 5116 73952 5180 73956
rect 35596 74012 35660 74016
rect 35596 73956 35600 74012
rect 35600 73956 35656 74012
rect 35656 73956 35660 74012
rect 35596 73952 35660 73956
rect 35676 74012 35740 74016
rect 35676 73956 35680 74012
rect 35680 73956 35736 74012
rect 35736 73956 35740 74012
rect 35676 73952 35740 73956
rect 35756 74012 35820 74016
rect 35756 73956 35760 74012
rect 35760 73956 35816 74012
rect 35816 73956 35820 74012
rect 35756 73952 35820 73956
rect 35836 74012 35900 74016
rect 35836 73956 35840 74012
rect 35840 73956 35896 74012
rect 35896 73956 35900 74012
rect 35836 73952 35900 73956
rect 66316 74012 66380 74016
rect 66316 73956 66320 74012
rect 66320 73956 66376 74012
rect 66376 73956 66380 74012
rect 66316 73952 66380 73956
rect 66396 74012 66460 74016
rect 66396 73956 66400 74012
rect 66400 73956 66456 74012
rect 66456 73956 66460 74012
rect 66396 73952 66460 73956
rect 66476 74012 66540 74016
rect 66476 73956 66480 74012
rect 66480 73956 66536 74012
rect 66536 73956 66540 74012
rect 66476 73952 66540 73956
rect 66556 74012 66620 74016
rect 66556 73956 66560 74012
rect 66560 73956 66616 74012
rect 66616 73956 66620 74012
rect 66556 73952 66620 73956
rect 97036 74012 97100 74016
rect 97036 73956 97040 74012
rect 97040 73956 97096 74012
rect 97096 73956 97100 74012
rect 97036 73952 97100 73956
rect 97116 74012 97180 74016
rect 97116 73956 97120 74012
rect 97120 73956 97176 74012
rect 97176 73956 97180 74012
rect 97116 73952 97180 73956
rect 97196 74012 97260 74016
rect 97196 73956 97200 74012
rect 97200 73956 97256 74012
rect 97256 73956 97260 74012
rect 97196 73952 97260 73956
rect 97276 74012 97340 74016
rect 97276 73956 97280 74012
rect 97280 73956 97336 74012
rect 97336 73956 97340 74012
rect 97276 73952 97340 73956
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 34936 73468 35000 73472
rect 34936 73412 34940 73468
rect 34940 73412 34996 73468
rect 34996 73412 35000 73468
rect 34936 73408 35000 73412
rect 35016 73468 35080 73472
rect 35016 73412 35020 73468
rect 35020 73412 35076 73468
rect 35076 73412 35080 73468
rect 35016 73408 35080 73412
rect 35096 73468 35160 73472
rect 35096 73412 35100 73468
rect 35100 73412 35156 73468
rect 35156 73412 35160 73468
rect 35096 73408 35160 73412
rect 35176 73468 35240 73472
rect 35176 73412 35180 73468
rect 35180 73412 35236 73468
rect 35236 73412 35240 73468
rect 35176 73408 35240 73412
rect 65656 73468 65720 73472
rect 65656 73412 65660 73468
rect 65660 73412 65716 73468
rect 65716 73412 65720 73468
rect 65656 73408 65720 73412
rect 65736 73468 65800 73472
rect 65736 73412 65740 73468
rect 65740 73412 65796 73468
rect 65796 73412 65800 73468
rect 65736 73408 65800 73412
rect 65816 73468 65880 73472
rect 65816 73412 65820 73468
rect 65820 73412 65876 73468
rect 65876 73412 65880 73468
rect 65816 73408 65880 73412
rect 65896 73468 65960 73472
rect 65896 73412 65900 73468
rect 65900 73412 65956 73468
rect 65956 73412 65960 73468
rect 65896 73408 65960 73412
rect 96376 73468 96440 73472
rect 96376 73412 96380 73468
rect 96380 73412 96436 73468
rect 96436 73412 96440 73468
rect 96376 73408 96440 73412
rect 96456 73468 96520 73472
rect 96456 73412 96460 73468
rect 96460 73412 96516 73468
rect 96516 73412 96520 73468
rect 96456 73408 96520 73412
rect 96536 73468 96600 73472
rect 96536 73412 96540 73468
rect 96540 73412 96596 73468
rect 96596 73412 96600 73468
rect 96536 73408 96600 73412
rect 96616 73468 96680 73472
rect 96616 73412 96620 73468
rect 96620 73412 96676 73468
rect 96676 73412 96680 73468
rect 96616 73408 96680 73412
rect 4876 72924 4940 72928
rect 4876 72868 4880 72924
rect 4880 72868 4936 72924
rect 4936 72868 4940 72924
rect 4876 72864 4940 72868
rect 4956 72924 5020 72928
rect 4956 72868 4960 72924
rect 4960 72868 5016 72924
rect 5016 72868 5020 72924
rect 4956 72864 5020 72868
rect 5036 72924 5100 72928
rect 5036 72868 5040 72924
rect 5040 72868 5096 72924
rect 5096 72868 5100 72924
rect 5036 72864 5100 72868
rect 5116 72924 5180 72928
rect 5116 72868 5120 72924
rect 5120 72868 5176 72924
rect 5176 72868 5180 72924
rect 5116 72864 5180 72868
rect 35596 72924 35660 72928
rect 35596 72868 35600 72924
rect 35600 72868 35656 72924
rect 35656 72868 35660 72924
rect 35596 72864 35660 72868
rect 35676 72924 35740 72928
rect 35676 72868 35680 72924
rect 35680 72868 35736 72924
rect 35736 72868 35740 72924
rect 35676 72864 35740 72868
rect 35756 72924 35820 72928
rect 35756 72868 35760 72924
rect 35760 72868 35816 72924
rect 35816 72868 35820 72924
rect 35756 72864 35820 72868
rect 35836 72924 35900 72928
rect 35836 72868 35840 72924
rect 35840 72868 35896 72924
rect 35896 72868 35900 72924
rect 35836 72864 35900 72868
rect 66316 72924 66380 72928
rect 66316 72868 66320 72924
rect 66320 72868 66376 72924
rect 66376 72868 66380 72924
rect 66316 72864 66380 72868
rect 66396 72924 66460 72928
rect 66396 72868 66400 72924
rect 66400 72868 66456 72924
rect 66456 72868 66460 72924
rect 66396 72864 66460 72868
rect 66476 72924 66540 72928
rect 66476 72868 66480 72924
rect 66480 72868 66536 72924
rect 66536 72868 66540 72924
rect 66476 72864 66540 72868
rect 66556 72924 66620 72928
rect 66556 72868 66560 72924
rect 66560 72868 66616 72924
rect 66616 72868 66620 72924
rect 66556 72864 66620 72868
rect 97036 72924 97100 72928
rect 97036 72868 97040 72924
rect 97040 72868 97096 72924
rect 97096 72868 97100 72924
rect 97036 72864 97100 72868
rect 97116 72924 97180 72928
rect 97116 72868 97120 72924
rect 97120 72868 97176 72924
rect 97176 72868 97180 72924
rect 97116 72864 97180 72868
rect 97196 72924 97260 72928
rect 97196 72868 97200 72924
rect 97200 72868 97256 72924
rect 97256 72868 97260 72924
rect 97196 72864 97260 72868
rect 97276 72924 97340 72928
rect 97276 72868 97280 72924
rect 97280 72868 97336 72924
rect 97336 72868 97340 72924
rect 97276 72864 97340 72868
rect 86172 72524 86236 72588
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 34936 72380 35000 72384
rect 34936 72324 34940 72380
rect 34940 72324 34996 72380
rect 34996 72324 35000 72380
rect 34936 72320 35000 72324
rect 35016 72380 35080 72384
rect 35016 72324 35020 72380
rect 35020 72324 35076 72380
rect 35076 72324 35080 72380
rect 35016 72320 35080 72324
rect 35096 72380 35160 72384
rect 35096 72324 35100 72380
rect 35100 72324 35156 72380
rect 35156 72324 35160 72380
rect 35096 72320 35160 72324
rect 35176 72380 35240 72384
rect 35176 72324 35180 72380
rect 35180 72324 35236 72380
rect 35236 72324 35240 72380
rect 35176 72320 35240 72324
rect 65656 72380 65720 72384
rect 65656 72324 65660 72380
rect 65660 72324 65716 72380
rect 65716 72324 65720 72380
rect 65656 72320 65720 72324
rect 65736 72380 65800 72384
rect 65736 72324 65740 72380
rect 65740 72324 65796 72380
rect 65796 72324 65800 72380
rect 65736 72320 65800 72324
rect 65816 72380 65880 72384
rect 65816 72324 65820 72380
rect 65820 72324 65876 72380
rect 65876 72324 65880 72380
rect 65816 72320 65880 72324
rect 65896 72380 65960 72384
rect 65896 72324 65900 72380
rect 65900 72324 65956 72380
rect 65956 72324 65960 72380
rect 65896 72320 65960 72324
rect 96376 72380 96440 72384
rect 96376 72324 96380 72380
rect 96380 72324 96436 72380
rect 96436 72324 96440 72380
rect 96376 72320 96440 72324
rect 96456 72380 96520 72384
rect 96456 72324 96460 72380
rect 96460 72324 96516 72380
rect 96516 72324 96520 72380
rect 96456 72320 96520 72324
rect 96536 72380 96600 72384
rect 96536 72324 96540 72380
rect 96540 72324 96596 72380
rect 96596 72324 96600 72380
rect 96536 72320 96600 72324
rect 96616 72380 96680 72384
rect 96616 72324 96620 72380
rect 96620 72324 96676 72380
rect 96676 72324 96680 72380
rect 96616 72320 96680 72324
rect 4876 71836 4940 71840
rect 4876 71780 4880 71836
rect 4880 71780 4936 71836
rect 4936 71780 4940 71836
rect 4876 71776 4940 71780
rect 4956 71836 5020 71840
rect 4956 71780 4960 71836
rect 4960 71780 5016 71836
rect 5016 71780 5020 71836
rect 4956 71776 5020 71780
rect 5036 71836 5100 71840
rect 5036 71780 5040 71836
rect 5040 71780 5096 71836
rect 5096 71780 5100 71836
rect 5036 71776 5100 71780
rect 5116 71836 5180 71840
rect 5116 71780 5120 71836
rect 5120 71780 5176 71836
rect 5176 71780 5180 71836
rect 5116 71776 5180 71780
rect 35596 71836 35660 71840
rect 35596 71780 35600 71836
rect 35600 71780 35656 71836
rect 35656 71780 35660 71836
rect 35596 71776 35660 71780
rect 35676 71836 35740 71840
rect 35676 71780 35680 71836
rect 35680 71780 35736 71836
rect 35736 71780 35740 71836
rect 35676 71776 35740 71780
rect 35756 71836 35820 71840
rect 35756 71780 35760 71836
rect 35760 71780 35816 71836
rect 35816 71780 35820 71836
rect 35756 71776 35820 71780
rect 35836 71836 35900 71840
rect 35836 71780 35840 71836
rect 35840 71780 35896 71836
rect 35896 71780 35900 71836
rect 35836 71776 35900 71780
rect 66316 71836 66380 71840
rect 66316 71780 66320 71836
rect 66320 71780 66376 71836
rect 66376 71780 66380 71836
rect 66316 71776 66380 71780
rect 66396 71836 66460 71840
rect 66396 71780 66400 71836
rect 66400 71780 66456 71836
rect 66456 71780 66460 71836
rect 66396 71776 66460 71780
rect 66476 71836 66540 71840
rect 66476 71780 66480 71836
rect 66480 71780 66536 71836
rect 66536 71780 66540 71836
rect 66476 71776 66540 71780
rect 66556 71836 66620 71840
rect 66556 71780 66560 71836
rect 66560 71780 66616 71836
rect 66616 71780 66620 71836
rect 66556 71776 66620 71780
rect 97036 71836 97100 71840
rect 97036 71780 97040 71836
rect 97040 71780 97096 71836
rect 97096 71780 97100 71836
rect 97036 71776 97100 71780
rect 97116 71836 97180 71840
rect 97116 71780 97120 71836
rect 97120 71780 97176 71836
rect 97176 71780 97180 71836
rect 97116 71776 97180 71780
rect 97196 71836 97260 71840
rect 97196 71780 97200 71836
rect 97200 71780 97256 71836
rect 97256 71780 97260 71836
rect 97196 71776 97260 71780
rect 97276 71836 97340 71840
rect 97276 71780 97280 71836
rect 97280 71780 97336 71836
rect 97336 71780 97340 71836
rect 97276 71776 97340 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 34936 71292 35000 71296
rect 34936 71236 34940 71292
rect 34940 71236 34996 71292
rect 34996 71236 35000 71292
rect 34936 71232 35000 71236
rect 35016 71292 35080 71296
rect 35016 71236 35020 71292
rect 35020 71236 35076 71292
rect 35076 71236 35080 71292
rect 35016 71232 35080 71236
rect 35096 71292 35160 71296
rect 35096 71236 35100 71292
rect 35100 71236 35156 71292
rect 35156 71236 35160 71292
rect 35096 71232 35160 71236
rect 35176 71292 35240 71296
rect 35176 71236 35180 71292
rect 35180 71236 35236 71292
rect 35236 71236 35240 71292
rect 35176 71232 35240 71236
rect 65656 71292 65720 71296
rect 65656 71236 65660 71292
rect 65660 71236 65716 71292
rect 65716 71236 65720 71292
rect 65656 71232 65720 71236
rect 65736 71292 65800 71296
rect 65736 71236 65740 71292
rect 65740 71236 65796 71292
rect 65796 71236 65800 71292
rect 65736 71232 65800 71236
rect 65816 71292 65880 71296
rect 65816 71236 65820 71292
rect 65820 71236 65876 71292
rect 65876 71236 65880 71292
rect 65816 71232 65880 71236
rect 65896 71292 65960 71296
rect 65896 71236 65900 71292
rect 65900 71236 65956 71292
rect 65956 71236 65960 71292
rect 65896 71232 65960 71236
rect 96376 71292 96440 71296
rect 96376 71236 96380 71292
rect 96380 71236 96436 71292
rect 96436 71236 96440 71292
rect 96376 71232 96440 71236
rect 96456 71292 96520 71296
rect 96456 71236 96460 71292
rect 96460 71236 96516 71292
rect 96516 71236 96520 71292
rect 96456 71232 96520 71236
rect 96536 71292 96600 71296
rect 96536 71236 96540 71292
rect 96540 71236 96596 71292
rect 96596 71236 96600 71292
rect 96536 71232 96600 71236
rect 96616 71292 96680 71296
rect 96616 71236 96620 71292
rect 96620 71236 96676 71292
rect 96676 71236 96680 71292
rect 96616 71232 96680 71236
rect 4876 70748 4940 70752
rect 4876 70692 4880 70748
rect 4880 70692 4936 70748
rect 4936 70692 4940 70748
rect 4876 70688 4940 70692
rect 4956 70748 5020 70752
rect 4956 70692 4960 70748
rect 4960 70692 5016 70748
rect 5016 70692 5020 70748
rect 4956 70688 5020 70692
rect 5036 70748 5100 70752
rect 5036 70692 5040 70748
rect 5040 70692 5096 70748
rect 5096 70692 5100 70748
rect 5036 70688 5100 70692
rect 5116 70748 5180 70752
rect 5116 70692 5120 70748
rect 5120 70692 5176 70748
rect 5176 70692 5180 70748
rect 5116 70688 5180 70692
rect 35596 70748 35660 70752
rect 35596 70692 35600 70748
rect 35600 70692 35656 70748
rect 35656 70692 35660 70748
rect 35596 70688 35660 70692
rect 35676 70748 35740 70752
rect 35676 70692 35680 70748
rect 35680 70692 35736 70748
rect 35736 70692 35740 70748
rect 35676 70688 35740 70692
rect 35756 70748 35820 70752
rect 35756 70692 35760 70748
rect 35760 70692 35816 70748
rect 35816 70692 35820 70748
rect 35756 70688 35820 70692
rect 35836 70748 35900 70752
rect 35836 70692 35840 70748
rect 35840 70692 35896 70748
rect 35896 70692 35900 70748
rect 35836 70688 35900 70692
rect 66316 70748 66380 70752
rect 66316 70692 66320 70748
rect 66320 70692 66376 70748
rect 66376 70692 66380 70748
rect 66316 70688 66380 70692
rect 66396 70748 66460 70752
rect 66396 70692 66400 70748
rect 66400 70692 66456 70748
rect 66456 70692 66460 70748
rect 66396 70688 66460 70692
rect 66476 70748 66540 70752
rect 66476 70692 66480 70748
rect 66480 70692 66536 70748
rect 66536 70692 66540 70748
rect 66476 70688 66540 70692
rect 66556 70748 66620 70752
rect 66556 70692 66560 70748
rect 66560 70692 66616 70748
rect 66616 70692 66620 70748
rect 66556 70688 66620 70692
rect 97036 70748 97100 70752
rect 97036 70692 97040 70748
rect 97040 70692 97096 70748
rect 97096 70692 97100 70748
rect 97036 70688 97100 70692
rect 97116 70748 97180 70752
rect 97116 70692 97120 70748
rect 97120 70692 97176 70748
rect 97176 70692 97180 70748
rect 97116 70688 97180 70692
rect 97196 70748 97260 70752
rect 97196 70692 97200 70748
rect 97200 70692 97256 70748
rect 97256 70692 97260 70748
rect 97196 70688 97260 70692
rect 97276 70748 97340 70752
rect 97276 70692 97280 70748
rect 97280 70692 97336 70748
rect 97336 70692 97340 70748
rect 97276 70688 97340 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 34936 70204 35000 70208
rect 34936 70148 34940 70204
rect 34940 70148 34996 70204
rect 34996 70148 35000 70204
rect 34936 70144 35000 70148
rect 35016 70204 35080 70208
rect 35016 70148 35020 70204
rect 35020 70148 35076 70204
rect 35076 70148 35080 70204
rect 35016 70144 35080 70148
rect 35096 70204 35160 70208
rect 35096 70148 35100 70204
rect 35100 70148 35156 70204
rect 35156 70148 35160 70204
rect 35096 70144 35160 70148
rect 35176 70204 35240 70208
rect 35176 70148 35180 70204
rect 35180 70148 35236 70204
rect 35236 70148 35240 70204
rect 35176 70144 35240 70148
rect 65656 70204 65720 70208
rect 65656 70148 65660 70204
rect 65660 70148 65716 70204
rect 65716 70148 65720 70204
rect 65656 70144 65720 70148
rect 65736 70204 65800 70208
rect 65736 70148 65740 70204
rect 65740 70148 65796 70204
rect 65796 70148 65800 70204
rect 65736 70144 65800 70148
rect 65816 70204 65880 70208
rect 65816 70148 65820 70204
rect 65820 70148 65876 70204
rect 65876 70148 65880 70204
rect 65816 70144 65880 70148
rect 65896 70204 65960 70208
rect 65896 70148 65900 70204
rect 65900 70148 65956 70204
rect 65956 70148 65960 70204
rect 65896 70144 65960 70148
rect 96376 70204 96440 70208
rect 96376 70148 96380 70204
rect 96380 70148 96436 70204
rect 96436 70148 96440 70204
rect 96376 70144 96440 70148
rect 96456 70204 96520 70208
rect 96456 70148 96460 70204
rect 96460 70148 96516 70204
rect 96516 70148 96520 70204
rect 96456 70144 96520 70148
rect 96536 70204 96600 70208
rect 96536 70148 96540 70204
rect 96540 70148 96596 70204
rect 96596 70148 96600 70204
rect 96536 70144 96600 70148
rect 96616 70204 96680 70208
rect 96616 70148 96620 70204
rect 96620 70148 96676 70204
rect 96676 70148 96680 70204
rect 96616 70144 96680 70148
rect 63540 69804 63604 69868
rect 73660 69804 73724 69868
rect 4876 69660 4940 69664
rect 4876 69604 4880 69660
rect 4880 69604 4936 69660
rect 4936 69604 4940 69660
rect 4876 69600 4940 69604
rect 4956 69660 5020 69664
rect 4956 69604 4960 69660
rect 4960 69604 5016 69660
rect 5016 69604 5020 69660
rect 4956 69600 5020 69604
rect 5036 69660 5100 69664
rect 5036 69604 5040 69660
rect 5040 69604 5096 69660
rect 5096 69604 5100 69660
rect 5036 69600 5100 69604
rect 5116 69660 5180 69664
rect 5116 69604 5120 69660
rect 5120 69604 5176 69660
rect 5176 69604 5180 69660
rect 5116 69600 5180 69604
rect 35596 69660 35660 69664
rect 35596 69604 35600 69660
rect 35600 69604 35656 69660
rect 35656 69604 35660 69660
rect 35596 69600 35660 69604
rect 35676 69660 35740 69664
rect 35676 69604 35680 69660
rect 35680 69604 35736 69660
rect 35736 69604 35740 69660
rect 35676 69600 35740 69604
rect 35756 69660 35820 69664
rect 35756 69604 35760 69660
rect 35760 69604 35816 69660
rect 35816 69604 35820 69660
rect 35756 69600 35820 69604
rect 35836 69660 35900 69664
rect 35836 69604 35840 69660
rect 35840 69604 35896 69660
rect 35896 69604 35900 69660
rect 35836 69600 35900 69604
rect 66316 69660 66380 69664
rect 66316 69604 66320 69660
rect 66320 69604 66376 69660
rect 66376 69604 66380 69660
rect 66316 69600 66380 69604
rect 66396 69660 66460 69664
rect 66396 69604 66400 69660
rect 66400 69604 66456 69660
rect 66456 69604 66460 69660
rect 66396 69600 66460 69604
rect 66476 69660 66540 69664
rect 66476 69604 66480 69660
rect 66480 69604 66536 69660
rect 66536 69604 66540 69660
rect 66476 69600 66540 69604
rect 66556 69660 66620 69664
rect 66556 69604 66560 69660
rect 66560 69604 66616 69660
rect 66616 69604 66620 69660
rect 66556 69600 66620 69604
rect 97036 69660 97100 69664
rect 97036 69604 97040 69660
rect 97040 69604 97096 69660
rect 97096 69604 97100 69660
rect 97036 69600 97100 69604
rect 97116 69660 97180 69664
rect 97116 69604 97120 69660
rect 97120 69604 97176 69660
rect 97176 69604 97180 69660
rect 97116 69600 97180 69604
rect 97196 69660 97260 69664
rect 97196 69604 97200 69660
rect 97200 69604 97256 69660
rect 97256 69604 97260 69660
rect 97196 69600 97260 69604
rect 97276 69660 97340 69664
rect 97276 69604 97280 69660
rect 97280 69604 97336 69660
rect 97336 69604 97340 69660
rect 97276 69600 97340 69604
rect 61148 69260 61212 69324
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 96376 69116 96440 69120
rect 96376 69060 96380 69116
rect 96380 69060 96436 69116
rect 96436 69060 96440 69116
rect 96376 69056 96440 69060
rect 96456 69116 96520 69120
rect 96456 69060 96460 69116
rect 96460 69060 96516 69116
rect 96516 69060 96520 69116
rect 96456 69056 96520 69060
rect 96536 69116 96600 69120
rect 96536 69060 96540 69116
rect 96540 69060 96596 69116
rect 96596 69060 96600 69116
rect 96536 69056 96600 69060
rect 96616 69116 96680 69120
rect 96616 69060 96620 69116
rect 96620 69060 96676 69116
rect 96676 69060 96680 69116
rect 96616 69056 96680 69060
rect 102732 68852 102796 68916
rect 53604 68716 53668 68780
rect 56180 68580 56244 68644
rect 4876 68572 4940 68576
rect 4876 68516 4880 68572
rect 4880 68516 4936 68572
rect 4936 68516 4940 68572
rect 4876 68512 4940 68516
rect 4956 68572 5020 68576
rect 4956 68516 4960 68572
rect 4960 68516 5016 68572
rect 5016 68516 5020 68572
rect 4956 68512 5020 68516
rect 5036 68572 5100 68576
rect 5036 68516 5040 68572
rect 5040 68516 5096 68572
rect 5096 68516 5100 68572
rect 5036 68512 5100 68516
rect 5116 68572 5180 68576
rect 5116 68516 5120 68572
rect 5120 68516 5176 68572
rect 5176 68516 5180 68572
rect 5116 68512 5180 68516
rect 35596 68572 35660 68576
rect 35596 68516 35600 68572
rect 35600 68516 35656 68572
rect 35656 68516 35660 68572
rect 35596 68512 35660 68516
rect 35676 68572 35740 68576
rect 35676 68516 35680 68572
rect 35680 68516 35736 68572
rect 35736 68516 35740 68572
rect 35676 68512 35740 68516
rect 35756 68572 35820 68576
rect 35756 68516 35760 68572
rect 35760 68516 35816 68572
rect 35816 68516 35820 68572
rect 35756 68512 35820 68516
rect 35836 68572 35900 68576
rect 35836 68516 35840 68572
rect 35840 68516 35896 68572
rect 35896 68516 35900 68572
rect 35836 68512 35900 68516
rect 66316 68572 66380 68576
rect 66316 68516 66320 68572
rect 66320 68516 66376 68572
rect 66376 68516 66380 68572
rect 66316 68512 66380 68516
rect 66396 68572 66460 68576
rect 66396 68516 66400 68572
rect 66400 68516 66456 68572
rect 66456 68516 66460 68572
rect 66396 68512 66460 68516
rect 66476 68572 66540 68576
rect 66476 68516 66480 68572
rect 66480 68516 66536 68572
rect 66536 68516 66540 68572
rect 66476 68512 66540 68516
rect 66556 68572 66620 68576
rect 66556 68516 66560 68572
rect 66560 68516 66616 68572
rect 66616 68516 66620 68572
rect 66556 68512 66620 68516
rect 97036 68572 97100 68576
rect 97036 68516 97040 68572
rect 97040 68516 97096 68572
rect 97096 68516 97100 68572
rect 97036 68512 97100 68516
rect 97116 68572 97180 68576
rect 97116 68516 97120 68572
rect 97120 68516 97176 68572
rect 97176 68516 97180 68572
rect 97116 68512 97180 68516
rect 97196 68572 97260 68576
rect 97196 68516 97200 68572
rect 97200 68516 97256 68572
rect 97256 68516 97260 68572
rect 97196 68512 97260 68516
rect 97276 68572 97340 68576
rect 97276 68516 97280 68572
rect 97280 68516 97336 68572
rect 97336 68516 97340 68572
rect 97276 68512 97340 68516
rect 48636 68172 48700 68236
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 96376 68028 96440 68032
rect 96376 67972 96380 68028
rect 96380 67972 96436 68028
rect 96436 67972 96440 68028
rect 96376 67968 96440 67972
rect 96456 68028 96520 68032
rect 96456 67972 96460 68028
rect 96460 67972 96516 68028
rect 96516 67972 96520 68028
rect 96456 67968 96520 67972
rect 96536 68028 96600 68032
rect 96536 67972 96540 68028
rect 96540 67972 96596 68028
rect 96596 67972 96600 68028
rect 96536 67968 96600 67972
rect 96616 68028 96680 68032
rect 96616 67972 96620 68028
rect 96620 67972 96676 68028
rect 96676 67972 96680 68028
rect 96616 67968 96680 67972
rect 4876 67484 4940 67488
rect 4876 67428 4880 67484
rect 4880 67428 4936 67484
rect 4936 67428 4940 67484
rect 4876 67424 4940 67428
rect 4956 67484 5020 67488
rect 4956 67428 4960 67484
rect 4960 67428 5016 67484
rect 5016 67428 5020 67484
rect 4956 67424 5020 67428
rect 5036 67484 5100 67488
rect 5036 67428 5040 67484
rect 5040 67428 5096 67484
rect 5096 67428 5100 67484
rect 5036 67424 5100 67428
rect 5116 67484 5180 67488
rect 5116 67428 5120 67484
rect 5120 67428 5176 67484
rect 5176 67428 5180 67484
rect 5116 67424 5180 67428
rect 35596 67484 35660 67488
rect 35596 67428 35600 67484
rect 35600 67428 35656 67484
rect 35656 67428 35660 67484
rect 35596 67424 35660 67428
rect 35676 67484 35740 67488
rect 35676 67428 35680 67484
rect 35680 67428 35736 67484
rect 35736 67428 35740 67484
rect 35676 67424 35740 67428
rect 35756 67484 35820 67488
rect 35756 67428 35760 67484
rect 35760 67428 35816 67484
rect 35816 67428 35820 67484
rect 35756 67424 35820 67428
rect 35836 67484 35900 67488
rect 35836 67428 35840 67484
rect 35840 67428 35896 67484
rect 35896 67428 35900 67484
rect 35836 67424 35900 67428
rect 66316 67484 66380 67488
rect 66316 67428 66320 67484
rect 66320 67428 66376 67484
rect 66376 67428 66380 67484
rect 66316 67424 66380 67428
rect 66396 67484 66460 67488
rect 66396 67428 66400 67484
rect 66400 67428 66456 67484
rect 66456 67428 66460 67484
rect 66396 67424 66460 67428
rect 66476 67484 66540 67488
rect 66476 67428 66480 67484
rect 66480 67428 66536 67484
rect 66536 67428 66540 67484
rect 66476 67424 66540 67428
rect 66556 67484 66620 67488
rect 66556 67428 66560 67484
rect 66560 67428 66616 67484
rect 66616 67428 66620 67484
rect 66556 67424 66620 67428
rect 97036 67484 97100 67488
rect 97036 67428 97040 67484
rect 97040 67428 97096 67484
rect 97096 67428 97100 67484
rect 97036 67424 97100 67428
rect 97116 67484 97180 67488
rect 97116 67428 97120 67484
rect 97120 67428 97176 67484
rect 97176 67428 97180 67484
rect 97116 67424 97180 67428
rect 97196 67484 97260 67488
rect 97196 67428 97200 67484
rect 97200 67428 97256 67484
rect 97256 67428 97260 67484
rect 97196 67424 97260 67428
rect 97276 67484 97340 67488
rect 97276 67428 97280 67484
rect 97280 67428 97336 67484
rect 97336 67428 97340 67484
rect 97276 67424 97340 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 96376 66940 96440 66944
rect 96376 66884 96380 66940
rect 96380 66884 96436 66940
rect 96436 66884 96440 66940
rect 96376 66880 96440 66884
rect 96456 66940 96520 66944
rect 96456 66884 96460 66940
rect 96460 66884 96516 66940
rect 96516 66884 96520 66940
rect 96456 66880 96520 66884
rect 96536 66940 96600 66944
rect 96536 66884 96540 66940
rect 96540 66884 96596 66940
rect 96596 66884 96600 66940
rect 96536 66880 96600 66884
rect 96616 66940 96680 66944
rect 96616 66884 96620 66940
rect 96620 66884 96676 66940
rect 96676 66884 96680 66940
rect 96616 66880 96680 66884
rect 4876 66396 4940 66400
rect 4876 66340 4880 66396
rect 4880 66340 4936 66396
rect 4936 66340 4940 66396
rect 4876 66336 4940 66340
rect 4956 66396 5020 66400
rect 4956 66340 4960 66396
rect 4960 66340 5016 66396
rect 5016 66340 5020 66396
rect 4956 66336 5020 66340
rect 5036 66396 5100 66400
rect 5036 66340 5040 66396
rect 5040 66340 5096 66396
rect 5096 66340 5100 66396
rect 5036 66336 5100 66340
rect 5116 66396 5180 66400
rect 5116 66340 5120 66396
rect 5120 66340 5176 66396
rect 5176 66340 5180 66396
rect 5116 66336 5180 66340
rect 35596 66396 35660 66400
rect 35596 66340 35600 66396
rect 35600 66340 35656 66396
rect 35656 66340 35660 66396
rect 35596 66336 35660 66340
rect 35676 66396 35740 66400
rect 35676 66340 35680 66396
rect 35680 66340 35736 66396
rect 35736 66340 35740 66396
rect 35676 66336 35740 66340
rect 35756 66396 35820 66400
rect 35756 66340 35760 66396
rect 35760 66340 35816 66396
rect 35816 66340 35820 66396
rect 35756 66336 35820 66340
rect 35836 66396 35900 66400
rect 35836 66340 35840 66396
rect 35840 66340 35896 66396
rect 35896 66340 35900 66396
rect 35836 66336 35900 66340
rect 66316 66396 66380 66400
rect 66316 66340 66320 66396
rect 66320 66340 66376 66396
rect 66376 66340 66380 66396
rect 66316 66336 66380 66340
rect 66396 66396 66460 66400
rect 66396 66340 66400 66396
rect 66400 66340 66456 66396
rect 66456 66340 66460 66396
rect 66396 66336 66460 66340
rect 66476 66396 66540 66400
rect 66476 66340 66480 66396
rect 66480 66340 66536 66396
rect 66536 66340 66540 66396
rect 66476 66336 66540 66340
rect 66556 66396 66620 66400
rect 66556 66340 66560 66396
rect 66560 66340 66616 66396
rect 66616 66340 66620 66396
rect 66556 66336 66620 66340
rect 97036 66396 97100 66400
rect 97036 66340 97040 66396
rect 97040 66340 97096 66396
rect 97096 66340 97100 66396
rect 97036 66336 97100 66340
rect 97116 66396 97180 66400
rect 97116 66340 97120 66396
rect 97120 66340 97176 66396
rect 97176 66340 97180 66396
rect 97116 66336 97180 66340
rect 97196 66396 97260 66400
rect 97196 66340 97200 66396
rect 97200 66340 97256 66396
rect 97256 66340 97260 66396
rect 97196 66336 97260 66340
rect 97276 66396 97340 66400
rect 97276 66340 97280 66396
rect 97280 66340 97336 66396
rect 97336 66340 97340 66396
rect 97276 66336 97340 66340
rect 106660 66396 106724 66400
rect 106660 66340 106664 66396
rect 106664 66340 106720 66396
rect 106720 66340 106724 66396
rect 106660 66336 106724 66340
rect 106740 66396 106804 66400
rect 106740 66340 106744 66396
rect 106744 66340 106800 66396
rect 106800 66340 106804 66396
rect 106740 66336 106804 66340
rect 106820 66396 106884 66400
rect 106820 66340 106824 66396
rect 106824 66340 106880 66396
rect 106880 66340 106884 66396
rect 106820 66336 106884 66340
rect 106900 66396 106964 66400
rect 106900 66340 106904 66396
rect 106904 66340 106960 66396
rect 106960 66340 106964 66396
rect 106900 66336 106964 66340
rect 68508 66132 68572 66196
rect 87276 65860 87340 65924
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 96376 65852 96440 65856
rect 96376 65796 96380 65852
rect 96380 65796 96436 65852
rect 96436 65796 96440 65852
rect 96376 65792 96440 65796
rect 96456 65852 96520 65856
rect 96456 65796 96460 65852
rect 96460 65796 96516 65852
rect 96516 65796 96520 65852
rect 96456 65792 96520 65796
rect 96536 65852 96600 65856
rect 96536 65796 96540 65852
rect 96540 65796 96596 65852
rect 96596 65796 96600 65852
rect 96536 65792 96600 65796
rect 96616 65852 96680 65856
rect 96616 65796 96620 65852
rect 96620 65796 96676 65852
rect 96676 65796 96680 65852
rect 96616 65792 96680 65796
rect 105924 65852 105988 65856
rect 105924 65796 105928 65852
rect 105928 65796 105984 65852
rect 105984 65796 105988 65852
rect 105924 65792 105988 65796
rect 106004 65852 106068 65856
rect 106004 65796 106008 65852
rect 106008 65796 106064 65852
rect 106064 65796 106068 65852
rect 106004 65792 106068 65796
rect 106084 65852 106148 65856
rect 106084 65796 106088 65852
rect 106088 65796 106144 65852
rect 106144 65796 106148 65852
rect 106084 65792 106148 65796
rect 106164 65852 106228 65856
rect 106164 65796 106168 65852
rect 106168 65796 106224 65852
rect 106224 65796 106228 65852
rect 106164 65792 106228 65796
rect 36124 65588 36188 65652
rect 46060 65588 46124 65652
rect 38516 65452 38580 65516
rect 4876 65308 4940 65312
rect 4876 65252 4880 65308
rect 4880 65252 4936 65308
rect 4936 65252 4940 65308
rect 4876 65248 4940 65252
rect 4956 65308 5020 65312
rect 4956 65252 4960 65308
rect 4960 65252 5016 65308
rect 5016 65252 5020 65308
rect 4956 65248 5020 65252
rect 5036 65308 5100 65312
rect 5036 65252 5040 65308
rect 5040 65252 5096 65308
rect 5096 65252 5100 65308
rect 5036 65248 5100 65252
rect 5116 65308 5180 65312
rect 5116 65252 5120 65308
rect 5120 65252 5176 65308
rect 5176 65252 5180 65308
rect 5116 65248 5180 65252
rect 106660 65308 106724 65312
rect 106660 65252 106664 65308
rect 106664 65252 106720 65308
rect 106720 65252 106724 65308
rect 106660 65248 106724 65252
rect 106740 65308 106804 65312
rect 106740 65252 106744 65308
rect 106744 65252 106800 65308
rect 106800 65252 106804 65308
rect 106740 65248 106804 65252
rect 106820 65308 106884 65312
rect 106820 65252 106824 65308
rect 106824 65252 106880 65308
rect 106880 65252 106884 65308
rect 106820 65248 106884 65252
rect 106900 65308 106964 65312
rect 106900 65252 106904 65308
rect 106904 65252 106960 65308
rect 106960 65252 106964 65308
rect 106900 65248 106964 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 105924 64764 105988 64768
rect 105924 64708 105928 64764
rect 105928 64708 105984 64764
rect 105984 64708 105988 64764
rect 105924 64704 105988 64708
rect 106004 64764 106068 64768
rect 106004 64708 106008 64764
rect 106008 64708 106064 64764
rect 106064 64708 106068 64764
rect 106004 64704 106068 64708
rect 106084 64764 106148 64768
rect 106084 64708 106088 64764
rect 106088 64708 106144 64764
rect 106144 64708 106148 64764
rect 106084 64704 106148 64708
rect 106164 64764 106228 64768
rect 106164 64708 106168 64764
rect 106168 64708 106224 64764
rect 106224 64708 106228 64764
rect 106164 64704 106228 64708
rect 41092 64288 41156 64292
rect 41092 64232 41142 64288
rect 41142 64232 41156 64288
rect 41092 64228 41156 64232
rect 4876 64220 4940 64224
rect 4876 64164 4880 64220
rect 4880 64164 4936 64220
rect 4936 64164 4940 64220
rect 4876 64160 4940 64164
rect 4956 64220 5020 64224
rect 4956 64164 4960 64220
rect 4960 64164 5016 64220
rect 5016 64164 5020 64220
rect 4956 64160 5020 64164
rect 5036 64220 5100 64224
rect 5036 64164 5040 64220
rect 5040 64164 5096 64220
rect 5096 64164 5100 64220
rect 5036 64160 5100 64164
rect 5116 64220 5180 64224
rect 5116 64164 5120 64220
rect 5120 64164 5176 64220
rect 5176 64164 5180 64220
rect 5116 64160 5180 64164
rect 106660 64220 106724 64224
rect 106660 64164 106664 64220
rect 106664 64164 106720 64220
rect 106720 64164 106724 64220
rect 106660 64160 106724 64164
rect 106740 64220 106804 64224
rect 106740 64164 106744 64220
rect 106744 64164 106800 64220
rect 106800 64164 106804 64220
rect 106740 64160 106804 64164
rect 106820 64220 106884 64224
rect 106820 64164 106824 64220
rect 106824 64164 106880 64220
rect 106880 64164 106884 64220
rect 106820 64160 106884 64164
rect 106900 64220 106964 64224
rect 106900 64164 106904 64220
rect 106904 64164 106960 64220
rect 106960 64164 106964 64220
rect 106900 64160 106964 64164
rect 43563 64092 43627 64156
rect 51051 64092 51115 64156
rect 58539 64092 58603 64156
rect 95858 64152 95922 64156
rect 95858 64096 95882 64152
rect 95882 64096 95922 64152
rect 95858 64092 95922 64096
rect 66027 63956 66091 64020
rect 71019 63820 71083 63884
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 105924 63676 105988 63680
rect 105924 63620 105928 63676
rect 105928 63620 105984 63676
rect 105984 63620 105988 63676
rect 105924 63616 105988 63620
rect 106004 63676 106068 63680
rect 106004 63620 106008 63676
rect 106008 63620 106064 63676
rect 106064 63620 106068 63676
rect 106004 63616 106068 63620
rect 106084 63676 106148 63680
rect 106084 63620 106088 63676
rect 106088 63620 106144 63676
rect 106144 63620 106148 63676
rect 106084 63616 106148 63620
rect 106164 63676 106228 63680
rect 106164 63620 106168 63676
rect 106168 63620 106224 63676
rect 106224 63620 106228 63676
rect 106164 63616 106228 63620
rect 4876 63132 4940 63136
rect 4876 63076 4880 63132
rect 4880 63076 4936 63132
rect 4936 63076 4940 63132
rect 4876 63072 4940 63076
rect 4956 63132 5020 63136
rect 4956 63076 4960 63132
rect 4960 63076 5016 63132
rect 5016 63076 5020 63132
rect 4956 63072 5020 63076
rect 5036 63132 5100 63136
rect 5036 63076 5040 63132
rect 5040 63076 5096 63132
rect 5096 63076 5100 63132
rect 5036 63072 5100 63076
rect 5116 63132 5180 63136
rect 5116 63076 5120 63132
rect 5120 63076 5176 63132
rect 5176 63076 5180 63132
rect 5116 63072 5180 63076
rect 106660 63132 106724 63136
rect 106660 63076 106664 63132
rect 106664 63076 106720 63132
rect 106720 63076 106724 63132
rect 106660 63072 106724 63076
rect 106740 63132 106804 63136
rect 106740 63076 106744 63132
rect 106744 63076 106800 63132
rect 106800 63076 106804 63132
rect 106740 63072 106804 63076
rect 106820 63132 106884 63136
rect 106820 63076 106824 63132
rect 106824 63076 106880 63132
rect 106880 63076 106884 63132
rect 106820 63072 106884 63076
rect 106900 63132 106964 63136
rect 106900 63076 106904 63132
rect 106904 63076 106960 63132
rect 106960 63076 106964 63132
rect 106900 63072 106964 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 105924 62588 105988 62592
rect 105924 62532 105928 62588
rect 105928 62532 105984 62588
rect 105984 62532 105988 62588
rect 105924 62528 105988 62532
rect 106004 62588 106068 62592
rect 106004 62532 106008 62588
rect 106008 62532 106064 62588
rect 106064 62532 106068 62588
rect 106004 62528 106068 62532
rect 106084 62588 106148 62592
rect 106084 62532 106088 62588
rect 106088 62532 106144 62588
rect 106144 62532 106148 62588
rect 106084 62528 106148 62532
rect 106164 62588 106228 62592
rect 106164 62532 106168 62588
rect 106168 62532 106224 62588
rect 106224 62532 106228 62588
rect 106164 62528 106228 62532
rect 4876 62044 4940 62048
rect 4876 61988 4880 62044
rect 4880 61988 4936 62044
rect 4936 61988 4940 62044
rect 4876 61984 4940 61988
rect 4956 62044 5020 62048
rect 4956 61988 4960 62044
rect 4960 61988 5016 62044
rect 5016 61988 5020 62044
rect 4956 61984 5020 61988
rect 5036 62044 5100 62048
rect 5036 61988 5040 62044
rect 5040 61988 5096 62044
rect 5096 61988 5100 62044
rect 5036 61984 5100 61988
rect 5116 62044 5180 62048
rect 5116 61988 5120 62044
rect 5120 61988 5176 62044
rect 5176 61988 5180 62044
rect 5116 61984 5180 61988
rect 106660 62044 106724 62048
rect 106660 61988 106664 62044
rect 106664 61988 106720 62044
rect 106720 61988 106724 62044
rect 106660 61984 106724 61988
rect 106740 62044 106804 62048
rect 106740 61988 106744 62044
rect 106744 61988 106800 62044
rect 106800 61988 106804 62044
rect 106740 61984 106804 61988
rect 106820 62044 106884 62048
rect 106820 61988 106824 62044
rect 106824 61988 106880 62044
rect 106880 61988 106884 62044
rect 106820 61984 106884 61988
rect 106900 62044 106964 62048
rect 106900 61988 106904 62044
rect 106904 61988 106960 62044
rect 106960 61988 106964 62044
rect 106900 61984 106964 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 105924 61500 105988 61504
rect 105924 61444 105928 61500
rect 105928 61444 105984 61500
rect 105984 61444 105988 61500
rect 105924 61440 105988 61444
rect 106004 61500 106068 61504
rect 106004 61444 106008 61500
rect 106008 61444 106064 61500
rect 106064 61444 106068 61500
rect 106004 61440 106068 61444
rect 106084 61500 106148 61504
rect 106084 61444 106088 61500
rect 106088 61444 106144 61500
rect 106144 61444 106148 61500
rect 106084 61440 106148 61444
rect 106164 61500 106228 61504
rect 106164 61444 106168 61500
rect 106168 61444 106224 61500
rect 106224 61444 106228 61500
rect 106164 61440 106228 61444
rect 4876 60956 4940 60960
rect 4876 60900 4880 60956
rect 4880 60900 4936 60956
rect 4936 60900 4940 60956
rect 4876 60896 4940 60900
rect 4956 60956 5020 60960
rect 4956 60900 4960 60956
rect 4960 60900 5016 60956
rect 5016 60900 5020 60956
rect 4956 60896 5020 60900
rect 5036 60956 5100 60960
rect 5036 60900 5040 60956
rect 5040 60900 5096 60956
rect 5096 60900 5100 60956
rect 5036 60896 5100 60900
rect 5116 60956 5180 60960
rect 5116 60900 5120 60956
rect 5120 60900 5176 60956
rect 5176 60900 5180 60956
rect 5116 60896 5180 60900
rect 106660 60956 106724 60960
rect 106660 60900 106664 60956
rect 106664 60900 106720 60956
rect 106720 60900 106724 60956
rect 106660 60896 106724 60900
rect 106740 60956 106804 60960
rect 106740 60900 106744 60956
rect 106744 60900 106800 60956
rect 106800 60900 106804 60956
rect 106740 60896 106804 60900
rect 106820 60956 106884 60960
rect 106820 60900 106824 60956
rect 106824 60900 106880 60956
rect 106880 60900 106884 60956
rect 106820 60896 106884 60900
rect 106900 60956 106964 60960
rect 106900 60900 106904 60956
rect 106904 60900 106960 60956
rect 106960 60900 106964 60956
rect 106900 60896 106964 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 105924 60412 105988 60416
rect 105924 60356 105928 60412
rect 105928 60356 105984 60412
rect 105984 60356 105988 60412
rect 105924 60352 105988 60356
rect 106004 60412 106068 60416
rect 106004 60356 106008 60412
rect 106008 60356 106064 60412
rect 106064 60356 106068 60412
rect 106004 60352 106068 60356
rect 106084 60412 106148 60416
rect 106084 60356 106088 60412
rect 106088 60356 106144 60412
rect 106144 60356 106148 60412
rect 106084 60352 106148 60356
rect 106164 60412 106228 60416
rect 106164 60356 106168 60412
rect 106168 60356 106224 60412
rect 106224 60356 106228 60412
rect 106164 60352 106228 60356
rect 4876 59868 4940 59872
rect 4876 59812 4880 59868
rect 4880 59812 4936 59868
rect 4936 59812 4940 59868
rect 4876 59808 4940 59812
rect 4956 59868 5020 59872
rect 4956 59812 4960 59868
rect 4960 59812 5016 59868
rect 5016 59812 5020 59868
rect 4956 59808 5020 59812
rect 5036 59868 5100 59872
rect 5036 59812 5040 59868
rect 5040 59812 5096 59868
rect 5096 59812 5100 59868
rect 5036 59808 5100 59812
rect 5116 59868 5180 59872
rect 5116 59812 5120 59868
rect 5120 59812 5176 59868
rect 5176 59812 5180 59868
rect 5116 59808 5180 59812
rect 106660 59868 106724 59872
rect 106660 59812 106664 59868
rect 106664 59812 106720 59868
rect 106720 59812 106724 59868
rect 106660 59808 106724 59812
rect 106740 59868 106804 59872
rect 106740 59812 106744 59868
rect 106744 59812 106800 59868
rect 106800 59812 106804 59868
rect 106740 59808 106804 59812
rect 106820 59868 106884 59872
rect 106820 59812 106824 59868
rect 106824 59812 106880 59868
rect 106880 59812 106884 59868
rect 106820 59808 106884 59812
rect 106900 59868 106964 59872
rect 106900 59812 106904 59868
rect 106904 59812 106960 59868
rect 106960 59812 106964 59868
rect 106900 59808 106964 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 105924 59324 105988 59328
rect 105924 59268 105928 59324
rect 105928 59268 105984 59324
rect 105984 59268 105988 59324
rect 105924 59264 105988 59268
rect 106004 59324 106068 59328
rect 106004 59268 106008 59324
rect 106008 59268 106064 59324
rect 106064 59268 106068 59324
rect 106004 59264 106068 59268
rect 106084 59324 106148 59328
rect 106084 59268 106088 59324
rect 106088 59268 106144 59324
rect 106144 59268 106148 59324
rect 106084 59264 106148 59268
rect 106164 59324 106228 59328
rect 106164 59268 106168 59324
rect 106168 59268 106224 59324
rect 106224 59268 106228 59324
rect 106164 59264 106228 59268
rect 4876 58780 4940 58784
rect 4876 58724 4880 58780
rect 4880 58724 4936 58780
rect 4936 58724 4940 58780
rect 4876 58720 4940 58724
rect 4956 58780 5020 58784
rect 4956 58724 4960 58780
rect 4960 58724 5016 58780
rect 5016 58724 5020 58780
rect 4956 58720 5020 58724
rect 5036 58780 5100 58784
rect 5036 58724 5040 58780
rect 5040 58724 5096 58780
rect 5096 58724 5100 58780
rect 5036 58720 5100 58724
rect 5116 58780 5180 58784
rect 5116 58724 5120 58780
rect 5120 58724 5176 58780
rect 5176 58724 5180 58780
rect 5116 58720 5180 58724
rect 106660 58780 106724 58784
rect 106660 58724 106664 58780
rect 106664 58724 106720 58780
rect 106720 58724 106724 58780
rect 106660 58720 106724 58724
rect 106740 58780 106804 58784
rect 106740 58724 106744 58780
rect 106744 58724 106800 58780
rect 106800 58724 106804 58780
rect 106740 58720 106804 58724
rect 106820 58780 106884 58784
rect 106820 58724 106824 58780
rect 106824 58724 106880 58780
rect 106880 58724 106884 58780
rect 106820 58720 106884 58724
rect 106900 58780 106964 58784
rect 106900 58724 106904 58780
rect 106904 58724 106960 58780
rect 106960 58724 106964 58780
rect 106900 58720 106964 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 105924 58236 105988 58240
rect 105924 58180 105928 58236
rect 105928 58180 105984 58236
rect 105984 58180 105988 58236
rect 105924 58176 105988 58180
rect 106004 58236 106068 58240
rect 106004 58180 106008 58236
rect 106008 58180 106064 58236
rect 106064 58180 106068 58236
rect 106004 58176 106068 58180
rect 106084 58236 106148 58240
rect 106084 58180 106088 58236
rect 106088 58180 106144 58236
rect 106144 58180 106148 58236
rect 106084 58176 106148 58180
rect 106164 58236 106228 58240
rect 106164 58180 106168 58236
rect 106168 58180 106224 58236
rect 106224 58180 106228 58236
rect 106164 58176 106228 58180
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 106660 57692 106724 57696
rect 106660 57636 106664 57692
rect 106664 57636 106720 57692
rect 106720 57636 106724 57692
rect 106660 57632 106724 57636
rect 106740 57692 106804 57696
rect 106740 57636 106744 57692
rect 106744 57636 106800 57692
rect 106800 57636 106804 57692
rect 106740 57632 106804 57636
rect 106820 57692 106884 57696
rect 106820 57636 106824 57692
rect 106824 57636 106880 57692
rect 106880 57636 106884 57692
rect 106820 57632 106884 57636
rect 106900 57692 106964 57696
rect 106900 57636 106904 57692
rect 106904 57636 106960 57692
rect 106960 57636 106964 57692
rect 106900 57632 106964 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 105924 57148 105988 57152
rect 105924 57092 105928 57148
rect 105928 57092 105984 57148
rect 105984 57092 105988 57148
rect 105924 57088 105988 57092
rect 106004 57148 106068 57152
rect 106004 57092 106008 57148
rect 106008 57092 106064 57148
rect 106064 57092 106068 57148
rect 106004 57088 106068 57092
rect 106084 57148 106148 57152
rect 106084 57092 106088 57148
rect 106088 57092 106144 57148
rect 106144 57092 106148 57148
rect 106084 57088 106148 57092
rect 106164 57148 106228 57152
rect 106164 57092 106168 57148
rect 106168 57092 106224 57148
rect 106224 57092 106228 57148
rect 106164 57088 106228 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 106660 56604 106724 56608
rect 106660 56548 106664 56604
rect 106664 56548 106720 56604
rect 106720 56548 106724 56604
rect 106660 56544 106724 56548
rect 106740 56604 106804 56608
rect 106740 56548 106744 56604
rect 106744 56548 106800 56604
rect 106800 56548 106804 56604
rect 106740 56544 106804 56548
rect 106820 56604 106884 56608
rect 106820 56548 106824 56604
rect 106824 56548 106880 56604
rect 106880 56548 106884 56604
rect 106820 56544 106884 56548
rect 106900 56604 106964 56608
rect 106900 56548 106904 56604
rect 106904 56548 106960 56604
rect 106960 56548 106964 56604
rect 106900 56544 106964 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 105924 56060 105988 56064
rect 105924 56004 105928 56060
rect 105928 56004 105984 56060
rect 105984 56004 105988 56060
rect 105924 56000 105988 56004
rect 106004 56060 106068 56064
rect 106004 56004 106008 56060
rect 106008 56004 106064 56060
rect 106064 56004 106068 56060
rect 106004 56000 106068 56004
rect 106084 56060 106148 56064
rect 106084 56004 106088 56060
rect 106088 56004 106144 56060
rect 106144 56004 106148 56060
rect 106084 56000 106148 56004
rect 106164 56060 106228 56064
rect 106164 56004 106168 56060
rect 106168 56004 106224 56060
rect 106224 56004 106228 56060
rect 106164 56000 106228 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 106660 55516 106724 55520
rect 106660 55460 106664 55516
rect 106664 55460 106720 55516
rect 106720 55460 106724 55516
rect 106660 55456 106724 55460
rect 106740 55516 106804 55520
rect 106740 55460 106744 55516
rect 106744 55460 106800 55516
rect 106800 55460 106804 55516
rect 106740 55456 106804 55460
rect 106820 55516 106884 55520
rect 106820 55460 106824 55516
rect 106824 55460 106880 55516
rect 106880 55460 106884 55516
rect 106820 55456 106884 55460
rect 106900 55516 106964 55520
rect 106900 55460 106904 55516
rect 106904 55460 106960 55516
rect 106960 55460 106964 55516
rect 106900 55456 106964 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 105924 54972 105988 54976
rect 105924 54916 105928 54972
rect 105928 54916 105984 54972
rect 105984 54916 105988 54972
rect 105924 54912 105988 54916
rect 106004 54972 106068 54976
rect 106004 54916 106008 54972
rect 106008 54916 106064 54972
rect 106064 54916 106068 54972
rect 106004 54912 106068 54916
rect 106084 54972 106148 54976
rect 106084 54916 106088 54972
rect 106088 54916 106144 54972
rect 106144 54916 106148 54972
rect 106084 54912 106148 54916
rect 106164 54972 106228 54976
rect 106164 54916 106168 54972
rect 106168 54916 106224 54972
rect 106224 54916 106228 54972
rect 106164 54912 106228 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 106660 54428 106724 54432
rect 106660 54372 106664 54428
rect 106664 54372 106720 54428
rect 106720 54372 106724 54428
rect 106660 54368 106724 54372
rect 106740 54428 106804 54432
rect 106740 54372 106744 54428
rect 106744 54372 106800 54428
rect 106800 54372 106804 54428
rect 106740 54368 106804 54372
rect 106820 54428 106884 54432
rect 106820 54372 106824 54428
rect 106824 54372 106880 54428
rect 106880 54372 106884 54428
rect 106820 54368 106884 54372
rect 106900 54428 106964 54432
rect 106900 54372 106904 54428
rect 106904 54372 106960 54428
rect 106960 54372 106964 54428
rect 106900 54368 106964 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 105924 53884 105988 53888
rect 105924 53828 105928 53884
rect 105928 53828 105984 53884
rect 105984 53828 105988 53884
rect 105924 53824 105988 53828
rect 106004 53884 106068 53888
rect 106004 53828 106008 53884
rect 106008 53828 106064 53884
rect 106064 53828 106068 53884
rect 106004 53824 106068 53828
rect 106084 53884 106148 53888
rect 106084 53828 106088 53884
rect 106088 53828 106144 53884
rect 106144 53828 106148 53884
rect 106084 53824 106148 53828
rect 106164 53884 106228 53888
rect 106164 53828 106168 53884
rect 106168 53828 106224 53884
rect 106224 53828 106228 53884
rect 106164 53824 106228 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 106660 53340 106724 53344
rect 106660 53284 106664 53340
rect 106664 53284 106720 53340
rect 106720 53284 106724 53340
rect 106660 53280 106724 53284
rect 106740 53340 106804 53344
rect 106740 53284 106744 53340
rect 106744 53284 106800 53340
rect 106800 53284 106804 53340
rect 106740 53280 106804 53284
rect 106820 53340 106884 53344
rect 106820 53284 106824 53340
rect 106824 53284 106880 53340
rect 106880 53284 106884 53340
rect 106820 53280 106884 53284
rect 106900 53340 106964 53344
rect 106900 53284 106904 53340
rect 106904 53284 106960 53340
rect 106960 53284 106964 53340
rect 106900 53280 106964 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 105924 52796 105988 52800
rect 105924 52740 105928 52796
rect 105928 52740 105984 52796
rect 105984 52740 105988 52796
rect 105924 52736 105988 52740
rect 106004 52796 106068 52800
rect 106004 52740 106008 52796
rect 106008 52740 106064 52796
rect 106064 52740 106068 52796
rect 106004 52736 106068 52740
rect 106084 52796 106148 52800
rect 106084 52740 106088 52796
rect 106088 52740 106144 52796
rect 106144 52740 106148 52796
rect 106084 52736 106148 52740
rect 106164 52796 106228 52800
rect 106164 52740 106168 52796
rect 106168 52740 106224 52796
rect 106224 52740 106228 52796
rect 106164 52736 106228 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 106660 52252 106724 52256
rect 106660 52196 106664 52252
rect 106664 52196 106720 52252
rect 106720 52196 106724 52252
rect 106660 52192 106724 52196
rect 106740 52252 106804 52256
rect 106740 52196 106744 52252
rect 106744 52196 106800 52252
rect 106800 52196 106804 52252
rect 106740 52192 106804 52196
rect 106820 52252 106884 52256
rect 106820 52196 106824 52252
rect 106824 52196 106880 52252
rect 106880 52196 106884 52252
rect 106820 52192 106884 52196
rect 106900 52252 106964 52256
rect 106900 52196 106904 52252
rect 106904 52196 106960 52252
rect 106960 52196 106964 52252
rect 106900 52192 106964 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 105924 51708 105988 51712
rect 105924 51652 105928 51708
rect 105928 51652 105984 51708
rect 105984 51652 105988 51708
rect 105924 51648 105988 51652
rect 106004 51708 106068 51712
rect 106004 51652 106008 51708
rect 106008 51652 106064 51708
rect 106064 51652 106068 51708
rect 106004 51648 106068 51652
rect 106084 51708 106148 51712
rect 106084 51652 106088 51708
rect 106088 51652 106144 51708
rect 106144 51652 106148 51708
rect 106084 51648 106148 51652
rect 106164 51708 106228 51712
rect 106164 51652 106168 51708
rect 106168 51652 106224 51708
rect 106224 51652 106228 51708
rect 106164 51648 106228 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 106660 51164 106724 51168
rect 106660 51108 106664 51164
rect 106664 51108 106720 51164
rect 106720 51108 106724 51164
rect 106660 51104 106724 51108
rect 106740 51164 106804 51168
rect 106740 51108 106744 51164
rect 106744 51108 106800 51164
rect 106800 51108 106804 51164
rect 106740 51104 106804 51108
rect 106820 51164 106884 51168
rect 106820 51108 106824 51164
rect 106824 51108 106880 51164
rect 106880 51108 106884 51164
rect 106820 51104 106884 51108
rect 106900 51164 106964 51168
rect 106900 51108 106904 51164
rect 106904 51108 106960 51164
rect 106960 51108 106964 51164
rect 106900 51104 106964 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 105924 50620 105988 50624
rect 105924 50564 105928 50620
rect 105928 50564 105984 50620
rect 105984 50564 105988 50620
rect 105924 50560 105988 50564
rect 106004 50620 106068 50624
rect 106004 50564 106008 50620
rect 106008 50564 106064 50620
rect 106064 50564 106068 50620
rect 106004 50560 106068 50564
rect 106084 50620 106148 50624
rect 106084 50564 106088 50620
rect 106088 50564 106144 50620
rect 106144 50564 106148 50620
rect 106084 50560 106148 50564
rect 106164 50620 106228 50624
rect 106164 50564 106168 50620
rect 106168 50564 106224 50620
rect 106224 50564 106228 50620
rect 106164 50560 106228 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 106660 50076 106724 50080
rect 106660 50020 106664 50076
rect 106664 50020 106720 50076
rect 106720 50020 106724 50076
rect 106660 50016 106724 50020
rect 106740 50076 106804 50080
rect 106740 50020 106744 50076
rect 106744 50020 106800 50076
rect 106800 50020 106804 50076
rect 106740 50016 106804 50020
rect 106820 50076 106884 50080
rect 106820 50020 106824 50076
rect 106824 50020 106880 50076
rect 106880 50020 106884 50076
rect 106820 50016 106884 50020
rect 106900 50076 106964 50080
rect 106900 50020 106904 50076
rect 106904 50020 106960 50076
rect 106960 50020 106964 50076
rect 106900 50016 106964 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 105924 49532 105988 49536
rect 105924 49476 105928 49532
rect 105928 49476 105984 49532
rect 105984 49476 105988 49532
rect 105924 49472 105988 49476
rect 106004 49532 106068 49536
rect 106004 49476 106008 49532
rect 106008 49476 106064 49532
rect 106064 49476 106068 49532
rect 106004 49472 106068 49476
rect 106084 49532 106148 49536
rect 106084 49476 106088 49532
rect 106088 49476 106144 49532
rect 106144 49476 106148 49532
rect 106084 49472 106148 49476
rect 106164 49532 106228 49536
rect 106164 49476 106168 49532
rect 106168 49476 106224 49532
rect 106224 49476 106228 49532
rect 106164 49472 106228 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 106660 48988 106724 48992
rect 106660 48932 106664 48988
rect 106664 48932 106720 48988
rect 106720 48932 106724 48988
rect 106660 48928 106724 48932
rect 106740 48988 106804 48992
rect 106740 48932 106744 48988
rect 106744 48932 106800 48988
rect 106800 48932 106804 48988
rect 106740 48928 106804 48932
rect 106820 48988 106884 48992
rect 106820 48932 106824 48988
rect 106824 48932 106880 48988
rect 106880 48932 106884 48988
rect 106820 48928 106884 48932
rect 106900 48988 106964 48992
rect 106900 48932 106904 48988
rect 106904 48932 106960 48988
rect 106960 48932 106964 48988
rect 106900 48928 106964 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 105924 48444 105988 48448
rect 105924 48388 105928 48444
rect 105928 48388 105984 48444
rect 105984 48388 105988 48444
rect 105924 48384 105988 48388
rect 106004 48444 106068 48448
rect 106004 48388 106008 48444
rect 106008 48388 106064 48444
rect 106064 48388 106068 48444
rect 106004 48384 106068 48388
rect 106084 48444 106148 48448
rect 106084 48388 106088 48444
rect 106088 48388 106144 48444
rect 106144 48388 106148 48444
rect 106084 48384 106148 48388
rect 106164 48444 106228 48448
rect 106164 48388 106168 48444
rect 106168 48388 106224 48444
rect 106224 48388 106228 48444
rect 106164 48384 106228 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 106660 47900 106724 47904
rect 106660 47844 106664 47900
rect 106664 47844 106720 47900
rect 106720 47844 106724 47900
rect 106660 47840 106724 47844
rect 106740 47900 106804 47904
rect 106740 47844 106744 47900
rect 106744 47844 106800 47900
rect 106800 47844 106804 47900
rect 106740 47840 106804 47844
rect 106820 47900 106884 47904
rect 106820 47844 106824 47900
rect 106824 47844 106880 47900
rect 106880 47844 106884 47900
rect 106820 47840 106884 47844
rect 106900 47900 106964 47904
rect 106900 47844 106904 47900
rect 106904 47844 106960 47900
rect 106960 47844 106964 47900
rect 106900 47840 106964 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 105924 47356 105988 47360
rect 105924 47300 105928 47356
rect 105928 47300 105984 47356
rect 105984 47300 105988 47356
rect 105924 47296 105988 47300
rect 106004 47356 106068 47360
rect 106004 47300 106008 47356
rect 106008 47300 106064 47356
rect 106064 47300 106068 47356
rect 106004 47296 106068 47300
rect 106084 47356 106148 47360
rect 106084 47300 106088 47356
rect 106088 47300 106144 47356
rect 106144 47300 106148 47356
rect 106084 47296 106148 47300
rect 106164 47356 106228 47360
rect 106164 47300 106168 47356
rect 106168 47300 106224 47356
rect 106224 47300 106228 47356
rect 106164 47296 106228 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 106660 46812 106724 46816
rect 106660 46756 106664 46812
rect 106664 46756 106720 46812
rect 106720 46756 106724 46812
rect 106660 46752 106724 46756
rect 106740 46812 106804 46816
rect 106740 46756 106744 46812
rect 106744 46756 106800 46812
rect 106800 46756 106804 46812
rect 106740 46752 106804 46756
rect 106820 46812 106884 46816
rect 106820 46756 106824 46812
rect 106824 46756 106880 46812
rect 106880 46756 106884 46812
rect 106820 46752 106884 46756
rect 106900 46812 106964 46816
rect 106900 46756 106904 46812
rect 106904 46756 106960 46812
rect 106960 46756 106964 46812
rect 106900 46752 106964 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 105924 46268 105988 46272
rect 105924 46212 105928 46268
rect 105928 46212 105984 46268
rect 105984 46212 105988 46268
rect 105924 46208 105988 46212
rect 106004 46268 106068 46272
rect 106004 46212 106008 46268
rect 106008 46212 106064 46268
rect 106064 46212 106068 46268
rect 106004 46208 106068 46212
rect 106084 46268 106148 46272
rect 106084 46212 106088 46268
rect 106088 46212 106144 46268
rect 106144 46212 106148 46268
rect 106084 46208 106148 46212
rect 106164 46268 106228 46272
rect 106164 46212 106168 46268
rect 106168 46212 106224 46268
rect 106224 46212 106228 46268
rect 106164 46208 106228 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 106660 45724 106724 45728
rect 106660 45668 106664 45724
rect 106664 45668 106720 45724
rect 106720 45668 106724 45724
rect 106660 45664 106724 45668
rect 106740 45724 106804 45728
rect 106740 45668 106744 45724
rect 106744 45668 106800 45724
rect 106800 45668 106804 45724
rect 106740 45664 106804 45668
rect 106820 45724 106884 45728
rect 106820 45668 106824 45724
rect 106824 45668 106880 45724
rect 106880 45668 106884 45724
rect 106820 45664 106884 45668
rect 106900 45724 106964 45728
rect 106900 45668 106904 45724
rect 106904 45668 106960 45724
rect 106960 45668 106964 45724
rect 106900 45664 106964 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 105924 45180 105988 45184
rect 105924 45124 105928 45180
rect 105928 45124 105984 45180
rect 105984 45124 105988 45180
rect 105924 45120 105988 45124
rect 106004 45180 106068 45184
rect 106004 45124 106008 45180
rect 106008 45124 106064 45180
rect 106064 45124 106068 45180
rect 106004 45120 106068 45124
rect 106084 45180 106148 45184
rect 106084 45124 106088 45180
rect 106088 45124 106144 45180
rect 106144 45124 106148 45180
rect 106084 45120 106148 45124
rect 106164 45180 106228 45184
rect 106164 45124 106168 45180
rect 106168 45124 106224 45180
rect 106224 45124 106228 45180
rect 106164 45120 106228 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 106660 44636 106724 44640
rect 106660 44580 106664 44636
rect 106664 44580 106720 44636
rect 106720 44580 106724 44636
rect 106660 44576 106724 44580
rect 106740 44636 106804 44640
rect 106740 44580 106744 44636
rect 106744 44580 106800 44636
rect 106800 44580 106804 44636
rect 106740 44576 106804 44580
rect 106820 44636 106884 44640
rect 106820 44580 106824 44636
rect 106824 44580 106880 44636
rect 106880 44580 106884 44636
rect 106820 44576 106884 44580
rect 106900 44636 106964 44640
rect 106900 44580 106904 44636
rect 106904 44580 106960 44636
rect 106960 44580 106964 44636
rect 106900 44576 106964 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 105924 44092 105988 44096
rect 105924 44036 105928 44092
rect 105928 44036 105984 44092
rect 105984 44036 105988 44092
rect 105924 44032 105988 44036
rect 106004 44092 106068 44096
rect 106004 44036 106008 44092
rect 106008 44036 106064 44092
rect 106064 44036 106068 44092
rect 106004 44032 106068 44036
rect 106084 44092 106148 44096
rect 106084 44036 106088 44092
rect 106088 44036 106144 44092
rect 106144 44036 106148 44092
rect 106084 44032 106148 44036
rect 106164 44092 106228 44096
rect 106164 44036 106168 44092
rect 106168 44036 106224 44092
rect 106224 44036 106228 44092
rect 106164 44032 106228 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 106660 43548 106724 43552
rect 106660 43492 106664 43548
rect 106664 43492 106720 43548
rect 106720 43492 106724 43548
rect 106660 43488 106724 43492
rect 106740 43548 106804 43552
rect 106740 43492 106744 43548
rect 106744 43492 106800 43548
rect 106800 43492 106804 43548
rect 106740 43488 106804 43492
rect 106820 43548 106884 43552
rect 106820 43492 106824 43548
rect 106824 43492 106880 43548
rect 106880 43492 106884 43548
rect 106820 43488 106884 43492
rect 106900 43548 106964 43552
rect 106900 43492 106904 43548
rect 106904 43492 106960 43548
rect 106960 43492 106964 43548
rect 106900 43488 106964 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 105924 43004 105988 43008
rect 105924 42948 105928 43004
rect 105928 42948 105984 43004
rect 105984 42948 105988 43004
rect 105924 42944 105988 42948
rect 106004 43004 106068 43008
rect 106004 42948 106008 43004
rect 106008 42948 106064 43004
rect 106064 42948 106068 43004
rect 106004 42944 106068 42948
rect 106084 43004 106148 43008
rect 106084 42948 106088 43004
rect 106088 42948 106144 43004
rect 106144 42948 106148 43004
rect 106084 42944 106148 42948
rect 106164 43004 106228 43008
rect 106164 42948 106168 43004
rect 106168 42948 106224 43004
rect 106224 42948 106228 43004
rect 106164 42944 106228 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 106660 42460 106724 42464
rect 106660 42404 106664 42460
rect 106664 42404 106720 42460
rect 106720 42404 106724 42460
rect 106660 42400 106724 42404
rect 106740 42460 106804 42464
rect 106740 42404 106744 42460
rect 106744 42404 106800 42460
rect 106800 42404 106804 42460
rect 106740 42400 106804 42404
rect 106820 42460 106884 42464
rect 106820 42404 106824 42460
rect 106824 42404 106880 42460
rect 106880 42404 106884 42460
rect 106820 42400 106884 42404
rect 106900 42460 106964 42464
rect 106900 42404 106904 42460
rect 106904 42404 106960 42460
rect 106960 42404 106964 42460
rect 106900 42400 106964 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 105924 41916 105988 41920
rect 105924 41860 105928 41916
rect 105928 41860 105984 41916
rect 105984 41860 105988 41916
rect 105924 41856 105988 41860
rect 106004 41916 106068 41920
rect 106004 41860 106008 41916
rect 106008 41860 106064 41916
rect 106064 41860 106068 41916
rect 106004 41856 106068 41860
rect 106084 41916 106148 41920
rect 106084 41860 106088 41916
rect 106088 41860 106144 41916
rect 106144 41860 106148 41916
rect 106084 41856 106148 41860
rect 106164 41916 106228 41920
rect 106164 41860 106168 41916
rect 106168 41860 106224 41916
rect 106224 41860 106228 41916
rect 106164 41856 106228 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 106660 41372 106724 41376
rect 106660 41316 106664 41372
rect 106664 41316 106720 41372
rect 106720 41316 106724 41372
rect 106660 41312 106724 41316
rect 106740 41372 106804 41376
rect 106740 41316 106744 41372
rect 106744 41316 106800 41372
rect 106800 41316 106804 41372
rect 106740 41312 106804 41316
rect 106820 41372 106884 41376
rect 106820 41316 106824 41372
rect 106824 41316 106880 41372
rect 106880 41316 106884 41372
rect 106820 41312 106884 41316
rect 106900 41372 106964 41376
rect 106900 41316 106904 41372
rect 106904 41316 106960 41372
rect 106960 41316 106964 41372
rect 106900 41312 106964 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 105924 40828 105988 40832
rect 105924 40772 105928 40828
rect 105928 40772 105984 40828
rect 105984 40772 105988 40828
rect 105924 40768 105988 40772
rect 106004 40828 106068 40832
rect 106004 40772 106008 40828
rect 106008 40772 106064 40828
rect 106064 40772 106068 40828
rect 106004 40768 106068 40772
rect 106084 40828 106148 40832
rect 106084 40772 106088 40828
rect 106088 40772 106144 40828
rect 106144 40772 106148 40828
rect 106084 40768 106148 40772
rect 106164 40828 106228 40832
rect 106164 40772 106168 40828
rect 106168 40772 106224 40828
rect 106224 40772 106228 40828
rect 106164 40768 106228 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 106660 40284 106724 40288
rect 106660 40228 106664 40284
rect 106664 40228 106720 40284
rect 106720 40228 106724 40284
rect 106660 40224 106724 40228
rect 106740 40284 106804 40288
rect 106740 40228 106744 40284
rect 106744 40228 106800 40284
rect 106800 40228 106804 40284
rect 106740 40224 106804 40228
rect 106820 40284 106884 40288
rect 106820 40228 106824 40284
rect 106824 40228 106880 40284
rect 106880 40228 106884 40284
rect 106820 40224 106884 40228
rect 106900 40284 106964 40288
rect 106900 40228 106904 40284
rect 106904 40228 106960 40284
rect 106960 40228 106964 40284
rect 106900 40224 106964 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 105924 39740 105988 39744
rect 105924 39684 105928 39740
rect 105928 39684 105984 39740
rect 105984 39684 105988 39740
rect 105924 39680 105988 39684
rect 106004 39740 106068 39744
rect 106004 39684 106008 39740
rect 106008 39684 106064 39740
rect 106064 39684 106068 39740
rect 106004 39680 106068 39684
rect 106084 39740 106148 39744
rect 106084 39684 106088 39740
rect 106088 39684 106144 39740
rect 106144 39684 106148 39740
rect 106084 39680 106148 39684
rect 106164 39740 106228 39744
rect 106164 39684 106168 39740
rect 106168 39684 106224 39740
rect 106224 39684 106228 39740
rect 106164 39680 106228 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 106660 39196 106724 39200
rect 106660 39140 106664 39196
rect 106664 39140 106720 39196
rect 106720 39140 106724 39196
rect 106660 39136 106724 39140
rect 106740 39196 106804 39200
rect 106740 39140 106744 39196
rect 106744 39140 106800 39196
rect 106800 39140 106804 39196
rect 106740 39136 106804 39140
rect 106820 39196 106884 39200
rect 106820 39140 106824 39196
rect 106824 39140 106880 39196
rect 106880 39140 106884 39196
rect 106820 39136 106884 39140
rect 106900 39196 106964 39200
rect 106900 39140 106904 39196
rect 106904 39140 106960 39196
rect 106960 39140 106964 39196
rect 106900 39136 106964 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 105924 38652 105988 38656
rect 105924 38596 105928 38652
rect 105928 38596 105984 38652
rect 105984 38596 105988 38652
rect 105924 38592 105988 38596
rect 106004 38652 106068 38656
rect 106004 38596 106008 38652
rect 106008 38596 106064 38652
rect 106064 38596 106068 38652
rect 106004 38592 106068 38596
rect 106084 38652 106148 38656
rect 106084 38596 106088 38652
rect 106088 38596 106144 38652
rect 106144 38596 106148 38652
rect 106084 38592 106148 38596
rect 106164 38652 106228 38656
rect 106164 38596 106168 38652
rect 106168 38596 106224 38652
rect 106224 38596 106228 38652
rect 106164 38592 106228 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 106660 38108 106724 38112
rect 106660 38052 106664 38108
rect 106664 38052 106720 38108
rect 106720 38052 106724 38108
rect 106660 38048 106724 38052
rect 106740 38108 106804 38112
rect 106740 38052 106744 38108
rect 106744 38052 106800 38108
rect 106800 38052 106804 38108
rect 106740 38048 106804 38052
rect 106820 38108 106884 38112
rect 106820 38052 106824 38108
rect 106824 38052 106880 38108
rect 106880 38052 106884 38108
rect 106820 38048 106884 38052
rect 106900 38108 106964 38112
rect 106900 38052 106904 38108
rect 106904 38052 106960 38108
rect 106960 38052 106964 38108
rect 106900 38048 106964 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 105924 37564 105988 37568
rect 105924 37508 105928 37564
rect 105928 37508 105984 37564
rect 105984 37508 105988 37564
rect 105924 37504 105988 37508
rect 106004 37564 106068 37568
rect 106004 37508 106008 37564
rect 106008 37508 106064 37564
rect 106064 37508 106068 37564
rect 106004 37504 106068 37508
rect 106084 37564 106148 37568
rect 106084 37508 106088 37564
rect 106088 37508 106144 37564
rect 106144 37508 106148 37564
rect 106084 37504 106148 37508
rect 106164 37564 106228 37568
rect 106164 37508 106168 37564
rect 106168 37508 106224 37564
rect 106224 37508 106228 37564
rect 106164 37504 106228 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 106660 37020 106724 37024
rect 106660 36964 106664 37020
rect 106664 36964 106720 37020
rect 106720 36964 106724 37020
rect 106660 36960 106724 36964
rect 106740 37020 106804 37024
rect 106740 36964 106744 37020
rect 106744 36964 106800 37020
rect 106800 36964 106804 37020
rect 106740 36960 106804 36964
rect 106820 37020 106884 37024
rect 106820 36964 106824 37020
rect 106824 36964 106880 37020
rect 106880 36964 106884 37020
rect 106820 36960 106884 36964
rect 106900 37020 106964 37024
rect 106900 36964 106904 37020
rect 106904 36964 106960 37020
rect 106960 36964 106964 37020
rect 106900 36960 106964 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 105924 36476 105988 36480
rect 105924 36420 105928 36476
rect 105928 36420 105984 36476
rect 105984 36420 105988 36476
rect 105924 36416 105988 36420
rect 106004 36476 106068 36480
rect 106004 36420 106008 36476
rect 106008 36420 106064 36476
rect 106064 36420 106068 36476
rect 106004 36416 106068 36420
rect 106084 36476 106148 36480
rect 106084 36420 106088 36476
rect 106088 36420 106144 36476
rect 106144 36420 106148 36476
rect 106084 36416 106148 36420
rect 106164 36476 106228 36480
rect 106164 36420 106168 36476
rect 106168 36420 106224 36476
rect 106224 36420 106228 36476
rect 106164 36416 106228 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 106660 35932 106724 35936
rect 106660 35876 106664 35932
rect 106664 35876 106720 35932
rect 106720 35876 106724 35932
rect 106660 35872 106724 35876
rect 106740 35932 106804 35936
rect 106740 35876 106744 35932
rect 106744 35876 106800 35932
rect 106800 35876 106804 35932
rect 106740 35872 106804 35876
rect 106820 35932 106884 35936
rect 106820 35876 106824 35932
rect 106824 35876 106880 35932
rect 106880 35876 106884 35932
rect 106820 35872 106884 35876
rect 106900 35932 106964 35936
rect 106900 35876 106904 35932
rect 106904 35876 106960 35932
rect 106960 35876 106964 35932
rect 106900 35872 106964 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 105924 35388 105988 35392
rect 105924 35332 105928 35388
rect 105928 35332 105984 35388
rect 105984 35332 105988 35388
rect 105924 35328 105988 35332
rect 106004 35388 106068 35392
rect 106004 35332 106008 35388
rect 106008 35332 106064 35388
rect 106064 35332 106068 35388
rect 106004 35328 106068 35332
rect 106084 35388 106148 35392
rect 106084 35332 106088 35388
rect 106088 35332 106144 35388
rect 106144 35332 106148 35388
rect 106084 35328 106148 35332
rect 106164 35388 106228 35392
rect 106164 35332 106168 35388
rect 106168 35332 106224 35388
rect 106224 35332 106228 35388
rect 106164 35328 106228 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 106660 34844 106724 34848
rect 106660 34788 106664 34844
rect 106664 34788 106720 34844
rect 106720 34788 106724 34844
rect 106660 34784 106724 34788
rect 106740 34844 106804 34848
rect 106740 34788 106744 34844
rect 106744 34788 106800 34844
rect 106800 34788 106804 34844
rect 106740 34784 106804 34788
rect 106820 34844 106884 34848
rect 106820 34788 106824 34844
rect 106824 34788 106880 34844
rect 106880 34788 106884 34844
rect 106820 34784 106884 34788
rect 106900 34844 106964 34848
rect 106900 34788 106904 34844
rect 106904 34788 106960 34844
rect 106960 34788 106964 34844
rect 106900 34784 106964 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 105924 34300 105988 34304
rect 105924 34244 105928 34300
rect 105928 34244 105984 34300
rect 105984 34244 105988 34300
rect 105924 34240 105988 34244
rect 106004 34300 106068 34304
rect 106004 34244 106008 34300
rect 106008 34244 106064 34300
rect 106064 34244 106068 34300
rect 106004 34240 106068 34244
rect 106084 34300 106148 34304
rect 106084 34244 106088 34300
rect 106088 34244 106144 34300
rect 106144 34244 106148 34300
rect 106084 34240 106148 34244
rect 106164 34300 106228 34304
rect 106164 34244 106168 34300
rect 106168 34244 106224 34300
rect 106224 34244 106228 34300
rect 106164 34240 106228 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 106660 33756 106724 33760
rect 106660 33700 106664 33756
rect 106664 33700 106720 33756
rect 106720 33700 106724 33756
rect 106660 33696 106724 33700
rect 106740 33756 106804 33760
rect 106740 33700 106744 33756
rect 106744 33700 106800 33756
rect 106800 33700 106804 33756
rect 106740 33696 106804 33700
rect 106820 33756 106884 33760
rect 106820 33700 106824 33756
rect 106824 33700 106880 33756
rect 106880 33700 106884 33756
rect 106820 33696 106884 33700
rect 106900 33756 106964 33760
rect 106900 33700 106904 33756
rect 106904 33700 106960 33756
rect 106960 33700 106964 33756
rect 106900 33696 106964 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 105924 33212 105988 33216
rect 105924 33156 105928 33212
rect 105928 33156 105984 33212
rect 105984 33156 105988 33212
rect 105924 33152 105988 33156
rect 106004 33212 106068 33216
rect 106004 33156 106008 33212
rect 106008 33156 106064 33212
rect 106064 33156 106068 33212
rect 106004 33152 106068 33156
rect 106084 33212 106148 33216
rect 106084 33156 106088 33212
rect 106088 33156 106144 33212
rect 106144 33156 106148 33212
rect 106084 33152 106148 33156
rect 106164 33212 106228 33216
rect 106164 33156 106168 33212
rect 106168 33156 106224 33212
rect 106224 33156 106228 33212
rect 106164 33152 106228 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 106660 32668 106724 32672
rect 106660 32612 106664 32668
rect 106664 32612 106720 32668
rect 106720 32612 106724 32668
rect 106660 32608 106724 32612
rect 106740 32668 106804 32672
rect 106740 32612 106744 32668
rect 106744 32612 106800 32668
rect 106800 32612 106804 32668
rect 106740 32608 106804 32612
rect 106820 32668 106884 32672
rect 106820 32612 106824 32668
rect 106824 32612 106880 32668
rect 106880 32612 106884 32668
rect 106820 32608 106884 32612
rect 106900 32668 106964 32672
rect 106900 32612 106904 32668
rect 106904 32612 106960 32668
rect 106960 32612 106964 32668
rect 106900 32608 106964 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 105924 32124 105988 32128
rect 105924 32068 105928 32124
rect 105928 32068 105984 32124
rect 105984 32068 105988 32124
rect 105924 32064 105988 32068
rect 106004 32124 106068 32128
rect 106004 32068 106008 32124
rect 106008 32068 106064 32124
rect 106064 32068 106068 32124
rect 106004 32064 106068 32068
rect 106084 32124 106148 32128
rect 106084 32068 106088 32124
rect 106088 32068 106144 32124
rect 106144 32068 106148 32124
rect 106084 32064 106148 32068
rect 106164 32124 106228 32128
rect 106164 32068 106168 32124
rect 106168 32068 106224 32124
rect 106224 32068 106228 32124
rect 106164 32064 106228 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 106660 31580 106724 31584
rect 106660 31524 106664 31580
rect 106664 31524 106720 31580
rect 106720 31524 106724 31580
rect 106660 31520 106724 31524
rect 106740 31580 106804 31584
rect 106740 31524 106744 31580
rect 106744 31524 106800 31580
rect 106800 31524 106804 31580
rect 106740 31520 106804 31524
rect 106820 31580 106884 31584
rect 106820 31524 106824 31580
rect 106824 31524 106880 31580
rect 106880 31524 106884 31580
rect 106820 31520 106884 31524
rect 106900 31580 106964 31584
rect 106900 31524 106904 31580
rect 106904 31524 106960 31580
rect 106960 31524 106964 31580
rect 106900 31520 106964 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 105924 31036 105988 31040
rect 105924 30980 105928 31036
rect 105928 30980 105984 31036
rect 105984 30980 105988 31036
rect 105924 30976 105988 30980
rect 106004 31036 106068 31040
rect 106004 30980 106008 31036
rect 106008 30980 106064 31036
rect 106064 30980 106068 31036
rect 106004 30976 106068 30980
rect 106084 31036 106148 31040
rect 106084 30980 106088 31036
rect 106088 30980 106144 31036
rect 106144 30980 106148 31036
rect 106084 30976 106148 30980
rect 106164 31036 106228 31040
rect 106164 30980 106168 31036
rect 106168 30980 106224 31036
rect 106224 30980 106228 31036
rect 106164 30976 106228 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 106660 30492 106724 30496
rect 106660 30436 106664 30492
rect 106664 30436 106720 30492
rect 106720 30436 106724 30492
rect 106660 30432 106724 30436
rect 106740 30492 106804 30496
rect 106740 30436 106744 30492
rect 106744 30436 106800 30492
rect 106800 30436 106804 30492
rect 106740 30432 106804 30436
rect 106820 30492 106884 30496
rect 106820 30436 106824 30492
rect 106824 30436 106880 30492
rect 106880 30436 106884 30492
rect 106820 30432 106884 30436
rect 106900 30492 106964 30496
rect 106900 30436 106904 30492
rect 106904 30436 106960 30492
rect 106960 30436 106964 30492
rect 106900 30432 106964 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 105924 29948 105988 29952
rect 105924 29892 105928 29948
rect 105928 29892 105984 29948
rect 105984 29892 105988 29948
rect 105924 29888 105988 29892
rect 106004 29948 106068 29952
rect 106004 29892 106008 29948
rect 106008 29892 106064 29948
rect 106064 29892 106068 29948
rect 106004 29888 106068 29892
rect 106084 29948 106148 29952
rect 106084 29892 106088 29948
rect 106088 29892 106144 29948
rect 106144 29892 106148 29948
rect 106084 29888 106148 29892
rect 106164 29948 106228 29952
rect 106164 29892 106168 29948
rect 106168 29892 106224 29948
rect 106224 29892 106228 29948
rect 106164 29888 106228 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 106660 29404 106724 29408
rect 106660 29348 106664 29404
rect 106664 29348 106720 29404
rect 106720 29348 106724 29404
rect 106660 29344 106724 29348
rect 106740 29404 106804 29408
rect 106740 29348 106744 29404
rect 106744 29348 106800 29404
rect 106800 29348 106804 29404
rect 106740 29344 106804 29348
rect 106820 29404 106884 29408
rect 106820 29348 106824 29404
rect 106824 29348 106880 29404
rect 106880 29348 106884 29404
rect 106820 29344 106884 29348
rect 106900 29404 106964 29408
rect 106900 29348 106904 29404
rect 106904 29348 106960 29404
rect 106960 29348 106964 29404
rect 106900 29344 106964 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 105924 28860 105988 28864
rect 105924 28804 105928 28860
rect 105928 28804 105984 28860
rect 105984 28804 105988 28860
rect 105924 28800 105988 28804
rect 106004 28860 106068 28864
rect 106004 28804 106008 28860
rect 106008 28804 106064 28860
rect 106064 28804 106068 28860
rect 106004 28800 106068 28804
rect 106084 28860 106148 28864
rect 106084 28804 106088 28860
rect 106088 28804 106144 28860
rect 106144 28804 106148 28860
rect 106084 28800 106148 28804
rect 106164 28860 106228 28864
rect 106164 28804 106168 28860
rect 106168 28804 106224 28860
rect 106224 28804 106228 28860
rect 106164 28800 106228 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 106660 28316 106724 28320
rect 106660 28260 106664 28316
rect 106664 28260 106720 28316
rect 106720 28260 106724 28316
rect 106660 28256 106724 28260
rect 106740 28316 106804 28320
rect 106740 28260 106744 28316
rect 106744 28260 106800 28316
rect 106800 28260 106804 28316
rect 106740 28256 106804 28260
rect 106820 28316 106884 28320
rect 106820 28260 106824 28316
rect 106824 28260 106880 28316
rect 106880 28260 106884 28316
rect 106820 28256 106884 28260
rect 106900 28316 106964 28320
rect 106900 28260 106904 28316
rect 106904 28260 106960 28316
rect 106960 28260 106964 28316
rect 106900 28256 106964 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 105924 27772 105988 27776
rect 105924 27716 105928 27772
rect 105928 27716 105984 27772
rect 105984 27716 105988 27772
rect 105924 27712 105988 27716
rect 106004 27772 106068 27776
rect 106004 27716 106008 27772
rect 106008 27716 106064 27772
rect 106064 27716 106068 27772
rect 106004 27712 106068 27716
rect 106084 27772 106148 27776
rect 106084 27716 106088 27772
rect 106088 27716 106144 27772
rect 106144 27716 106148 27772
rect 106084 27712 106148 27716
rect 106164 27772 106228 27776
rect 106164 27716 106168 27772
rect 106168 27716 106224 27772
rect 106224 27716 106228 27772
rect 106164 27712 106228 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 106660 27228 106724 27232
rect 106660 27172 106664 27228
rect 106664 27172 106720 27228
rect 106720 27172 106724 27228
rect 106660 27168 106724 27172
rect 106740 27228 106804 27232
rect 106740 27172 106744 27228
rect 106744 27172 106800 27228
rect 106800 27172 106804 27228
rect 106740 27168 106804 27172
rect 106820 27228 106884 27232
rect 106820 27172 106824 27228
rect 106824 27172 106880 27228
rect 106880 27172 106884 27228
rect 106820 27168 106884 27172
rect 106900 27228 106964 27232
rect 106900 27172 106904 27228
rect 106904 27172 106960 27228
rect 106960 27172 106964 27228
rect 106900 27168 106964 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 105924 26684 105988 26688
rect 105924 26628 105928 26684
rect 105928 26628 105984 26684
rect 105984 26628 105988 26684
rect 105924 26624 105988 26628
rect 106004 26684 106068 26688
rect 106004 26628 106008 26684
rect 106008 26628 106064 26684
rect 106064 26628 106068 26684
rect 106004 26624 106068 26628
rect 106084 26684 106148 26688
rect 106084 26628 106088 26684
rect 106088 26628 106144 26684
rect 106144 26628 106148 26684
rect 106084 26624 106148 26628
rect 106164 26684 106228 26688
rect 106164 26628 106168 26684
rect 106168 26628 106224 26684
rect 106224 26628 106228 26684
rect 106164 26624 106228 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 106660 26140 106724 26144
rect 106660 26084 106664 26140
rect 106664 26084 106720 26140
rect 106720 26084 106724 26140
rect 106660 26080 106724 26084
rect 106740 26140 106804 26144
rect 106740 26084 106744 26140
rect 106744 26084 106800 26140
rect 106800 26084 106804 26140
rect 106740 26080 106804 26084
rect 106820 26140 106884 26144
rect 106820 26084 106824 26140
rect 106824 26084 106880 26140
rect 106880 26084 106884 26140
rect 106820 26080 106884 26084
rect 106900 26140 106964 26144
rect 106900 26084 106904 26140
rect 106904 26084 106960 26140
rect 106960 26084 106964 26140
rect 106900 26080 106964 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 105924 25596 105988 25600
rect 105924 25540 105928 25596
rect 105928 25540 105984 25596
rect 105984 25540 105988 25596
rect 105924 25536 105988 25540
rect 106004 25596 106068 25600
rect 106004 25540 106008 25596
rect 106008 25540 106064 25596
rect 106064 25540 106068 25596
rect 106004 25536 106068 25540
rect 106084 25596 106148 25600
rect 106084 25540 106088 25596
rect 106088 25540 106144 25596
rect 106144 25540 106148 25596
rect 106084 25536 106148 25540
rect 106164 25596 106228 25600
rect 106164 25540 106168 25596
rect 106168 25540 106224 25596
rect 106224 25540 106228 25596
rect 106164 25536 106228 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 106660 25052 106724 25056
rect 106660 24996 106664 25052
rect 106664 24996 106720 25052
rect 106720 24996 106724 25052
rect 106660 24992 106724 24996
rect 106740 25052 106804 25056
rect 106740 24996 106744 25052
rect 106744 24996 106800 25052
rect 106800 24996 106804 25052
rect 106740 24992 106804 24996
rect 106820 25052 106884 25056
rect 106820 24996 106824 25052
rect 106824 24996 106880 25052
rect 106880 24996 106884 25052
rect 106820 24992 106884 24996
rect 106900 25052 106964 25056
rect 106900 24996 106904 25052
rect 106904 24996 106960 25052
rect 106960 24996 106964 25052
rect 106900 24992 106964 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 105924 24508 105988 24512
rect 105924 24452 105928 24508
rect 105928 24452 105984 24508
rect 105984 24452 105988 24508
rect 105924 24448 105988 24452
rect 106004 24508 106068 24512
rect 106004 24452 106008 24508
rect 106008 24452 106064 24508
rect 106064 24452 106068 24508
rect 106004 24448 106068 24452
rect 106084 24508 106148 24512
rect 106084 24452 106088 24508
rect 106088 24452 106144 24508
rect 106144 24452 106148 24508
rect 106084 24448 106148 24452
rect 106164 24508 106228 24512
rect 106164 24452 106168 24508
rect 106168 24452 106224 24508
rect 106224 24452 106228 24508
rect 106164 24448 106228 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 106660 23964 106724 23968
rect 106660 23908 106664 23964
rect 106664 23908 106720 23964
rect 106720 23908 106724 23964
rect 106660 23904 106724 23908
rect 106740 23964 106804 23968
rect 106740 23908 106744 23964
rect 106744 23908 106800 23964
rect 106800 23908 106804 23964
rect 106740 23904 106804 23908
rect 106820 23964 106884 23968
rect 106820 23908 106824 23964
rect 106824 23908 106880 23964
rect 106880 23908 106884 23964
rect 106820 23904 106884 23908
rect 106900 23964 106964 23968
rect 106900 23908 106904 23964
rect 106904 23908 106960 23964
rect 106960 23908 106964 23964
rect 106900 23904 106964 23908
rect 102732 23488 102796 23492
rect 102732 23432 102782 23488
rect 102782 23432 102796 23488
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 102732 23428 102796 23432
rect 105924 23420 105988 23424
rect 105924 23364 105928 23420
rect 105928 23364 105984 23420
rect 105984 23364 105988 23420
rect 105924 23360 105988 23364
rect 106004 23420 106068 23424
rect 106004 23364 106008 23420
rect 106008 23364 106064 23420
rect 106064 23364 106068 23420
rect 106004 23360 106068 23364
rect 106084 23420 106148 23424
rect 106084 23364 106088 23420
rect 106088 23364 106144 23420
rect 106144 23364 106148 23420
rect 106084 23360 106148 23364
rect 106164 23420 106228 23424
rect 106164 23364 106168 23420
rect 106168 23364 106224 23420
rect 106224 23364 106228 23420
rect 106164 23360 106228 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 106660 22876 106724 22880
rect 106660 22820 106664 22876
rect 106664 22820 106720 22876
rect 106720 22820 106724 22876
rect 106660 22816 106724 22820
rect 106740 22876 106804 22880
rect 106740 22820 106744 22876
rect 106744 22820 106800 22876
rect 106800 22820 106804 22876
rect 106740 22816 106804 22820
rect 106820 22876 106884 22880
rect 106820 22820 106824 22876
rect 106824 22820 106880 22876
rect 106880 22820 106884 22876
rect 106820 22816 106884 22820
rect 106900 22876 106964 22880
rect 106900 22820 106904 22876
rect 106904 22820 106960 22876
rect 106960 22820 106964 22876
rect 106900 22816 106964 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 105924 22332 105988 22336
rect 105924 22276 105928 22332
rect 105928 22276 105984 22332
rect 105984 22276 105988 22332
rect 105924 22272 105988 22276
rect 106004 22332 106068 22336
rect 106004 22276 106008 22332
rect 106008 22276 106064 22332
rect 106064 22276 106068 22332
rect 106004 22272 106068 22276
rect 106084 22332 106148 22336
rect 106084 22276 106088 22332
rect 106088 22276 106144 22332
rect 106144 22276 106148 22332
rect 106084 22272 106148 22276
rect 106164 22332 106228 22336
rect 106164 22276 106168 22332
rect 106168 22276 106224 22332
rect 106224 22276 106228 22332
rect 106164 22272 106228 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 106660 21788 106724 21792
rect 106660 21732 106664 21788
rect 106664 21732 106720 21788
rect 106720 21732 106724 21788
rect 106660 21728 106724 21732
rect 106740 21788 106804 21792
rect 106740 21732 106744 21788
rect 106744 21732 106800 21788
rect 106800 21732 106804 21788
rect 106740 21728 106804 21732
rect 106820 21788 106884 21792
rect 106820 21732 106824 21788
rect 106824 21732 106880 21788
rect 106880 21732 106884 21788
rect 106820 21728 106884 21732
rect 106900 21788 106964 21792
rect 106900 21732 106904 21788
rect 106904 21732 106960 21788
rect 106960 21732 106964 21788
rect 106900 21728 106964 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 105924 21244 105988 21248
rect 105924 21188 105928 21244
rect 105928 21188 105984 21244
rect 105984 21188 105988 21244
rect 105924 21184 105988 21188
rect 106004 21244 106068 21248
rect 106004 21188 106008 21244
rect 106008 21188 106064 21244
rect 106064 21188 106068 21244
rect 106004 21184 106068 21188
rect 106084 21244 106148 21248
rect 106084 21188 106088 21244
rect 106088 21188 106144 21244
rect 106144 21188 106148 21244
rect 106084 21184 106148 21188
rect 106164 21244 106228 21248
rect 106164 21188 106168 21244
rect 106168 21188 106224 21244
rect 106224 21188 106228 21244
rect 106164 21184 106228 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 106660 20700 106724 20704
rect 106660 20644 106664 20700
rect 106664 20644 106720 20700
rect 106720 20644 106724 20700
rect 106660 20640 106724 20644
rect 106740 20700 106804 20704
rect 106740 20644 106744 20700
rect 106744 20644 106800 20700
rect 106800 20644 106804 20700
rect 106740 20640 106804 20644
rect 106820 20700 106884 20704
rect 106820 20644 106824 20700
rect 106824 20644 106880 20700
rect 106880 20644 106884 20700
rect 106820 20640 106884 20644
rect 106900 20700 106964 20704
rect 106900 20644 106904 20700
rect 106904 20644 106960 20700
rect 106960 20644 106964 20700
rect 106900 20640 106964 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 105924 20156 105988 20160
rect 105924 20100 105928 20156
rect 105928 20100 105984 20156
rect 105984 20100 105988 20156
rect 105924 20096 105988 20100
rect 106004 20156 106068 20160
rect 106004 20100 106008 20156
rect 106008 20100 106064 20156
rect 106064 20100 106068 20156
rect 106004 20096 106068 20100
rect 106084 20156 106148 20160
rect 106084 20100 106088 20156
rect 106088 20100 106144 20156
rect 106144 20100 106148 20156
rect 106084 20096 106148 20100
rect 106164 20156 106228 20160
rect 106164 20100 106168 20156
rect 106168 20100 106224 20156
rect 106224 20100 106228 20156
rect 106164 20096 106228 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 106660 19612 106724 19616
rect 106660 19556 106664 19612
rect 106664 19556 106720 19612
rect 106720 19556 106724 19612
rect 106660 19552 106724 19556
rect 106740 19612 106804 19616
rect 106740 19556 106744 19612
rect 106744 19556 106800 19612
rect 106800 19556 106804 19612
rect 106740 19552 106804 19556
rect 106820 19612 106884 19616
rect 106820 19556 106824 19612
rect 106824 19556 106880 19612
rect 106880 19556 106884 19612
rect 106820 19552 106884 19556
rect 106900 19612 106964 19616
rect 106900 19556 106904 19612
rect 106904 19556 106960 19612
rect 106960 19556 106964 19612
rect 106900 19552 106964 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 105924 19068 105988 19072
rect 105924 19012 105928 19068
rect 105928 19012 105984 19068
rect 105984 19012 105988 19068
rect 105924 19008 105988 19012
rect 106004 19068 106068 19072
rect 106004 19012 106008 19068
rect 106008 19012 106064 19068
rect 106064 19012 106068 19068
rect 106004 19008 106068 19012
rect 106084 19068 106148 19072
rect 106084 19012 106088 19068
rect 106088 19012 106144 19068
rect 106144 19012 106148 19068
rect 106084 19008 106148 19012
rect 106164 19068 106228 19072
rect 106164 19012 106168 19068
rect 106168 19012 106224 19068
rect 106224 19012 106228 19068
rect 106164 19008 106228 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 106660 18524 106724 18528
rect 106660 18468 106664 18524
rect 106664 18468 106720 18524
rect 106720 18468 106724 18524
rect 106660 18464 106724 18468
rect 106740 18524 106804 18528
rect 106740 18468 106744 18524
rect 106744 18468 106800 18524
rect 106800 18468 106804 18524
rect 106740 18464 106804 18468
rect 106820 18524 106884 18528
rect 106820 18468 106824 18524
rect 106824 18468 106880 18524
rect 106880 18468 106884 18524
rect 106820 18464 106884 18468
rect 106900 18524 106964 18528
rect 106900 18468 106904 18524
rect 106904 18468 106960 18524
rect 106960 18468 106964 18524
rect 106900 18464 106964 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 105924 17980 105988 17984
rect 105924 17924 105928 17980
rect 105928 17924 105984 17980
rect 105984 17924 105988 17980
rect 105924 17920 105988 17924
rect 106004 17980 106068 17984
rect 106004 17924 106008 17980
rect 106008 17924 106064 17980
rect 106064 17924 106068 17980
rect 106004 17920 106068 17924
rect 106084 17980 106148 17984
rect 106084 17924 106088 17980
rect 106088 17924 106144 17980
rect 106144 17924 106148 17980
rect 106084 17920 106148 17924
rect 106164 17980 106228 17984
rect 106164 17924 106168 17980
rect 106168 17924 106224 17980
rect 106224 17924 106228 17980
rect 106164 17920 106228 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 106660 17436 106724 17440
rect 106660 17380 106664 17436
rect 106664 17380 106720 17436
rect 106720 17380 106724 17436
rect 106660 17376 106724 17380
rect 106740 17436 106804 17440
rect 106740 17380 106744 17436
rect 106744 17380 106800 17436
rect 106800 17380 106804 17436
rect 106740 17376 106804 17380
rect 106820 17436 106884 17440
rect 106820 17380 106824 17436
rect 106824 17380 106880 17436
rect 106880 17380 106884 17436
rect 106820 17376 106884 17380
rect 106900 17436 106964 17440
rect 106900 17380 106904 17436
rect 106904 17380 106960 17436
rect 106960 17380 106964 17436
rect 106900 17376 106964 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 105924 16892 105988 16896
rect 105924 16836 105928 16892
rect 105928 16836 105984 16892
rect 105984 16836 105988 16892
rect 105924 16832 105988 16836
rect 106004 16892 106068 16896
rect 106004 16836 106008 16892
rect 106008 16836 106064 16892
rect 106064 16836 106068 16892
rect 106004 16832 106068 16836
rect 106084 16892 106148 16896
rect 106084 16836 106088 16892
rect 106088 16836 106144 16892
rect 106144 16836 106148 16892
rect 106084 16832 106148 16836
rect 106164 16892 106228 16896
rect 106164 16836 106168 16892
rect 106168 16836 106224 16892
rect 106224 16836 106228 16892
rect 106164 16832 106228 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 106660 16348 106724 16352
rect 106660 16292 106664 16348
rect 106664 16292 106720 16348
rect 106720 16292 106724 16348
rect 106660 16288 106724 16292
rect 106740 16348 106804 16352
rect 106740 16292 106744 16348
rect 106744 16292 106800 16348
rect 106800 16292 106804 16348
rect 106740 16288 106804 16292
rect 106820 16348 106884 16352
rect 106820 16292 106824 16348
rect 106824 16292 106880 16348
rect 106880 16292 106884 16348
rect 106820 16288 106884 16292
rect 106900 16348 106964 16352
rect 106900 16292 106904 16348
rect 106904 16292 106960 16348
rect 106960 16292 106964 16348
rect 106900 16288 106964 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 105924 15804 105988 15808
rect 105924 15748 105928 15804
rect 105928 15748 105984 15804
rect 105984 15748 105988 15804
rect 105924 15744 105988 15748
rect 106004 15804 106068 15808
rect 106004 15748 106008 15804
rect 106008 15748 106064 15804
rect 106064 15748 106068 15804
rect 106004 15744 106068 15748
rect 106084 15804 106148 15808
rect 106084 15748 106088 15804
rect 106088 15748 106144 15804
rect 106144 15748 106148 15804
rect 106084 15744 106148 15748
rect 106164 15804 106228 15808
rect 106164 15748 106168 15804
rect 106168 15748 106224 15804
rect 106224 15748 106228 15804
rect 106164 15744 106228 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 106660 15260 106724 15264
rect 106660 15204 106664 15260
rect 106664 15204 106720 15260
rect 106720 15204 106724 15260
rect 106660 15200 106724 15204
rect 106740 15260 106804 15264
rect 106740 15204 106744 15260
rect 106744 15204 106800 15260
rect 106800 15204 106804 15260
rect 106740 15200 106804 15204
rect 106820 15260 106884 15264
rect 106820 15204 106824 15260
rect 106824 15204 106880 15260
rect 106880 15204 106884 15260
rect 106820 15200 106884 15204
rect 106900 15260 106964 15264
rect 106900 15204 106904 15260
rect 106904 15204 106960 15260
rect 106960 15204 106964 15260
rect 106900 15200 106964 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 105924 14716 105988 14720
rect 105924 14660 105928 14716
rect 105928 14660 105984 14716
rect 105984 14660 105988 14716
rect 105924 14656 105988 14660
rect 106004 14716 106068 14720
rect 106004 14660 106008 14716
rect 106008 14660 106064 14716
rect 106064 14660 106068 14716
rect 106004 14656 106068 14660
rect 106084 14716 106148 14720
rect 106084 14660 106088 14716
rect 106088 14660 106144 14716
rect 106144 14660 106148 14716
rect 106084 14656 106148 14660
rect 106164 14716 106228 14720
rect 106164 14660 106168 14716
rect 106168 14660 106224 14716
rect 106224 14660 106228 14716
rect 106164 14656 106228 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 106660 14172 106724 14176
rect 106660 14116 106664 14172
rect 106664 14116 106720 14172
rect 106720 14116 106724 14172
rect 106660 14112 106724 14116
rect 106740 14172 106804 14176
rect 106740 14116 106744 14172
rect 106744 14116 106800 14172
rect 106800 14116 106804 14172
rect 106740 14112 106804 14116
rect 106820 14172 106884 14176
rect 106820 14116 106824 14172
rect 106824 14116 106880 14172
rect 106880 14116 106884 14172
rect 106820 14112 106884 14116
rect 106900 14172 106964 14176
rect 106900 14116 106904 14172
rect 106904 14116 106960 14172
rect 106960 14116 106964 14172
rect 106900 14112 106964 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 105924 13628 105988 13632
rect 105924 13572 105928 13628
rect 105928 13572 105984 13628
rect 105984 13572 105988 13628
rect 105924 13568 105988 13572
rect 106004 13628 106068 13632
rect 106004 13572 106008 13628
rect 106008 13572 106064 13628
rect 106064 13572 106068 13628
rect 106004 13568 106068 13572
rect 106084 13628 106148 13632
rect 106084 13572 106088 13628
rect 106088 13572 106144 13628
rect 106144 13572 106148 13628
rect 106084 13568 106148 13572
rect 106164 13628 106228 13632
rect 106164 13572 106168 13628
rect 106168 13572 106224 13628
rect 106224 13572 106228 13628
rect 106164 13568 106228 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 106660 13084 106724 13088
rect 106660 13028 106664 13084
rect 106664 13028 106720 13084
rect 106720 13028 106724 13084
rect 106660 13024 106724 13028
rect 106740 13084 106804 13088
rect 106740 13028 106744 13084
rect 106744 13028 106800 13084
rect 106800 13028 106804 13084
rect 106740 13024 106804 13028
rect 106820 13084 106884 13088
rect 106820 13028 106824 13084
rect 106824 13028 106880 13084
rect 106880 13028 106884 13084
rect 106820 13024 106884 13028
rect 106900 13084 106964 13088
rect 106900 13028 106904 13084
rect 106904 13028 106960 13084
rect 106960 13028 106964 13084
rect 106900 13024 106964 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 105924 12540 105988 12544
rect 105924 12484 105928 12540
rect 105928 12484 105984 12540
rect 105984 12484 105988 12540
rect 105924 12480 105988 12484
rect 106004 12540 106068 12544
rect 106004 12484 106008 12540
rect 106008 12484 106064 12540
rect 106064 12484 106068 12540
rect 106004 12480 106068 12484
rect 106084 12540 106148 12544
rect 106084 12484 106088 12540
rect 106088 12484 106144 12540
rect 106144 12484 106148 12540
rect 106084 12480 106148 12484
rect 106164 12540 106228 12544
rect 106164 12484 106168 12540
rect 106168 12484 106224 12540
rect 106224 12484 106228 12540
rect 106164 12480 106228 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 106660 11996 106724 12000
rect 106660 11940 106664 11996
rect 106664 11940 106720 11996
rect 106720 11940 106724 11996
rect 106660 11936 106724 11940
rect 106740 11996 106804 12000
rect 106740 11940 106744 11996
rect 106744 11940 106800 11996
rect 106800 11940 106804 11996
rect 106740 11936 106804 11940
rect 106820 11996 106884 12000
rect 106820 11940 106824 11996
rect 106824 11940 106880 11996
rect 106880 11940 106884 11996
rect 106820 11936 106884 11940
rect 106900 11996 106964 12000
rect 106900 11940 106904 11996
rect 106904 11940 106960 11996
rect 106960 11940 106964 11996
rect 106900 11936 106964 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 105924 11452 105988 11456
rect 105924 11396 105928 11452
rect 105928 11396 105984 11452
rect 105984 11396 105988 11452
rect 105924 11392 105988 11396
rect 106004 11452 106068 11456
rect 106004 11396 106008 11452
rect 106008 11396 106064 11452
rect 106064 11396 106068 11452
rect 106004 11392 106068 11396
rect 106084 11452 106148 11456
rect 106084 11396 106088 11452
rect 106088 11396 106144 11452
rect 106144 11396 106148 11452
rect 106084 11392 106148 11396
rect 106164 11452 106228 11456
rect 106164 11396 106168 11452
rect 106168 11396 106224 11452
rect 106224 11396 106228 11452
rect 106164 11392 106228 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 106660 10908 106724 10912
rect 106660 10852 106664 10908
rect 106664 10852 106720 10908
rect 106720 10852 106724 10908
rect 106660 10848 106724 10852
rect 106740 10908 106804 10912
rect 106740 10852 106744 10908
rect 106744 10852 106800 10908
rect 106800 10852 106804 10908
rect 106740 10848 106804 10852
rect 106820 10908 106884 10912
rect 106820 10852 106824 10908
rect 106824 10852 106880 10908
rect 106880 10852 106884 10908
rect 106820 10848 106884 10852
rect 106900 10908 106964 10912
rect 106900 10852 106904 10908
rect 106904 10852 106960 10908
rect 106960 10852 106964 10908
rect 106900 10848 106964 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 105924 10364 105988 10368
rect 105924 10308 105928 10364
rect 105928 10308 105984 10364
rect 105984 10308 105988 10364
rect 105924 10304 105988 10308
rect 106004 10364 106068 10368
rect 106004 10308 106008 10364
rect 106008 10308 106064 10364
rect 106064 10308 106068 10364
rect 106004 10304 106068 10308
rect 106084 10364 106148 10368
rect 106084 10308 106088 10364
rect 106088 10308 106144 10364
rect 106144 10308 106148 10364
rect 106084 10304 106148 10308
rect 106164 10364 106228 10368
rect 106164 10308 106168 10364
rect 106168 10308 106224 10364
rect 106224 10308 106228 10364
rect 106164 10304 106228 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 106660 9820 106724 9824
rect 106660 9764 106664 9820
rect 106664 9764 106720 9820
rect 106720 9764 106724 9820
rect 106660 9760 106724 9764
rect 106740 9820 106804 9824
rect 106740 9764 106744 9820
rect 106744 9764 106800 9820
rect 106800 9764 106804 9820
rect 106740 9760 106804 9764
rect 106820 9820 106884 9824
rect 106820 9764 106824 9820
rect 106824 9764 106880 9820
rect 106880 9764 106884 9820
rect 106820 9760 106884 9764
rect 106900 9820 106964 9824
rect 106900 9764 106904 9820
rect 106904 9764 106960 9820
rect 106960 9764 106964 9820
rect 106900 9760 106964 9764
rect 23438 9752 23502 9756
rect 23438 9696 23478 9752
rect 23478 9696 23502 9752
rect 23438 9692 23502 9696
rect 25774 9752 25838 9756
rect 25774 9696 25778 9752
rect 25778 9696 25834 9752
rect 25834 9696 25838 9752
rect 25774 9692 25838 9696
rect 28120 9752 28184 9756
rect 28120 9696 28170 9752
rect 28170 9696 28184 9752
rect 28120 9692 28184 9696
rect 29278 9692 29342 9756
rect 30446 9752 30510 9756
rect 30446 9696 30470 9752
rect 30470 9696 30510 9752
rect 30446 9692 30510 9696
rect 16058 9616 16122 9620
rect 16058 9560 16082 9616
rect 16082 9560 16122 9616
rect 16058 9556 16122 9560
rect 24624 9616 24688 9620
rect 24624 9560 24674 9616
rect 24674 9560 24688 9616
rect 24624 9556 24688 9560
rect 90665 9616 90729 9620
rect 90665 9560 90694 9616
rect 90694 9560 90729 9616
rect 90665 9556 90729 9560
rect 90814 9616 90878 9620
rect 90814 9560 90822 9616
rect 90822 9560 90878 9616
rect 90814 9556 90878 9560
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 105924 9276 105988 9280
rect 105924 9220 105928 9276
rect 105928 9220 105984 9276
rect 105984 9220 105988 9276
rect 105924 9216 105988 9220
rect 106004 9276 106068 9280
rect 106004 9220 106008 9276
rect 106008 9220 106064 9276
rect 106064 9220 106068 9276
rect 106004 9216 106068 9220
rect 106084 9276 106148 9280
rect 106084 9220 106088 9276
rect 106088 9220 106144 9276
rect 106144 9220 106148 9276
rect 106084 9216 106148 9220
rect 106164 9276 106228 9280
rect 106164 9220 106168 9276
rect 106168 9220 106224 9276
rect 106224 9220 106228 9276
rect 106164 9216 106228 9220
rect 26924 8876 26988 8940
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 106660 8732 106724 8736
rect 106660 8676 106664 8732
rect 106664 8676 106720 8732
rect 106720 8676 106724 8732
rect 106660 8672 106724 8676
rect 106740 8732 106804 8736
rect 106740 8676 106744 8732
rect 106744 8676 106800 8732
rect 106800 8676 106804 8732
rect 106740 8672 106804 8676
rect 106820 8732 106884 8736
rect 106820 8676 106824 8732
rect 106824 8676 106880 8732
rect 106880 8676 106884 8732
rect 106820 8672 106884 8676
rect 106900 8732 106964 8736
rect 106900 8676 106904 8732
rect 106904 8676 106960 8732
rect 106960 8676 106964 8732
rect 106900 8672 106964 8676
rect 90404 8332 90468 8396
rect 31708 8256 31772 8260
rect 31708 8200 31722 8256
rect 31722 8200 31772 8256
rect 31708 8196 31772 8200
rect 32812 8196 32876 8260
rect 33916 8196 33980 8260
rect 35204 8196 35268 8260
rect 36308 8256 36372 8260
rect 36308 8200 36358 8256
rect 36358 8200 36372 8256
rect 36308 8196 36372 8200
rect 37412 8256 37476 8260
rect 37412 8200 37462 8256
rect 37462 8200 37476 8256
rect 37412 8196 37476 8200
rect 38700 8256 38764 8260
rect 38700 8200 38750 8256
rect 38750 8200 38764 8256
rect 38700 8196 38764 8200
rect 40908 8196 40972 8260
rect 42196 8256 42260 8260
rect 42196 8200 42210 8256
rect 42210 8200 42260 8256
rect 42196 8196 42260 8200
rect 43300 8196 43364 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 105924 8188 105988 8192
rect 105924 8132 105928 8188
rect 105928 8132 105984 8188
rect 105984 8132 105988 8188
rect 105924 8128 105988 8132
rect 106004 8188 106068 8192
rect 106004 8132 106008 8188
rect 106008 8132 106064 8188
rect 106064 8132 106068 8188
rect 106004 8128 106068 8132
rect 106084 8188 106148 8192
rect 106084 8132 106088 8188
rect 106088 8132 106144 8188
rect 106144 8132 106148 8188
rect 106084 8128 106148 8132
rect 106164 8188 106228 8192
rect 106164 8132 106168 8188
rect 106168 8132 106224 8188
rect 106224 8132 106228 8188
rect 106164 8128 106228 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 66316 7644 66380 7648
rect 66316 7588 66320 7644
rect 66320 7588 66376 7644
rect 66376 7588 66380 7644
rect 66316 7584 66380 7588
rect 66396 7644 66460 7648
rect 66396 7588 66400 7644
rect 66400 7588 66456 7644
rect 66456 7588 66460 7644
rect 66396 7584 66460 7588
rect 66476 7644 66540 7648
rect 66476 7588 66480 7644
rect 66480 7588 66536 7644
rect 66536 7588 66540 7644
rect 66476 7584 66540 7588
rect 66556 7644 66620 7648
rect 66556 7588 66560 7644
rect 66560 7588 66616 7644
rect 66616 7588 66620 7644
rect 66556 7584 66620 7588
rect 97036 7644 97100 7648
rect 97036 7588 97040 7644
rect 97040 7588 97096 7644
rect 97096 7588 97100 7644
rect 97036 7584 97100 7588
rect 97116 7644 97180 7648
rect 97116 7588 97120 7644
rect 97120 7588 97176 7644
rect 97176 7588 97180 7644
rect 97116 7584 97180 7588
rect 97196 7644 97260 7648
rect 97196 7588 97200 7644
rect 97200 7588 97256 7644
rect 97256 7588 97260 7644
rect 97196 7584 97260 7588
rect 97276 7644 97340 7648
rect 97276 7588 97280 7644
rect 97280 7588 97336 7644
rect 97336 7588 97340 7644
rect 97276 7584 97340 7588
rect 106660 7644 106724 7648
rect 106660 7588 106664 7644
rect 106664 7588 106720 7644
rect 106720 7588 106724 7644
rect 106660 7584 106724 7588
rect 106740 7644 106804 7648
rect 106740 7588 106744 7644
rect 106744 7588 106800 7644
rect 106800 7588 106804 7644
rect 106740 7584 106804 7588
rect 106820 7644 106884 7648
rect 106820 7588 106824 7644
rect 106824 7588 106880 7644
rect 106880 7588 106884 7644
rect 106820 7584 106884 7588
rect 106900 7644 106964 7648
rect 106900 7588 106904 7644
rect 106904 7588 106960 7644
rect 106960 7588 106964 7644
rect 106900 7584 106964 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 105924 7100 105988 7104
rect 105924 7044 105928 7100
rect 105928 7044 105984 7100
rect 105984 7044 105988 7100
rect 105924 7040 105988 7044
rect 106004 7100 106068 7104
rect 106004 7044 106008 7100
rect 106008 7044 106064 7100
rect 106064 7044 106068 7100
rect 106004 7040 106068 7044
rect 106084 7100 106148 7104
rect 106084 7044 106088 7100
rect 106088 7044 106144 7100
rect 106144 7044 106148 7100
rect 106084 7040 106148 7044
rect 106164 7100 106228 7104
rect 106164 7044 106168 7100
rect 106168 7044 106224 7100
rect 106224 7044 106228 7100
rect 106164 7040 106228 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 66316 6556 66380 6560
rect 66316 6500 66320 6556
rect 66320 6500 66376 6556
rect 66376 6500 66380 6556
rect 66316 6496 66380 6500
rect 66396 6556 66460 6560
rect 66396 6500 66400 6556
rect 66400 6500 66456 6556
rect 66456 6500 66460 6556
rect 66396 6496 66460 6500
rect 66476 6556 66540 6560
rect 66476 6500 66480 6556
rect 66480 6500 66536 6556
rect 66536 6500 66540 6556
rect 66476 6496 66540 6500
rect 66556 6556 66620 6560
rect 66556 6500 66560 6556
rect 66560 6500 66616 6556
rect 66616 6500 66620 6556
rect 66556 6496 66620 6500
rect 97036 6556 97100 6560
rect 97036 6500 97040 6556
rect 97040 6500 97096 6556
rect 97096 6500 97100 6556
rect 97036 6496 97100 6500
rect 97116 6556 97180 6560
rect 97116 6500 97120 6556
rect 97120 6500 97176 6556
rect 97176 6500 97180 6556
rect 97116 6496 97180 6500
rect 97196 6556 97260 6560
rect 97196 6500 97200 6556
rect 97200 6500 97256 6556
rect 97256 6500 97260 6556
rect 97196 6496 97260 6500
rect 97276 6556 97340 6560
rect 97276 6500 97280 6556
rect 97280 6500 97336 6556
rect 97336 6500 97340 6556
rect 97276 6496 97340 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 66316 5468 66380 5472
rect 66316 5412 66320 5468
rect 66320 5412 66376 5468
rect 66376 5412 66380 5468
rect 66316 5408 66380 5412
rect 66396 5468 66460 5472
rect 66396 5412 66400 5468
rect 66400 5412 66456 5468
rect 66456 5412 66460 5468
rect 66396 5408 66460 5412
rect 66476 5468 66540 5472
rect 66476 5412 66480 5468
rect 66480 5412 66536 5468
rect 66536 5412 66540 5468
rect 66476 5408 66540 5412
rect 66556 5468 66620 5472
rect 66556 5412 66560 5468
rect 66560 5412 66616 5468
rect 66616 5412 66620 5468
rect 66556 5408 66620 5412
rect 97036 5468 97100 5472
rect 97036 5412 97040 5468
rect 97040 5412 97096 5468
rect 97096 5412 97100 5468
rect 97036 5408 97100 5412
rect 97116 5468 97180 5472
rect 97116 5412 97120 5468
rect 97120 5412 97176 5468
rect 97176 5412 97180 5468
rect 97116 5408 97180 5412
rect 97196 5468 97260 5472
rect 97196 5412 97200 5468
rect 97200 5412 97256 5468
rect 97256 5412 97260 5468
rect 97196 5408 97260 5412
rect 97276 5468 97340 5472
rect 97276 5412 97280 5468
rect 97280 5412 97336 5468
rect 97336 5412 97340 5468
rect 97276 5408 97340 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 39804 4524 39868 4588
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 66316 4380 66380 4384
rect 66316 4324 66320 4380
rect 66320 4324 66376 4380
rect 66376 4324 66380 4380
rect 66316 4320 66380 4324
rect 66396 4380 66460 4384
rect 66396 4324 66400 4380
rect 66400 4324 66456 4380
rect 66456 4324 66460 4380
rect 66396 4320 66460 4324
rect 66476 4380 66540 4384
rect 66476 4324 66480 4380
rect 66480 4324 66536 4380
rect 66536 4324 66540 4380
rect 66476 4320 66540 4324
rect 66556 4380 66620 4384
rect 66556 4324 66560 4380
rect 66560 4324 66616 4380
rect 66616 4324 66620 4380
rect 66556 4320 66620 4324
rect 97036 4380 97100 4384
rect 97036 4324 97040 4380
rect 97040 4324 97096 4380
rect 97096 4324 97100 4380
rect 97036 4320 97100 4324
rect 97116 4380 97180 4384
rect 97116 4324 97120 4380
rect 97120 4324 97176 4380
rect 97176 4324 97180 4380
rect 97116 4320 97180 4324
rect 97196 4380 97260 4384
rect 97196 4324 97200 4380
rect 97200 4324 97256 4380
rect 97256 4324 97260 4380
rect 97196 4320 97260 4324
rect 97276 4380 97340 4384
rect 97276 4324 97280 4380
rect 97280 4324 97336 4380
rect 97336 4324 97340 4380
rect 97276 4320 97340 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 66316 3292 66380 3296
rect 66316 3236 66320 3292
rect 66320 3236 66376 3292
rect 66376 3236 66380 3292
rect 66316 3232 66380 3236
rect 66396 3292 66460 3296
rect 66396 3236 66400 3292
rect 66400 3236 66456 3292
rect 66456 3236 66460 3292
rect 66396 3232 66460 3236
rect 66476 3292 66540 3296
rect 66476 3236 66480 3292
rect 66480 3236 66536 3292
rect 66536 3236 66540 3292
rect 66476 3232 66540 3236
rect 66556 3292 66620 3296
rect 66556 3236 66560 3292
rect 66560 3236 66616 3292
rect 66616 3236 66620 3292
rect 66556 3232 66620 3236
rect 97036 3292 97100 3296
rect 97036 3236 97040 3292
rect 97040 3236 97096 3292
rect 97096 3236 97100 3292
rect 97036 3232 97100 3236
rect 97116 3292 97180 3296
rect 97116 3236 97120 3292
rect 97120 3236 97176 3292
rect 97176 3236 97180 3292
rect 97116 3232 97180 3236
rect 97196 3292 97260 3296
rect 97196 3236 97200 3292
rect 97200 3236 97256 3292
rect 97256 3236 97260 3292
rect 97196 3232 97260 3236
rect 97276 3292 97340 3296
rect 97276 3236 97280 3292
rect 97280 3236 97336 3292
rect 97336 3236 97340 3292
rect 97276 3232 97340 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
rect 66316 2204 66380 2208
rect 66316 2148 66320 2204
rect 66320 2148 66376 2204
rect 66376 2148 66380 2204
rect 66316 2144 66380 2148
rect 66396 2204 66460 2208
rect 66396 2148 66400 2204
rect 66400 2148 66456 2204
rect 66456 2148 66460 2204
rect 66396 2144 66460 2148
rect 66476 2204 66540 2208
rect 66476 2148 66480 2204
rect 66480 2148 66536 2204
rect 66536 2148 66540 2204
rect 66476 2144 66540 2148
rect 66556 2204 66620 2208
rect 66556 2148 66560 2204
rect 66560 2148 66616 2204
rect 66616 2148 66620 2204
rect 66556 2144 66620 2148
rect 97036 2204 97100 2208
rect 97036 2148 97040 2204
rect 97040 2148 97096 2204
rect 97096 2148 97100 2204
rect 97036 2144 97100 2148
rect 97116 2204 97180 2208
rect 97116 2148 97120 2204
rect 97120 2148 97176 2204
rect 97176 2148 97180 2204
rect 97116 2144 97180 2148
rect 97196 2204 97260 2208
rect 97196 2148 97200 2204
rect 97200 2148 97256 2204
rect 97256 2148 97260 2204
rect 97196 2144 97260 2148
rect 97276 2204 97340 2208
rect 97276 2148 97280 2204
rect 97280 2148 97336 2204
rect 97336 2148 97340 2204
rect 97276 2144 97340 2148
<< metal4 >>
rect 4208 147456 4528 147472
rect 4208 147392 4216 147456
rect 4280 147392 4296 147456
rect 4360 147392 4376 147456
rect 4440 147392 4456 147456
rect 4520 147392 4528 147456
rect 4208 146368 4528 147392
rect 4208 146304 4216 146368
rect 4280 146304 4296 146368
rect 4360 146304 4376 146368
rect 4440 146304 4456 146368
rect 4520 146304 4528 146368
rect 4208 145280 4528 146304
rect 4208 145216 4216 145280
rect 4280 145216 4296 145280
rect 4360 145216 4376 145280
rect 4440 145216 4456 145280
rect 4520 145216 4528 145280
rect 4208 144192 4528 145216
rect 4208 144128 4216 144192
rect 4280 144128 4296 144192
rect 4360 144128 4376 144192
rect 4440 144128 4456 144192
rect 4520 144128 4528 144192
rect 4208 143104 4528 144128
rect 4208 143040 4216 143104
rect 4280 143040 4296 143104
rect 4360 143040 4376 143104
rect 4440 143040 4456 143104
rect 4520 143040 4528 143104
rect 4208 142016 4528 143040
rect 4208 141952 4216 142016
rect 4280 141952 4296 142016
rect 4360 141952 4376 142016
rect 4440 141952 4456 142016
rect 4520 141952 4528 142016
rect 4208 141218 4528 141952
rect 4208 140982 4250 141218
rect 4486 140982 4528 141218
rect 4208 140928 4528 140982
rect 4208 140864 4216 140928
rect 4280 140864 4296 140928
rect 4360 140864 4376 140928
rect 4440 140864 4456 140928
rect 4520 140864 4528 140928
rect 4208 139840 4528 140864
rect 4208 139776 4216 139840
rect 4280 139776 4296 139840
rect 4360 139776 4376 139840
rect 4440 139776 4456 139840
rect 4520 139776 4528 139840
rect 4208 138752 4528 139776
rect 4208 138688 4216 138752
rect 4280 138688 4296 138752
rect 4360 138688 4376 138752
rect 4440 138688 4456 138752
rect 4520 138688 4528 138752
rect 4208 137664 4528 138688
rect 4208 137600 4216 137664
rect 4280 137600 4296 137664
rect 4360 137600 4376 137664
rect 4440 137600 4456 137664
rect 4520 137600 4528 137664
rect 4208 136576 4528 137600
rect 4208 136512 4216 136576
rect 4280 136512 4296 136576
rect 4360 136512 4376 136576
rect 4440 136512 4456 136576
rect 4520 136512 4528 136576
rect 4208 135488 4528 136512
rect 4208 135424 4216 135488
rect 4280 135424 4296 135488
rect 4360 135424 4376 135488
rect 4440 135424 4456 135488
rect 4520 135424 4528 135488
rect 4208 134400 4528 135424
rect 4208 134336 4216 134400
rect 4280 134336 4296 134400
rect 4360 134336 4376 134400
rect 4440 134336 4456 134400
rect 4520 134336 4528 134400
rect 4208 133312 4528 134336
rect 4208 133248 4216 133312
rect 4280 133248 4296 133312
rect 4360 133248 4376 133312
rect 4440 133248 4456 133312
rect 4520 133248 4528 133312
rect 4208 132224 4528 133248
rect 4208 132160 4216 132224
rect 4280 132160 4296 132224
rect 4360 132160 4376 132224
rect 4440 132160 4456 132224
rect 4520 132160 4528 132224
rect 4208 131136 4528 132160
rect 4208 131072 4216 131136
rect 4280 131072 4296 131136
rect 4360 131072 4376 131136
rect 4440 131072 4456 131136
rect 4520 131072 4528 131136
rect 4208 130048 4528 131072
rect 4208 129984 4216 130048
rect 4280 129984 4296 130048
rect 4360 129984 4376 130048
rect 4440 129984 4456 130048
rect 4520 129984 4528 130048
rect 4208 128960 4528 129984
rect 4208 128896 4216 128960
rect 4280 128896 4296 128960
rect 4360 128896 4376 128960
rect 4440 128896 4456 128960
rect 4520 128896 4528 128960
rect 4208 128168 4528 128896
rect 4208 127932 4250 128168
rect 4486 127932 4528 128168
rect 4208 127872 4528 127932
rect 4208 127808 4216 127872
rect 4280 127808 4296 127872
rect 4360 127808 4376 127872
rect 4440 127808 4456 127872
rect 4520 127808 4528 127872
rect 4208 126784 4528 127808
rect 4208 126720 4216 126784
rect 4280 126720 4296 126784
rect 4360 126720 4376 126784
rect 4440 126720 4456 126784
rect 4520 126720 4528 126784
rect 4208 125696 4528 126720
rect 4208 125632 4216 125696
rect 4280 125632 4296 125696
rect 4360 125632 4376 125696
rect 4440 125632 4456 125696
rect 4520 125632 4528 125696
rect 4208 124608 4528 125632
rect 4208 124544 4216 124608
rect 4280 124544 4296 124608
rect 4360 124544 4376 124608
rect 4440 124544 4456 124608
rect 4520 124544 4528 124608
rect 4208 123520 4528 124544
rect 4208 123456 4216 123520
rect 4280 123456 4296 123520
rect 4360 123456 4376 123520
rect 4440 123456 4456 123520
rect 4520 123456 4528 123520
rect 4208 122432 4528 123456
rect 4208 122368 4216 122432
rect 4280 122368 4296 122432
rect 4360 122368 4376 122432
rect 4440 122368 4456 122432
rect 4520 122368 4528 122432
rect 4208 121344 4528 122368
rect 4208 121280 4216 121344
rect 4280 121280 4296 121344
rect 4360 121280 4376 121344
rect 4440 121280 4456 121344
rect 4520 121280 4528 121344
rect 4208 120256 4528 121280
rect 4208 120192 4216 120256
rect 4280 120192 4296 120256
rect 4360 120192 4376 120256
rect 4440 120192 4456 120256
rect 4520 120192 4528 120256
rect 4208 119168 4528 120192
rect 4208 119104 4216 119168
rect 4280 119104 4296 119168
rect 4360 119104 4376 119168
rect 4440 119104 4456 119168
rect 4520 119104 4528 119168
rect 4208 118080 4528 119104
rect 4208 118016 4216 118080
rect 4280 118016 4296 118080
rect 4360 118016 4376 118080
rect 4440 118016 4456 118080
rect 4520 118016 4528 118080
rect 4208 116992 4528 118016
rect 4208 116928 4216 116992
rect 4280 116928 4296 116992
rect 4360 116928 4376 116992
rect 4440 116928 4456 116992
rect 4520 116928 4528 116992
rect 4208 115904 4528 116928
rect 4208 115840 4216 115904
rect 4280 115840 4296 115904
rect 4360 115840 4376 115904
rect 4440 115840 4456 115904
rect 4520 115840 4528 115904
rect 4208 114816 4528 115840
rect 4208 114752 4216 114816
rect 4280 114752 4296 114816
rect 4360 114752 4376 114816
rect 4440 114752 4456 114816
rect 4520 114752 4528 114816
rect 4208 113728 4528 114752
rect 4208 113664 4216 113728
rect 4280 113664 4296 113728
rect 4360 113664 4376 113728
rect 4440 113664 4456 113728
rect 4520 113664 4528 113728
rect 4208 112640 4528 113664
rect 4208 112576 4216 112640
rect 4280 112576 4296 112640
rect 4360 112576 4376 112640
rect 4440 112576 4456 112640
rect 4520 112576 4528 112640
rect 4208 111552 4528 112576
rect 4208 111488 4216 111552
rect 4280 111488 4296 111552
rect 4360 111488 4376 111552
rect 4440 111488 4456 111552
rect 4520 111488 4528 111552
rect 4208 110464 4528 111488
rect 4208 110400 4216 110464
rect 4280 110400 4296 110464
rect 4360 110400 4376 110464
rect 4440 110400 4456 110464
rect 4520 110400 4528 110464
rect 4208 109376 4528 110400
rect 4208 109312 4216 109376
rect 4280 109312 4296 109376
rect 4360 109312 4376 109376
rect 4440 109312 4456 109376
rect 4520 109312 4528 109376
rect 4208 108288 4528 109312
rect 4208 108224 4216 108288
rect 4280 108224 4296 108288
rect 4360 108224 4376 108288
rect 4440 108224 4456 108288
rect 4520 108224 4528 108288
rect 4208 107200 4528 108224
rect 4208 107136 4216 107200
rect 4280 107136 4296 107200
rect 4360 107136 4376 107200
rect 4440 107136 4456 107200
rect 4520 107136 4528 107200
rect 4208 106112 4528 107136
rect 4208 106048 4216 106112
rect 4280 106048 4296 106112
rect 4360 106048 4376 106112
rect 4440 106048 4456 106112
rect 4520 106048 4528 106112
rect 4208 105024 4528 106048
rect 4208 104960 4216 105024
rect 4280 104960 4296 105024
rect 4360 104960 4376 105024
rect 4440 104960 4456 105024
rect 4520 104960 4528 105024
rect 4208 103936 4528 104960
rect 4208 103872 4216 103936
rect 4280 103872 4296 103936
rect 4360 103872 4376 103936
rect 4440 103872 4456 103936
rect 4520 103872 4528 103936
rect 4208 102848 4528 103872
rect 4208 102784 4216 102848
rect 4280 102784 4296 102848
rect 4360 102784 4376 102848
rect 4440 102784 4456 102848
rect 4520 102784 4528 102848
rect 4208 101760 4528 102784
rect 4208 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4528 101760
rect 4208 100672 4528 101696
rect 4208 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4528 100672
rect 4208 99584 4528 100608
rect 4208 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4528 99584
rect 4208 98496 4528 99520
rect 4208 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4528 98496
rect 4208 97532 4528 98432
rect 4208 97408 4250 97532
rect 4486 97408 4528 97532
rect 4208 97344 4216 97408
rect 4520 97344 4528 97408
rect 4208 97296 4250 97344
rect 4486 97296 4528 97344
rect 4208 96320 4528 97296
rect 4208 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4528 96320
rect 4208 95232 4528 96256
rect 4208 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4528 95232
rect 4208 94144 4528 95168
rect 4208 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4528 94144
rect 4208 93056 4528 94080
rect 4208 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4528 93056
rect 4208 91968 4528 92992
rect 4208 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4528 91968
rect 4208 90880 4528 91904
rect 4208 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4528 90880
rect 4208 89792 4528 90816
rect 4208 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4528 89792
rect 4208 88704 4528 89728
rect 4208 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4528 88704
rect 4208 87616 4528 88640
rect 4208 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4528 87616
rect 4208 86528 4528 87552
rect 4208 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4528 86528
rect 4208 85440 4528 86464
rect 4208 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4528 85440
rect 4208 84352 4528 85376
rect 4208 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4528 84352
rect 4208 83264 4528 84288
rect 4208 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4528 83264
rect 4208 82176 4528 83200
rect 4208 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4528 82176
rect 4208 81088 4528 82112
rect 4208 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4528 81088
rect 4208 80000 4528 81024
rect 4208 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4528 80000
rect 4208 78912 4528 79936
rect 4208 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4528 78912
rect 4208 77824 4528 78848
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 76736 4528 77760
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 75648 4528 76672
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 4208 74560 4528 75584
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 73472 4528 74496
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66896 4296 66944
rect 4360 66896 4376 66944
rect 4440 66896 4456 66944
rect 4520 66880 4528 66944
rect 4208 66660 4250 66880
rect 4486 66660 4528 66880
rect 4208 65856 4528 66660
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 146912 5188 147472
rect 4868 146848 4876 146912
rect 4940 146848 4956 146912
rect 5020 146848 5036 146912
rect 5100 146848 5116 146912
rect 5180 146848 5188 146912
rect 4868 145824 5188 146848
rect 4868 145760 4876 145824
rect 4940 145760 4956 145824
rect 5020 145760 5036 145824
rect 5100 145760 5116 145824
rect 5180 145760 5188 145824
rect 4868 144736 5188 145760
rect 4868 144672 4876 144736
rect 4940 144672 4956 144736
rect 5020 144672 5036 144736
rect 5100 144672 5116 144736
rect 5180 144672 5188 144736
rect 4868 143648 5188 144672
rect 4868 143584 4876 143648
rect 4940 143584 4956 143648
rect 5020 143584 5036 143648
rect 5100 143584 5116 143648
rect 5180 143584 5188 143648
rect 4868 142560 5188 143584
rect 4868 142496 4876 142560
rect 4940 142496 4956 142560
rect 5020 142496 5036 142560
rect 5100 142496 5116 142560
rect 5180 142496 5188 142560
rect 4868 141898 5188 142496
rect 4868 141662 4910 141898
rect 5146 141662 5188 141898
rect 4868 141472 5188 141662
rect 4868 141408 4876 141472
rect 4940 141408 4956 141472
rect 5020 141408 5036 141472
rect 5100 141408 5116 141472
rect 5180 141408 5188 141472
rect 4868 140384 5188 141408
rect 4868 140320 4876 140384
rect 4940 140320 4956 140384
rect 5020 140320 5036 140384
rect 5100 140320 5116 140384
rect 5180 140320 5188 140384
rect 4868 139296 5188 140320
rect 4868 139232 4876 139296
rect 4940 139232 4956 139296
rect 5020 139232 5036 139296
rect 5100 139232 5116 139296
rect 5180 139232 5188 139296
rect 4868 138208 5188 139232
rect 4868 138144 4876 138208
rect 4940 138144 4956 138208
rect 5020 138144 5036 138208
rect 5100 138144 5116 138208
rect 5180 138144 5188 138208
rect 4868 137120 5188 138144
rect 4868 137056 4876 137120
rect 4940 137056 4956 137120
rect 5020 137056 5036 137120
rect 5100 137056 5116 137120
rect 5180 137056 5188 137120
rect 4868 136032 5188 137056
rect 4868 135968 4876 136032
rect 4940 135968 4956 136032
rect 5020 135968 5036 136032
rect 5100 135968 5116 136032
rect 5180 135968 5188 136032
rect 4868 134944 5188 135968
rect 34928 147456 35248 147472
rect 34928 147392 34936 147456
rect 35000 147392 35016 147456
rect 35080 147392 35096 147456
rect 35160 147392 35176 147456
rect 35240 147392 35248 147456
rect 34928 146368 35248 147392
rect 34928 146304 34936 146368
rect 35000 146304 35016 146368
rect 35080 146304 35096 146368
rect 35160 146304 35176 146368
rect 35240 146304 35248 146368
rect 34928 145280 35248 146304
rect 34928 145216 34936 145280
rect 35000 145216 35016 145280
rect 35080 145216 35096 145280
rect 35160 145216 35176 145280
rect 35240 145216 35248 145280
rect 34928 144192 35248 145216
rect 34928 144128 34936 144192
rect 35000 144128 35016 144192
rect 35080 144128 35096 144192
rect 35160 144128 35176 144192
rect 35240 144128 35248 144192
rect 34928 143104 35248 144128
rect 34928 143040 34936 143104
rect 35000 143040 35016 143104
rect 35080 143040 35096 143104
rect 35160 143040 35176 143104
rect 35240 143040 35248 143104
rect 34928 142016 35248 143040
rect 34928 141952 34936 142016
rect 35000 141952 35016 142016
rect 35080 141952 35096 142016
rect 35160 141952 35176 142016
rect 35240 141952 35248 142016
rect 34928 141218 35248 141952
rect 34928 140982 34970 141218
rect 35206 140982 35248 141218
rect 34928 140928 35248 140982
rect 34928 140864 34936 140928
rect 35000 140864 35016 140928
rect 35080 140864 35096 140928
rect 35160 140864 35176 140928
rect 35240 140864 35248 140928
rect 34928 139840 35248 140864
rect 34928 139776 34936 139840
rect 35000 139776 35016 139840
rect 35080 139776 35096 139840
rect 35160 139776 35176 139840
rect 35240 139776 35248 139840
rect 34928 138752 35248 139776
rect 34928 138688 34936 138752
rect 35000 138688 35016 138752
rect 35080 138688 35096 138752
rect 35160 138688 35176 138752
rect 35240 138688 35248 138752
rect 34928 137664 35248 138688
rect 34928 137600 34936 137664
rect 35000 137600 35016 137664
rect 35080 137600 35096 137664
rect 35160 137600 35176 137664
rect 35240 137600 35248 137664
rect 34928 136576 35248 137600
rect 34928 136512 34936 136576
rect 35000 136512 35016 136576
rect 35080 136512 35096 136576
rect 35160 136512 35176 136576
rect 35240 136512 35248 136576
rect 34928 135650 35248 136512
rect 35588 146912 35908 147472
rect 35588 146848 35596 146912
rect 35660 146848 35676 146912
rect 35740 146848 35756 146912
rect 35820 146848 35836 146912
rect 35900 146848 35908 146912
rect 35588 145824 35908 146848
rect 35588 145760 35596 145824
rect 35660 145760 35676 145824
rect 35740 145760 35756 145824
rect 35820 145760 35836 145824
rect 35900 145760 35908 145824
rect 35588 144736 35908 145760
rect 35588 144672 35596 144736
rect 35660 144672 35676 144736
rect 35740 144672 35756 144736
rect 35820 144672 35836 144736
rect 35900 144672 35908 144736
rect 35588 143648 35908 144672
rect 35588 143584 35596 143648
rect 35660 143584 35676 143648
rect 35740 143584 35756 143648
rect 35820 143584 35836 143648
rect 35900 143584 35908 143648
rect 35588 142560 35908 143584
rect 35588 142496 35596 142560
rect 35660 142496 35676 142560
rect 35740 142496 35756 142560
rect 35820 142496 35836 142560
rect 35900 142496 35908 142560
rect 35588 141898 35908 142496
rect 35588 141662 35630 141898
rect 35866 141662 35908 141898
rect 35588 141472 35908 141662
rect 35588 141408 35596 141472
rect 35660 141408 35676 141472
rect 35740 141408 35756 141472
rect 35820 141408 35836 141472
rect 35900 141408 35908 141472
rect 35588 140384 35908 141408
rect 35588 140320 35596 140384
rect 35660 140320 35676 140384
rect 35740 140320 35756 140384
rect 35820 140320 35836 140384
rect 35900 140320 35908 140384
rect 35588 139296 35908 140320
rect 35588 139232 35596 139296
rect 35660 139232 35676 139296
rect 35740 139232 35756 139296
rect 35820 139232 35836 139296
rect 35900 139232 35908 139296
rect 35588 138208 35908 139232
rect 35588 138144 35596 138208
rect 35660 138144 35676 138208
rect 35740 138144 35756 138208
rect 35820 138144 35836 138208
rect 35900 138144 35908 138208
rect 35588 137120 35908 138144
rect 35588 137056 35596 137120
rect 35660 137056 35676 137120
rect 35740 137056 35756 137120
rect 35820 137056 35836 137120
rect 35900 137056 35908 137120
rect 35588 136032 35908 137056
rect 35588 135968 35596 136032
rect 35660 135968 35676 136032
rect 35740 135968 35756 136032
rect 35820 135968 35836 136032
rect 35900 135968 35908 136032
rect 35588 135650 35908 135968
rect 65648 147456 65968 147472
rect 65648 147392 65656 147456
rect 65720 147392 65736 147456
rect 65800 147392 65816 147456
rect 65880 147392 65896 147456
rect 65960 147392 65968 147456
rect 65648 146368 65968 147392
rect 65648 146304 65656 146368
rect 65720 146304 65736 146368
rect 65800 146304 65816 146368
rect 65880 146304 65896 146368
rect 65960 146304 65968 146368
rect 65648 145280 65968 146304
rect 65648 145216 65656 145280
rect 65720 145216 65736 145280
rect 65800 145216 65816 145280
rect 65880 145216 65896 145280
rect 65960 145216 65968 145280
rect 65648 144192 65968 145216
rect 65648 144128 65656 144192
rect 65720 144128 65736 144192
rect 65800 144128 65816 144192
rect 65880 144128 65896 144192
rect 65960 144128 65968 144192
rect 65648 143104 65968 144128
rect 65648 143040 65656 143104
rect 65720 143040 65736 143104
rect 65800 143040 65816 143104
rect 65880 143040 65896 143104
rect 65960 143040 65968 143104
rect 65648 142016 65968 143040
rect 65648 141952 65656 142016
rect 65720 141952 65736 142016
rect 65800 141952 65816 142016
rect 65880 141952 65896 142016
rect 65960 141952 65968 142016
rect 65648 141218 65968 141952
rect 65648 140982 65690 141218
rect 65926 140982 65968 141218
rect 65648 140928 65968 140982
rect 65648 140864 65656 140928
rect 65720 140864 65736 140928
rect 65800 140864 65816 140928
rect 65880 140864 65896 140928
rect 65960 140864 65968 140928
rect 65648 139840 65968 140864
rect 65648 139776 65656 139840
rect 65720 139776 65736 139840
rect 65800 139776 65816 139840
rect 65880 139776 65896 139840
rect 65960 139776 65968 139840
rect 65648 138752 65968 139776
rect 65648 138688 65656 138752
rect 65720 138688 65736 138752
rect 65800 138688 65816 138752
rect 65880 138688 65896 138752
rect 65960 138688 65968 138752
rect 65648 137664 65968 138688
rect 65648 137600 65656 137664
rect 65720 137600 65736 137664
rect 65800 137600 65816 137664
rect 65880 137600 65896 137664
rect 65960 137600 65968 137664
rect 65648 136576 65968 137600
rect 65648 136512 65656 136576
rect 65720 136512 65736 136576
rect 65800 136512 65816 136576
rect 65880 136512 65896 136576
rect 65960 136512 65968 136576
rect 65648 135834 65968 136512
rect 66308 146912 66628 147472
rect 66308 146848 66316 146912
rect 66380 146848 66396 146912
rect 66460 146848 66476 146912
rect 66540 146848 66556 146912
rect 66620 146848 66628 146912
rect 66308 145824 66628 146848
rect 66308 145760 66316 145824
rect 66380 145760 66396 145824
rect 66460 145760 66476 145824
rect 66540 145760 66556 145824
rect 66620 145760 66628 145824
rect 66308 144736 66628 145760
rect 66308 144672 66316 144736
rect 66380 144672 66396 144736
rect 66460 144672 66476 144736
rect 66540 144672 66556 144736
rect 66620 144672 66628 144736
rect 66308 143648 66628 144672
rect 66308 143584 66316 143648
rect 66380 143584 66396 143648
rect 66460 143584 66476 143648
rect 66540 143584 66556 143648
rect 66620 143584 66628 143648
rect 66308 142560 66628 143584
rect 66308 142496 66316 142560
rect 66380 142496 66396 142560
rect 66460 142496 66476 142560
rect 66540 142496 66556 142560
rect 66620 142496 66628 142560
rect 66308 141898 66628 142496
rect 66308 141662 66350 141898
rect 66586 141662 66628 141898
rect 66308 141472 66628 141662
rect 66308 141408 66316 141472
rect 66380 141408 66396 141472
rect 66460 141408 66476 141472
rect 66540 141408 66556 141472
rect 66620 141408 66628 141472
rect 66308 140384 66628 141408
rect 66308 140320 66316 140384
rect 66380 140320 66396 140384
rect 66460 140320 66476 140384
rect 66540 140320 66556 140384
rect 66620 140320 66628 140384
rect 66308 139296 66628 140320
rect 66308 139232 66316 139296
rect 66380 139232 66396 139296
rect 66460 139232 66476 139296
rect 66540 139232 66556 139296
rect 66620 139232 66628 139296
rect 66308 138208 66628 139232
rect 66308 138144 66316 138208
rect 66380 138144 66396 138208
rect 66460 138144 66476 138208
rect 66540 138144 66556 138208
rect 66620 138144 66628 138208
rect 66308 137120 66628 138144
rect 66308 137056 66316 137120
rect 66380 137056 66396 137120
rect 66460 137056 66476 137120
rect 66540 137056 66556 137120
rect 66620 137056 66628 137120
rect 66308 136032 66628 137056
rect 66308 135968 66316 136032
rect 66380 135968 66396 136032
rect 66460 135968 66476 136032
rect 66540 135968 66556 136032
rect 66620 135968 66628 136032
rect 66308 135650 66628 135968
rect 96368 147456 96688 147472
rect 96368 147392 96376 147456
rect 96440 147392 96456 147456
rect 96520 147392 96536 147456
rect 96600 147392 96616 147456
rect 96680 147392 96688 147456
rect 96368 146368 96688 147392
rect 96368 146304 96376 146368
rect 96440 146304 96456 146368
rect 96520 146304 96536 146368
rect 96600 146304 96616 146368
rect 96680 146304 96688 146368
rect 96368 145280 96688 146304
rect 96368 145216 96376 145280
rect 96440 145216 96456 145280
rect 96520 145216 96536 145280
rect 96600 145216 96616 145280
rect 96680 145216 96688 145280
rect 96368 144192 96688 145216
rect 96368 144128 96376 144192
rect 96440 144128 96456 144192
rect 96520 144128 96536 144192
rect 96600 144128 96616 144192
rect 96680 144128 96688 144192
rect 96368 143104 96688 144128
rect 96368 143040 96376 143104
rect 96440 143040 96456 143104
rect 96520 143040 96536 143104
rect 96600 143040 96616 143104
rect 96680 143040 96688 143104
rect 96368 142016 96688 143040
rect 96368 141952 96376 142016
rect 96440 141952 96456 142016
rect 96520 141952 96536 142016
rect 96600 141952 96616 142016
rect 96680 141952 96688 142016
rect 96368 141218 96688 141952
rect 96368 140982 96410 141218
rect 96646 140982 96688 141218
rect 96368 140928 96688 140982
rect 96368 140864 96376 140928
rect 96440 140864 96456 140928
rect 96520 140864 96536 140928
rect 96600 140864 96616 140928
rect 96680 140864 96688 140928
rect 96368 139840 96688 140864
rect 96368 139776 96376 139840
rect 96440 139776 96456 139840
rect 96520 139776 96536 139840
rect 96600 139776 96616 139840
rect 96680 139776 96688 139840
rect 96368 138752 96688 139776
rect 96368 138688 96376 138752
rect 96440 138688 96456 138752
rect 96520 138688 96536 138752
rect 96600 138688 96616 138752
rect 96680 138688 96688 138752
rect 96368 137664 96688 138688
rect 96368 137600 96376 137664
rect 96440 137600 96456 137664
rect 96520 137600 96536 137664
rect 96600 137600 96616 137664
rect 96680 137600 96688 137664
rect 96368 136576 96688 137600
rect 96368 136512 96376 136576
rect 96440 136512 96456 136576
rect 96520 136512 96536 136576
rect 96600 136512 96616 136576
rect 96680 136512 96688 136576
rect 95923 135692 95989 135693
rect 95923 135628 95924 135692
rect 95988 135628 95989 135692
rect 96368 135650 96688 136512
rect 97028 146912 97348 147472
rect 97028 146848 97036 146912
rect 97100 146848 97116 146912
rect 97180 146848 97196 146912
rect 97260 146848 97276 146912
rect 97340 146848 97348 146912
rect 97028 145824 97348 146848
rect 97028 145760 97036 145824
rect 97100 145760 97116 145824
rect 97180 145760 97196 145824
rect 97260 145760 97276 145824
rect 97340 145760 97348 145824
rect 97028 144736 97348 145760
rect 97028 144672 97036 144736
rect 97100 144672 97116 144736
rect 97180 144672 97196 144736
rect 97260 144672 97276 144736
rect 97340 144672 97348 144736
rect 97028 143648 97348 144672
rect 97028 143584 97036 143648
rect 97100 143584 97116 143648
rect 97180 143584 97196 143648
rect 97260 143584 97276 143648
rect 97340 143584 97348 143648
rect 97028 142560 97348 143584
rect 97028 142496 97036 142560
rect 97100 142496 97116 142560
rect 97180 142496 97196 142560
rect 97260 142496 97276 142560
rect 97340 142496 97348 142560
rect 97028 141898 97348 142496
rect 97028 141662 97070 141898
rect 97306 141662 97348 141898
rect 97028 141472 97348 141662
rect 97028 141408 97036 141472
rect 97100 141408 97116 141472
rect 97180 141408 97196 141472
rect 97260 141408 97276 141472
rect 97340 141408 97348 141472
rect 97028 140384 97348 141408
rect 97028 140320 97036 140384
rect 97100 140320 97116 140384
rect 97180 140320 97196 140384
rect 97260 140320 97276 140384
rect 97340 140320 97348 140384
rect 97028 139296 97348 140320
rect 97028 139232 97036 139296
rect 97100 139232 97116 139296
rect 97180 139232 97196 139296
rect 97260 139232 97276 139296
rect 97340 139232 97348 139296
rect 97028 138208 97348 139232
rect 97028 138144 97036 138208
rect 97100 138144 97116 138208
rect 97180 138144 97196 138208
rect 97260 138144 97276 138208
rect 97340 138144 97348 138208
rect 97028 137120 97348 138144
rect 97028 137056 97036 137120
rect 97100 137056 97116 137120
rect 97180 137056 97196 137120
rect 97260 137056 97276 137120
rect 97340 137056 97348 137120
rect 97028 136032 97348 137056
rect 97028 135968 97036 136032
rect 97100 135968 97116 136032
rect 97180 135968 97196 136032
rect 97260 135968 97276 136032
rect 97340 135968 97348 136032
rect 97028 135650 97348 135968
rect 105916 136576 106236 136592
rect 105916 136512 105924 136576
rect 105988 136512 106004 136576
rect 106068 136512 106084 136576
rect 106148 136512 106164 136576
rect 106228 136512 106236 136576
rect 95923 135627 95989 135628
rect 58571 135284 58637 135285
rect 58571 135220 58572 135284
rect 58636 135220 58637 135284
rect 58571 135219 58637 135220
rect 61147 135284 61213 135285
rect 61147 135220 61148 135284
rect 61212 135220 61213 135284
rect 61147 135219 61213 135220
rect 71083 135284 71149 135285
rect 71083 135220 71084 135284
rect 71148 135220 71149 135284
rect 71083 135219 71149 135220
rect 4868 134880 4876 134944
rect 4940 134880 4956 134944
rect 5020 134880 5036 134944
rect 5100 134880 5116 134944
rect 5180 134880 5188 134944
rect 4868 133856 5188 134880
rect 58574 134330 58634 135219
rect 61150 134330 61210 135219
rect 63539 135148 63605 135149
rect 63539 135084 63540 135148
rect 63604 135084 63605 135148
rect 63539 135083 63605 135084
rect 58541 134270 58634 134330
rect 61058 134270 61210 134330
rect 41066 134196 41132 134197
rect 41066 134132 41067 134196
rect 41131 134132 41132 134196
rect 41066 134131 41132 134132
rect 43562 134196 43628 134197
rect 43562 134132 43563 134196
rect 43627 134132 43628 134196
rect 43562 134131 43628 134132
rect 53546 134196 53612 134197
rect 53546 134132 53547 134196
rect 53611 134132 53612 134196
rect 53546 134131 53612 134132
rect 56042 134196 56108 134197
rect 56042 134132 56043 134196
rect 56107 134132 56108 134196
rect 56042 134131 56108 134132
rect 36074 133924 36140 133925
rect 36074 133860 36075 133924
rect 36139 133860 36140 133924
rect 36074 133859 36140 133860
rect 38570 133924 38636 133925
rect 38570 133860 38571 133924
rect 38635 133860 38636 133924
rect 38570 133859 38636 133860
rect 4868 133792 4876 133856
rect 4940 133792 4956 133856
rect 5020 133792 5036 133856
rect 5100 133792 5116 133856
rect 5180 133792 5188 133856
rect 4868 132768 5188 133792
rect 36077 133676 36137 133859
rect 38573 133676 38633 133859
rect 41069 133676 41129 134131
rect 43565 133676 43625 134131
rect 46059 133924 46125 133925
rect 46059 133860 46060 133924
rect 46124 133860 46125 133924
rect 46059 133859 46125 133860
rect 48543 133924 48609 133925
rect 48543 133860 48544 133924
rect 48608 133860 48609 133924
rect 48543 133859 48609 133860
rect 51050 133924 51116 133925
rect 51050 133860 51051 133924
rect 51115 133860 51116 133924
rect 51050 133859 51116 133860
rect 46062 133676 46122 133859
rect 48546 133676 48606 133859
rect 51053 133676 51113 133859
rect 53549 133676 53609 134131
rect 56045 133676 56105 134131
rect 58541 133676 58601 134270
rect 61058 133676 61118 134270
rect 63542 133676 63602 135083
rect 71086 134330 71146 135219
rect 73475 134468 73541 134469
rect 73475 134404 73476 134468
rect 73540 134404 73541 134468
rect 73475 134403 73541 134404
rect 71021 134270 71146 134330
rect 73478 134330 73538 134403
rect 95926 134330 95986 135627
rect 73478 134270 73577 134330
rect 66026 134196 66092 134197
rect 66026 134132 66027 134196
rect 66091 134132 66092 134196
rect 66026 134131 66092 134132
rect 66029 133676 66089 134131
rect 68522 133924 68588 133925
rect 68522 133860 68523 133924
rect 68587 133860 68588 133924
rect 68522 133859 68588 133860
rect 68525 133676 68585 133859
rect 71021 133676 71081 134270
rect 73517 133676 73577 134270
rect 95860 134270 95986 134330
rect 105916 135488 106236 136512
rect 105916 135424 105924 135488
rect 105988 135424 106004 135488
rect 106068 135424 106084 135488
rect 106148 135424 106164 135488
rect 106228 135424 106236 135488
rect 105916 134400 106236 135424
rect 105916 134336 105924 134400
rect 105988 134336 106004 134400
rect 106068 134336 106084 134400
rect 106148 134336 106164 134400
rect 106228 134336 106236 134400
rect 86141 133924 86207 133925
rect 86141 133860 86142 133924
rect 86206 133860 86207 133924
rect 86141 133859 86207 133860
rect 87309 133924 87375 133925
rect 87309 133860 87310 133924
rect 87374 133860 87375 133924
rect 87309 133859 87375 133860
rect 86144 133676 86204 133859
rect 87312 133676 87372 133859
rect 95860 133676 95920 134270
rect 4868 132704 4876 132768
rect 4940 132704 4956 132768
rect 5020 132704 5036 132768
rect 5100 132704 5116 132768
rect 5180 132704 5188 132768
rect 4868 131680 5188 132704
rect 4868 131616 4876 131680
rect 4940 131616 4956 131680
rect 5020 131616 5036 131680
rect 5100 131616 5116 131680
rect 5180 131616 5188 131680
rect 4868 130592 5188 131616
rect 4868 130528 4876 130592
rect 4940 130528 4956 130592
rect 5020 130528 5036 130592
rect 5100 130528 5116 130592
rect 5180 130528 5188 130592
rect 4868 129504 5188 130528
rect 4868 129440 4876 129504
rect 4940 129440 4956 129504
rect 5020 129440 5036 129504
rect 5100 129440 5116 129504
rect 5180 129440 5188 129504
rect 4868 128828 5188 129440
rect 105916 133312 106236 134336
rect 105916 133248 105924 133312
rect 105988 133248 106004 133312
rect 106068 133248 106084 133312
rect 106148 133248 106164 133312
rect 106228 133248 106236 133312
rect 105916 132224 106236 133248
rect 105916 132160 105924 132224
rect 105988 132160 106004 132224
rect 106068 132160 106084 132224
rect 106148 132160 106164 132224
rect 106228 132160 106236 132224
rect 105916 131136 106236 132160
rect 105916 131072 105924 131136
rect 105988 131072 106004 131136
rect 106068 131072 106084 131136
rect 106148 131072 106164 131136
rect 106228 131072 106236 131136
rect 105916 130048 106236 131072
rect 105916 129984 105924 130048
rect 105988 129984 106004 130048
rect 106068 129984 106084 130048
rect 106148 129984 106164 130048
rect 106228 129984 106236 130048
rect 105916 128960 106236 129984
rect 105916 128896 105924 128960
rect 105988 128896 106004 128960
rect 106068 128896 106084 128960
rect 106148 128896 106164 128960
rect 106228 128896 106236 128960
rect 4868 128592 4910 128828
rect 5146 128592 5188 128828
rect 4868 128416 5188 128592
rect 10696 128828 11044 128870
rect 10696 128592 10752 128828
rect 10988 128592 11044 128828
rect 10696 128550 11044 128592
rect 100936 128828 101284 128870
rect 100936 128592 100992 128828
rect 101228 128592 101284 128828
rect 100936 128550 101284 128592
rect 4868 128352 4876 128416
rect 4940 128352 4956 128416
rect 5020 128352 5036 128416
rect 5100 128352 5116 128416
rect 5180 128352 5188 128416
rect 4868 127328 5188 128352
rect 10000 128168 10348 128210
rect 10000 127932 10056 128168
rect 10292 127932 10348 128168
rect 10000 127890 10348 127932
rect 101632 128168 101980 128210
rect 101632 127932 101688 128168
rect 101924 127932 101980 128168
rect 101632 127890 101980 127932
rect 105916 128168 106236 128896
rect 105916 127932 105958 128168
rect 106194 127932 106236 128168
rect 4868 127264 4876 127328
rect 4940 127264 4956 127328
rect 5020 127264 5036 127328
rect 5100 127264 5116 127328
rect 5180 127264 5188 127328
rect 4868 126240 5188 127264
rect 4868 126176 4876 126240
rect 4940 126176 4956 126240
rect 5020 126176 5036 126240
rect 5100 126176 5116 126240
rect 5180 126176 5188 126240
rect 4868 125152 5188 126176
rect 4868 125088 4876 125152
rect 4940 125088 4956 125152
rect 5020 125088 5036 125152
rect 5100 125088 5116 125152
rect 5180 125088 5188 125152
rect 4868 124064 5188 125088
rect 4868 124000 4876 124064
rect 4940 124000 4956 124064
rect 5020 124000 5036 124064
rect 5100 124000 5116 124064
rect 5180 124000 5188 124064
rect 4868 122976 5188 124000
rect 4868 122912 4876 122976
rect 4940 122912 4956 122976
rect 5020 122912 5036 122976
rect 5100 122912 5116 122976
rect 5180 122912 5188 122976
rect 4868 121888 5188 122912
rect 4868 121824 4876 121888
rect 4940 121824 4956 121888
rect 5020 121824 5036 121888
rect 5100 121824 5116 121888
rect 5180 121824 5188 121888
rect 4868 120800 5188 121824
rect 4868 120736 4876 120800
rect 4940 120736 4956 120800
rect 5020 120736 5036 120800
rect 5100 120736 5116 120800
rect 5180 120736 5188 120800
rect 4868 119712 5188 120736
rect 4868 119648 4876 119712
rect 4940 119648 4956 119712
rect 5020 119648 5036 119712
rect 5100 119648 5116 119712
rect 5180 119648 5188 119712
rect 4868 118624 5188 119648
rect 4868 118560 4876 118624
rect 4940 118560 4956 118624
rect 5020 118560 5036 118624
rect 5100 118560 5116 118624
rect 5180 118560 5188 118624
rect 4868 117536 5188 118560
rect 4868 117472 4876 117536
rect 4940 117472 4956 117536
rect 5020 117472 5036 117536
rect 5100 117472 5116 117536
rect 5180 117472 5188 117536
rect 4868 116448 5188 117472
rect 4868 116384 4876 116448
rect 4940 116384 4956 116448
rect 5020 116384 5036 116448
rect 5100 116384 5116 116448
rect 5180 116384 5188 116448
rect 4868 115360 5188 116384
rect 4868 115296 4876 115360
rect 4940 115296 4956 115360
rect 5020 115296 5036 115360
rect 5100 115296 5116 115360
rect 5180 115296 5188 115360
rect 4868 114272 5188 115296
rect 4868 114208 4876 114272
rect 4940 114208 4956 114272
rect 5020 114208 5036 114272
rect 5100 114208 5116 114272
rect 5180 114208 5188 114272
rect 4868 113184 5188 114208
rect 4868 113120 4876 113184
rect 4940 113120 4956 113184
rect 5020 113120 5036 113184
rect 5100 113120 5116 113184
rect 5180 113120 5188 113184
rect 4868 112096 5188 113120
rect 4868 112032 4876 112096
rect 4940 112032 4956 112096
rect 5020 112032 5036 112096
rect 5100 112032 5116 112096
rect 5180 112032 5188 112096
rect 4868 111008 5188 112032
rect 4868 110944 4876 111008
rect 4940 110944 4956 111008
rect 5020 110944 5036 111008
rect 5100 110944 5116 111008
rect 5180 110944 5188 111008
rect 4868 109920 5188 110944
rect 4868 109856 4876 109920
rect 4940 109856 4956 109920
rect 5020 109856 5036 109920
rect 5100 109856 5116 109920
rect 5180 109856 5188 109920
rect 4868 108832 5188 109856
rect 4868 108768 4876 108832
rect 4940 108768 4956 108832
rect 5020 108768 5036 108832
rect 5100 108768 5116 108832
rect 5180 108768 5188 108832
rect 4868 107744 5188 108768
rect 4868 107680 4876 107744
rect 4940 107680 4956 107744
rect 5020 107680 5036 107744
rect 5100 107680 5116 107744
rect 5180 107680 5188 107744
rect 4868 106656 5188 107680
rect 4868 106592 4876 106656
rect 4940 106592 4956 106656
rect 5020 106592 5036 106656
rect 5100 106592 5116 106656
rect 5180 106592 5188 106656
rect 4868 105568 5188 106592
rect 4868 105504 4876 105568
rect 4940 105504 4956 105568
rect 5020 105504 5036 105568
rect 5100 105504 5116 105568
rect 5180 105504 5188 105568
rect 4868 104480 5188 105504
rect 4868 104416 4876 104480
rect 4940 104416 4956 104480
rect 5020 104416 5036 104480
rect 5100 104416 5116 104480
rect 5180 104416 5188 104480
rect 4868 103392 5188 104416
rect 4868 103328 4876 103392
rect 4940 103328 4956 103392
rect 5020 103328 5036 103392
rect 5100 103328 5116 103392
rect 5180 103328 5188 103392
rect 4868 102304 5188 103328
rect 4868 102240 4876 102304
rect 4940 102240 4956 102304
rect 5020 102240 5036 102304
rect 5100 102240 5116 102304
rect 5180 102240 5188 102304
rect 4868 101216 5188 102240
rect 4868 101152 4876 101216
rect 4940 101152 4956 101216
rect 5020 101152 5036 101216
rect 5100 101152 5116 101216
rect 5180 101152 5188 101216
rect 4868 100128 5188 101152
rect 4868 100064 4876 100128
rect 4940 100064 4956 100128
rect 5020 100064 5036 100128
rect 5100 100064 5116 100128
rect 5180 100064 5188 100128
rect 4868 99040 5188 100064
rect 4868 98976 4876 99040
rect 4940 98976 4956 99040
rect 5020 98976 5036 99040
rect 5100 98976 5116 99040
rect 5180 98976 5188 99040
rect 4868 98192 5188 98976
rect 105916 127872 106236 127932
rect 105916 127808 105924 127872
rect 105988 127808 106004 127872
rect 106068 127808 106084 127872
rect 106148 127808 106164 127872
rect 106228 127808 106236 127872
rect 105916 126784 106236 127808
rect 105916 126720 105924 126784
rect 105988 126720 106004 126784
rect 106068 126720 106084 126784
rect 106148 126720 106164 126784
rect 106228 126720 106236 126784
rect 105916 125696 106236 126720
rect 105916 125632 105924 125696
rect 105988 125632 106004 125696
rect 106068 125632 106084 125696
rect 106148 125632 106164 125696
rect 106228 125632 106236 125696
rect 105916 124608 106236 125632
rect 105916 124544 105924 124608
rect 105988 124544 106004 124608
rect 106068 124544 106084 124608
rect 106148 124544 106164 124608
rect 106228 124544 106236 124608
rect 105916 123520 106236 124544
rect 105916 123456 105924 123520
rect 105988 123456 106004 123520
rect 106068 123456 106084 123520
rect 106148 123456 106164 123520
rect 106228 123456 106236 123520
rect 105916 122432 106236 123456
rect 105916 122368 105924 122432
rect 105988 122368 106004 122432
rect 106068 122368 106084 122432
rect 106148 122368 106164 122432
rect 106228 122368 106236 122432
rect 105916 121344 106236 122368
rect 105916 121280 105924 121344
rect 105988 121280 106004 121344
rect 106068 121280 106084 121344
rect 106148 121280 106164 121344
rect 106228 121280 106236 121344
rect 105916 120256 106236 121280
rect 105916 120192 105924 120256
rect 105988 120192 106004 120256
rect 106068 120192 106084 120256
rect 106148 120192 106164 120256
rect 106228 120192 106236 120256
rect 105916 119168 106236 120192
rect 105916 119104 105924 119168
rect 105988 119104 106004 119168
rect 106068 119104 106084 119168
rect 106148 119104 106164 119168
rect 106228 119104 106236 119168
rect 105916 118080 106236 119104
rect 105916 118016 105924 118080
rect 105988 118016 106004 118080
rect 106068 118016 106084 118080
rect 106148 118016 106164 118080
rect 106228 118016 106236 118080
rect 105916 116992 106236 118016
rect 105916 116928 105924 116992
rect 105988 116928 106004 116992
rect 106068 116928 106084 116992
rect 106148 116928 106164 116992
rect 106228 116928 106236 116992
rect 105916 115904 106236 116928
rect 105916 115840 105924 115904
rect 105988 115840 106004 115904
rect 106068 115840 106084 115904
rect 106148 115840 106164 115904
rect 106228 115840 106236 115904
rect 105916 114816 106236 115840
rect 105916 114752 105924 114816
rect 105988 114752 106004 114816
rect 106068 114752 106084 114816
rect 106148 114752 106164 114816
rect 106228 114752 106236 114816
rect 105916 113728 106236 114752
rect 105916 113664 105924 113728
rect 105988 113664 106004 113728
rect 106068 113664 106084 113728
rect 106148 113664 106164 113728
rect 106228 113664 106236 113728
rect 105916 112640 106236 113664
rect 105916 112576 105924 112640
rect 105988 112576 106004 112640
rect 106068 112576 106084 112640
rect 106148 112576 106164 112640
rect 106228 112576 106236 112640
rect 105916 111552 106236 112576
rect 105916 111488 105924 111552
rect 105988 111488 106004 111552
rect 106068 111488 106084 111552
rect 106148 111488 106164 111552
rect 106228 111488 106236 111552
rect 105916 110464 106236 111488
rect 105916 110400 105924 110464
rect 105988 110400 106004 110464
rect 106068 110400 106084 110464
rect 106148 110400 106164 110464
rect 106228 110400 106236 110464
rect 105916 109376 106236 110400
rect 105916 109312 105924 109376
rect 105988 109312 106004 109376
rect 106068 109312 106084 109376
rect 106148 109312 106164 109376
rect 106228 109312 106236 109376
rect 105916 108288 106236 109312
rect 105916 108224 105924 108288
rect 105988 108224 106004 108288
rect 106068 108224 106084 108288
rect 106148 108224 106164 108288
rect 106228 108224 106236 108288
rect 105916 107200 106236 108224
rect 105916 107136 105924 107200
rect 105988 107136 106004 107200
rect 106068 107136 106084 107200
rect 106148 107136 106164 107200
rect 106228 107136 106236 107200
rect 105916 106112 106236 107136
rect 105916 106048 105924 106112
rect 105988 106048 106004 106112
rect 106068 106048 106084 106112
rect 106148 106048 106164 106112
rect 106228 106048 106236 106112
rect 105916 105024 106236 106048
rect 105916 104960 105924 105024
rect 105988 104960 106004 105024
rect 106068 104960 106084 105024
rect 106148 104960 106164 105024
rect 106228 104960 106236 105024
rect 105916 103936 106236 104960
rect 105916 103872 105924 103936
rect 105988 103872 106004 103936
rect 106068 103872 106084 103936
rect 106148 103872 106164 103936
rect 106228 103872 106236 103936
rect 105916 102848 106236 103872
rect 105916 102784 105924 102848
rect 105988 102784 106004 102848
rect 106068 102784 106084 102848
rect 106148 102784 106164 102848
rect 106228 102784 106236 102848
rect 105916 101760 106236 102784
rect 105916 101696 105924 101760
rect 105988 101696 106004 101760
rect 106068 101696 106084 101760
rect 106148 101696 106164 101760
rect 106228 101696 106236 101760
rect 105916 100672 106236 101696
rect 105916 100608 105924 100672
rect 105988 100608 106004 100672
rect 106068 100608 106084 100672
rect 106148 100608 106164 100672
rect 106228 100608 106236 100672
rect 105916 99584 106236 100608
rect 105916 99520 105924 99584
rect 105988 99520 106004 99584
rect 106068 99520 106084 99584
rect 106148 99520 106164 99584
rect 106228 99520 106236 99584
rect 105916 98496 106236 99520
rect 105916 98432 105924 98496
rect 105988 98432 106004 98496
rect 106068 98432 106084 98496
rect 106148 98432 106164 98496
rect 106228 98432 106236 98496
rect 4868 97956 4910 98192
rect 5146 97956 5188 98192
rect 4868 97952 5188 97956
rect 4868 97888 4876 97952
rect 4940 97888 4956 97952
rect 5020 97888 5036 97952
rect 5100 97888 5116 97952
rect 5180 97888 5188 97952
rect 10696 98192 11044 98234
rect 10696 97956 10752 98192
rect 10988 97956 11044 98192
rect 10696 97914 11044 97956
rect 100936 98192 101284 98234
rect 100936 97956 100992 98192
rect 101228 97956 101284 98192
rect 100936 97914 101284 97956
rect 4868 96864 5188 97888
rect 10000 97532 10348 97574
rect 10000 97296 10056 97532
rect 10292 97296 10348 97532
rect 10000 97254 10348 97296
rect 101632 97532 101980 97574
rect 101632 97296 101688 97532
rect 101924 97296 101980 97532
rect 101632 97254 101980 97296
rect 105916 97532 106236 98432
rect 105916 97408 105958 97532
rect 106194 97408 106236 97532
rect 105916 97344 105924 97408
rect 106228 97344 106236 97408
rect 105916 97296 105958 97344
rect 106194 97296 106236 97344
rect 4868 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5188 96864
rect 4868 95776 5188 96800
rect 4868 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5188 95776
rect 4868 94688 5188 95712
rect 4868 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5188 94688
rect 4868 93600 5188 94624
rect 4868 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5188 93600
rect 4868 92512 5188 93536
rect 105916 96320 106236 97296
rect 105916 96256 105924 96320
rect 105988 96256 106004 96320
rect 106068 96256 106084 96320
rect 106148 96256 106164 96320
rect 106228 96256 106236 96320
rect 105916 95232 106236 96256
rect 105916 95168 105924 95232
rect 105988 95168 106004 95232
rect 106068 95168 106084 95232
rect 106148 95168 106164 95232
rect 106228 95168 106236 95232
rect 105916 94144 106236 95168
rect 105916 94080 105924 94144
rect 105988 94080 106004 94144
rect 106068 94080 106084 94144
rect 106148 94080 106164 94144
rect 106228 94080 106236 94144
rect 102179 93392 102245 93393
rect 102179 93328 102180 93392
rect 102244 93328 102245 93392
rect 102179 93327 102245 93328
rect 4868 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5188 92512
rect 4868 91424 5188 92448
rect 4868 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5188 91424
rect 4868 90336 5188 91360
rect 4868 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5188 90336
rect 4868 89248 5188 90272
rect 4868 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5188 89248
rect 4868 88160 5188 89184
rect 4868 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5188 88160
rect 4868 87072 5188 88096
rect 4868 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5188 87072
rect 4868 85984 5188 87008
rect 4868 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5188 85984
rect 4868 84896 5188 85920
rect 4868 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5188 84896
rect 4868 83808 5188 84832
rect 4868 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5188 83808
rect 4868 82720 5188 83744
rect 4868 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5188 82720
rect 4868 81632 5188 82656
rect 4868 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5188 81632
rect 4868 80544 5188 81568
rect 4868 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5188 80544
rect 4868 79456 5188 80480
rect 16070 79933 16130 80038
rect 23440 79933 23500 80038
rect 16067 79932 16133 79933
rect 16067 79868 16068 79932
rect 16132 79868 16133 79932
rect 16067 79867 16133 79868
rect 23437 79932 23503 79933
rect 23437 79868 23438 79932
rect 23502 79868 23503 79932
rect 23437 79867 23503 79868
rect 24626 79525 24686 80038
rect 25776 79525 25836 80038
rect 26944 79525 27004 80038
rect 28122 79525 28182 80038
rect 29280 79525 29340 80038
rect 30448 79661 30508 80038
rect 31618 79661 31678 80038
rect 32784 79797 32844 80038
rect 32781 79796 32847 79797
rect 32781 79732 32782 79796
rect 32846 79732 32847 79796
rect 32781 79731 32847 79732
rect 30445 79660 30511 79661
rect 30445 79596 30446 79660
rect 30510 79596 30511 79660
rect 30445 79595 30511 79596
rect 31615 79660 31681 79661
rect 31615 79596 31616 79660
rect 31680 79596 31681 79660
rect 32784 79658 32844 79731
rect 32784 79598 32874 79658
rect 31615 79595 31681 79596
rect 24623 79524 24689 79525
rect 24623 79460 24624 79524
rect 24688 79460 24689 79524
rect 24623 79459 24689 79460
rect 25773 79524 25839 79525
rect 25773 79460 25774 79524
rect 25838 79460 25839 79524
rect 25773 79459 25839 79460
rect 26941 79524 27007 79525
rect 26941 79460 26942 79524
rect 27006 79460 27007 79524
rect 26941 79459 27007 79460
rect 28119 79524 28185 79525
rect 28119 79460 28120 79524
rect 28184 79460 28185 79524
rect 28119 79459 28185 79460
rect 29277 79524 29343 79525
rect 29277 79460 29278 79524
rect 29342 79460 29343 79524
rect 29277 79459 29343 79460
rect 4868 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5188 79456
rect 4868 78368 5188 79392
rect 32814 79117 32874 79598
rect 33952 79525 34012 80038
rect 35120 79525 35180 80038
rect 36288 79933 36348 80038
rect 36285 79932 36351 79933
rect 36285 79868 36286 79932
rect 36350 79868 36351 79932
rect 36285 79867 36351 79868
rect 37456 79661 37516 80038
rect 38624 79797 38684 80038
rect 39792 79933 39852 80038
rect 40960 79933 41020 80038
rect 39789 79932 39855 79933
rect 39789 79868 39790 79932
rect 39854 79868 39855 79932
rect 39789 79867 39855 79868
rect 40957 79932 41023 79933
rect 40957 79868 40958 79932
rect 41022 79868 41023 79932
rect 40957 79867 41023 79868
rect 38621 79796 38687 79797
rect 38621 79732 38622 79796
rect 38686 79732 38687 79796
rect 38621 79731 38687 79732
rect 37453 79660 37519 79661
rect 37453 79596 37454 79660
rect 37518 79596 37519 79660
rect 37453 79595 37519 79596
rect 42128 79525 42188 80038
rect 43296 79933 43356 80038
rect 43293 79932 43359 79933
rect 43293 79868 43294 79932
rect 43358 79868 43359 79932
rect 90529 79930 90589 80038
rect 43293 79867 43359 79868
rect 90406 79870 90589 79930
rect 33949 79524 34015 79525
rect 33949 79460 33950 79524
rect 34014 79460 34015 79524
rect 33949 79459 34015 79460
rect 35117 79524 35183 79525
rect 35117 79460 35118 79524
rect 35182 79460 35183 79524
rect 35117 79459 35183 79460
rect 42125 79524 42191 79525
rect 42125 79460 42126 79524
rect 42190 79460 42191 79524
rect 42125 79459 42191 79460
rect 32811 79116 32877 79117
rect 32811 79052 32812 79116
rect 32876 79052 32877 79116
rect 32811 79051 32877 79052
rect 4868 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5188 78368
rect 4868 77280 5188 78304
rect 4868 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5188 77280
rect 4868 76192 5188 77216
rect 4868 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5188 76192
rect 4868 75104 5188 76128
rect 4868 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5188 75104
rect 4868 74016 5188 75040
rect 4868 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5188 74016
rect 4868 72928 5188 73952
rect 4868 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5188 72928
rect 4868 71840 5188 72864
rect 4868 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5188 71840
rect 4868 70752 5188 71776
rect 4868 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5188 70752
rect 4868 69664 5188 70688
rect 4868 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5188 69664
rect 4868 68576 5188 69600
rect 4868 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5188 68576
rect 4868 67556 5188 68512
rect 4868 67488 4910 67556
rect 5146 67488 5188 67556
rect 4868 67424 4876 67488
rect 5180 67424 5188 67488
rect 4868 67320 4910 67424
rect 5146 67320 5188 67424
rect 4868 66400 5188 67320
rect 4868 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5188 66400
rect 4868 65312 5188 66336
rect 34928 77824 35248 77880
rect 34928 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35248 77824
rect 34928 76736 35248 77760
rect 34928 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35248 76736
rect 34928 75648 35248 76672
rect 34928 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35248 75648
rect 34928 74560 35248 75584
rect 34928 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35248 74560
rect 34928 73472 35248 74496
rect 34928 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35248 73472
rect 34928 72384 35248 73408
rect 34928 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35248 72384
rect 34928 71296 35248 72320
rect 34928 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35248 71296
rect 34928 70208 35248 71232
rect 34928 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35248 70208
rect 34928 69120 35248 70144
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66896 35016 66944
rect 35080 66896 35096 66944
rect 35160 66896 35176 66944
rect 35240 66880 35248 66944
rect 34928 66660 34970 66880
rect 35206 66660 35248 66880
rect 34928 65856 35248 66660
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 65650 35248 65792
rect 35588 77280 35908 78064
rect 35588 77216 35596 77280
rect 35660 77216 35676 77280
rect 35740 77216 35756 77280
rect 35820 77216 35836 77280
rect 35900 77216 35908 77280
rect 35588 76192 35908 77216
rect 35588 76128 35596 76192
rect 35660 76128 35676 76192
rect 35740 76128 35756 76192
rect 35820 76128 35836 76192
rect 35900 76128 35908 76192
rect 35588 75104 35908 76128
rect 35588 75040 35596 75104
rect 35660 75040 35676 75104
rect 35740 75040 35756 75104
rect 35820 75040 35836 75104
rect 35900 75040 35908 75104
rect 35588 74016 35908 75040
rect 35588 73952 35596 74016
rect 35660 73952 35676 74016
rect 35740 73952 35756 74016
rect 35820 73952 35836 74016
rect 35900 73952 35908 74016
rect 35588 72928 35908 73952
rect 35588 72864 35596 72928
rect 35660 72864 35676 72928
rect 35740 72864 35756 72928
rect 35820 72864 35836 72928
rect 35900 72864 35908 72928
rect 35588 71840 35908 72864
rect 35588 71776 35596 71840
rect 35660 71776 35676 71840
rect 35740 71776 35756 71840
rect 35820 71776 35836 71840
rect 35900 71776 35908 71840
rect 35588 70752 35908 71776
rect 35588 70688 35596 70752
rect 35660 70688 35676 70752
rect 35740 70688 35756 70752
rect 35820 70688 35836 70752
rect 35900 70688 35908 70752
rect 35588 69664 35908 70688
rect 65648 77824 65968 78064
rect 65648 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65968 77824
rect 65648 76736 65968 77760
rect 65648 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65968 76736
rect 65648 75648 65968 76672
rect 65648 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65968 75648
rect 65648 74560 65968 75584
rect 65648 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65968 74560
rect 65648 73472 65968 74496
rect 65648 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65968 73472
rect 65648 72384 65968 73408
rect 65648 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65968 72384
rect 65648 71296 65968 72320
rect 65648 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65968 71296
rect 65648 70208 65968 71232
rect 65648 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65968 70208
rect 63539 69868 63605 69869
rect 63539 69804 63540 69868
rect 63604 69804 63605 69868
rect 63539 69803 63605 69804
rect 35588 69600 35596 69664
rect 35660 69600 35676 69664
rect 35740 69600 35756 69664
rect 35820 69600 35836 69664
rect 35900 69600 35908 69664
rect 35588 68576 35908 69600
rect 61147 69324 61213 69325
rect 61147 69260 61148 69324
rect 61212 69260 61213 69324
rect 61147 69259 61213 69260
rect 53603 68780 53669 68781
rect 53603 68716 53604 68780
rect 53668 68716 53669 68780
rect 53603 68715 53669 68716
rect 35588 68512 35596 68576
rect 35660 68512 35676 68576
rect 35740 68512 35756 68576
rect 35820 68512 35836 68576
rect 35900 68512 35908 68576
rect 35588 67556 35908 68512
rect 48635 68236 48701 68237
rect 48635 68172 48636 68236
rect 48700 68172 48701 68236
rect 48635 68171 48701 68172
rect 35588 67488 35630 67556
rect 35866 67488 35908 67556
rect 35588 67424 35596 67488
rect 35900 67424 35908 67488
rect 35588 67320 35630 67424
rect 35866 67320 35908 67424
rect 35588 66400 35908 67320
rect 35588 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35908 66400
rect 35588 65650 35908 66336
rect 36123 65652 36189 65653
rect 36123 65588 36124 65652
rect 36188 65588 36189 65652
rect 36123 65587 36189 65588
rect 46059 65652 46125 65653
rect 46059 65588 46060 65652
rect 46124 65588 46125 65652
rect 46059 65587 46125 65588
rect 4868 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5188 65312
rect 4868 64224 5188 65248
rect 36126 64290 36186 65587
rect 38515 65516 38581 65517
rect 38515 65452 38516 65516
rect 38580 65452 38581 65516
rect 38515 65451 38581 65452
rect 4868 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5188 64224
rect 4868 63136 5188 64160
rect 36077 64230 36186 64290
rect 38518 64290 38578 65451
rect 41091 64292 41157 64293
rect 41091 64290 41092 64292
rect 38518 64230 38633 64290
rect 36077 63676 36137 64230
rect 38573 63676 38633 64230
rect 41069 64228 41092 64290
rect 41156 64228 41157 64292
rect 41069 64227 41157 64228
rect 41069 63676 41129 64227
rect 43562 64156 43628 64157
rect 43562 64092 43563 64156
rect 43627 64092 43628 64156
rect 43562 64091 43628 64092
rect 43565 63676 43625 64091
rect 46062 63676 46122 65587
rect 48638 64290 48698 68171
rect 53606 64290 53666 68715
rect 56179 68644 56245 68645
rect 56179 68580 56180 68644
rect 56244 68580 56245 68644
rect 56179 68579 56245 68580
rect 56182 64290 56242 68579
rect 61150 64290 61210 69259
rect 48557 64230 48698 64290
rect 53549 64230 53666 64290
rect 56045 64230 56242 64290
rect 61058 64230 61210 64290
rect 48557 63676 48617 64230
rect 51050 64156 51116 64157
rect 51050 64092 51051 64156
rect 51115 64092 51116 64156
rect 51050 64091 51116 64092
rect 51053 63676 51113 64091
rect 53549 63676 53609 64230
rect 56045 63676 56105 64230
rect 58538 64156 58604 64157
rect 58538 64092 58539 64156
rect 58603 64092 58604 64156
rect 58538 64091 58604 64092
rect 58541 63676 58601 64091
rect 61058 63676 61118 64230
rect 63542 63676 63602 69803
rect 65648 69120 65968 70144
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66896 65736 66944
rect 65800 66896 65816 66944
rect 65880 66896 65896 66944
rect 65960 66880 65968 66944
rect 65648 66660 65690 66880
rect 65926 66660 65968 66880
rect 65648 65856 65968 66660
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 65776 65968 65792
rect 66308 77280 66628 78064
rect 90406 77757 90466 79870
rect 90682 79250 90742 80038
rect 90816 79930 90876 80038
rect 90816 79870 91018 79930
rect 90682 79190 90834 79250
rect 90403 77756 90469 77757
rect 90403 77692 90404 77756
rect 90468 77692 90469 77756
rect 90403 77691 90469 77692
rect 90774 77485 90834 79190
rect 90958 77621 91018 79870
rect 96368 77824 96688 78064
rect 96368 77760 96376 77824
rect 96440 77760 96456 77824
rect 96520 77760 96536 77824
rect 96600 77760 96616 77824
rect 96680 77760 96688 77824
rect 90955 77620 91021 77621
rect 90955 77556 90956 77620
rect 91020 77556 91021 77620
rect 90955 77555 91021 77556
rect 90771 77484 90837 77485
rect 90771 77420 90772 77484
rect 90836 77420 90837 77484
rect 90771 77419 90837 77420
rect 66308 77216 66316 77280
rect 66380 77216 66396 77280
rect 66460 77216 66476 77280
rect 66540 77216 66556 77280
rect 66620 77216 66628 77280
rect 66308 76192 66628 77216
rect 66308 76128 66316 76192
rect 66380 76128 66396 76192
rect 66460 76128 66476 76192
rect 66540 76128 66556 76192
rect 66620 76128 66628 76192
rect 66308 75104 66628 76128
rect 66308 75040 66316 75104
rect 66380 75040 66396 75104
rect 66460 75040 66476 75104
rect 66540 75040 66556 75104
rect 66620 75040 66628 75104
rect 66308 74016 66628 75040
rect 66308 73952 66316 74016
rect 66380 73952 66396 74016
rect 66460 73952 66476 74016
rect 66540 73952 66556 74016
rect 66620 73952 66628 74016
rect 66308 72928 66628 73952
rect 66308 72864 66316 72928
rect 66380 72864 66396 72928
rect 66460 72864 66476 72928
rect 66540 72864 66556 72928
rect 66620 72864 66628 72928
rect 66308 71840 66628 72864
rect 96368 76736 96688 77760
rect 96368 76672 96376 76736
rect 96440 76672 96456 76736
rect 96520 76672 96536 76736
rect 96600 76672 96616 76736
rect 96680 76672 96688 76736
rect 96368 75648 96688 76672
rect 96368 75584 96376 75648
rect 96440 75584 96456 75648
rect 96520 75584 96536 75648
rect 96600 75584 96616 75648
rect 96680 75584 96688 75648
rect 96368 74560 96688 75584
rect 96368 74496 96376 74560
rect 96440 74496 96456 74560
rect 96520 74496 96536 74560
rect 96600 74496 96616 74560
rect 96680 74496 96688 74560
rect 96368 73472 96688 74496
rect 96368 73408 96376 73472
rect 96440 73408 96456 73472
rect 96520 73408 96536 73472
rect 96600 73408 96616 73472
rect 96680 73408 96688 73472
rect 86171 72588 86237 72589
rect 86171 72524 86172 72588
rect 86236 72524 86237 72588
rect 86171 72523 86237 72524
rect 66308 71776 66316 71840
rect 66380 71776 66396 71840
rect 66460 71776 66476 71840
rect 66540 71776 66556 71840
rect 66620 71776 66628 71840
rect 66308 70752 66628 71776
rect 66308 70688 66316 70752
rect 66380 70688 66396 70752
rect 66460 70688 66476 70752
rect 66540 70688 66556 70752
rect 66620 70688 66628 70752
rect 66308 69664 66628 70688
rect 73659 69868 73725 69869
rect 73659 69804 73660 69868
rect 73724 69804 73725 69868
rect 73659 69803 73725 69804
rect 66308 69600 66316 69664
rect 66380 69600 66396 69664
rect 66460 69600 66476 69664
rect 66540 69600 66556 69664
rect 66620 69600 66628 69664
rect 66308 68576 66628 69600
rect 66308 68512 66316 68576
rect 66380 68512 66396 68576
rect 66460 68512 66476 68576
rect 66540 68512 66556 68576
rect 66620 68512 66628 68576
rect 66308 67556 66628 68512
rect 66308 67488 66350 67556
rect 66586 67488 66628 67556
rect 66308 67424 66316 67488
rect 66620 67424 66628 67488
rect 66308 67320 66350 67424
rect 66586 67320 66628 67424
rect 66308 66400 66628 67320
rect 66308 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66628 66400
rect 66308 65650 66628 66336
rect 68507 66196 68573 66197
rect 68507 66132 68508 66196
rect 68572 66132 68573 66196
rect 68507 66131 68573 66132
rect 66026 64020 66092 64021
rect 66026 63956 66027 64020
rect 66091 63956 66092 64020
rect 66026 63955 66092 63956
rect 66029 63676 66089 63955
rect 68510 63676 68570 66131
rect 73662 64290 73722 69803
rect 86174 64290 86234 72523
rect 96368 72384 96688 73408
rect 96368 72320 96376 72384
rect 96440 72320 96456 72384
rect 96520 72320 96536 72384
rect 96600 72320 96616 72384
rect 96680 72320 96688 72384
rect 96368 71296 96688 72320
rect 96368 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96688 71296
rect 96368 70208 96688 71232
rect 96368 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96688 70208
rect 96368 69120 96688 70144
rect 96368 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96688 69120
rect 96368 68032 96688 69056
rect 96368 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96688 68032
rect 96368 66944 96688 67968
rect 96368 66880 96376 66944
rect 96440 66896 96456 66944
rect 96520 66896 96536 66944
rect 96600 66896 96616 66944
rect 96680 66880 96688 66944
rect 96368 66660 96410 66880
rect 96646 66660 96688 66880
rect 87275 65924 87341 65925
rect 87275 65860 87276 65924
rect 87340 65860 87341 65924
rect 87275 65859 87341 65860
rect 73517 64230 73722 64290
rect 86144 64230 86234 64290
rect 87278 64290 87338 65859
rect 96368 65856 96688 66660
rect 96368 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96688 65856
rect 96368 65650 96688 65792
rect 97028 77280 97348 78064
rect 97028 77216 97036 77280
rect 97100 77216 97116 77280
rect 97180 77216 97196 77280
rect 97260 77216 97276 77280
rect 97340 77216 97348 77280
rect 97028 76192 97348 77216
rect 97028 76128 97036 76192
rect 97100 76128 97116 76192
rect 97180 76128 97196 76192
rect 97260 76128 97276 76192
rect 97340 76128 97348 76192
rect 97028 75104 97348 76128
rect 97028 75040 97036 75104
rect 97100 75040 97116 75104
rect 97180 75040 97196 75104
rect 97260 75040 97276 75104
rect 97340 75040 97348 75104
rect 97028 74016 97348 75040
rect 97028 73952 97036 74016
rect 97100 73952 97116 74016
rect 97180 73952 97196 74016
rect 97260 73952 97276 74016
rect 97340 73952 97348 74016
rect 97028 72928 97348 73952
rect 97028 72864 97036 72928
rect 97100 72864 97116 72928
rect 97180 72864 97196 72928
rect 97260 72864 97276 72928
rect 97340 72864 97348 72928
rect 97028 71840 97348 72864
rect 97028 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97348 71840
rect 97028 70752 97348 71776
rect 97028 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97348 70752
rect 97028 69664 97348 70688
rect 102182 70410 102242 93327
rect 105916 93056 106236 94080
rect 105916 92992 105924 93056
rect 105988 92992 106004 93056
rect 106068 92992 106084 93056
rect 106148 92992 106164 93056
rect 106228 92992 106236 93056
rect 105916 91968 106236 92992
rect 105916 91904 105924 91968
rect 105988 91904 106004 91968
rect 106068 91904 106084 91968
rect 106148 91904 106164 91968
rect 106228 91904 106236 91968
rect 105916 90880 106236 91904
rect 105916 90816 105924 90880
rect 105988 90816 106004 90880
rect 106068 90816 106084 90880
rect 106148 90816 106164 90880
rect 106228 90816 106236 90880
rect 105916 89792 106236 90816
rect 105916 89728 105924 89792
rect 105988 89728 106004 89792
rect 106068 89728 106084 89792
rect 106148 89728 106164 89792
rect 106228 89728 106236 89792
rect 105916 88704 106236 89728
rect 105916 88640 105924 88704
rect 105988 88640 106004 88704
rect 106068 88640 106084 88704
rect 106148 88640 106164 88704
rect 106228 88640 106236 88704
rect 105916 87616 106236 88640
rect 105916 87552 105924 87616
rect 105988 87552 106004 87616
rect 106068 87552 106084 87616
rect 106148 87552 106164 87616
rect 106228 87552 106236 87616
rect 105916 86528 106236 87552
rect 105916 86464 105924 86528
rect 105988 86464 106004 86528
rect 106068 86464 106084 86528
rect 106148 86464 106164 86528
rect 106228 86464 106236 86528
rect 105916 85440 106236 86464
rect 105916 85376 105924 85440
rect 105988 85376 106004 85440
rect 106068 85376 106084 85440
rect 106148 85376 106164 85440
rect 106228 85376 106236 85440
rect 105916 84352 106236 85376
rect 105916 84288 105924 84352
rect 105988 84288 106004 84352
rect 106068 84288 106084 84352
rect 106148 84288 106164 84352
rect 106228 84288 106236 84352
rect 105916 83264 106236 84288
rect 105916 83200 105924 83264
rect 105988 83200 106004 83264
rect 106068 83200 106084 83264
rect 106148 83200 106164 83264
rect 106228 83200 106236 83264
rect 105916 82176 106236 83200
rect 105916 82112 105924 82176
rect 105988 82112 106004 82176
rect 106068 82112 106084 82176
rect 106148 82112 106164 82176
rect 106228 82112 106236 82176
rect 105916 81088 106236 82112
rect 105916 81024 105924 81088
rect 105988 81024 106004 81088
rect 106068 81024 106084 81088
rect 106148 81024 106164 81088
rect 106228 81024 106236 81088
rect 105916 80000 106236 81024
rect 105916 79936 105924 80000
rect 105988 79936 106004 80000
rect 106068 79936 106084 80000
rect 106148 79936 106164 80000
rect 106228 79936 106236 80000
rect 105916 78912 106236 79936
rect 105916 78848 105924 78912
rect 105988 78848 106004 78912
rect 106068 78848 106084 78912
rect 106148 78848 106164 78912
rect 106228 78848 106236 78912
rect 105916 77824 106236 78848
rect 105916 77760 105924 77824
rect 105988 77760 106004 77824
rect 106068 77760 106084 77824
rect 106148 77760 106164 77824
rect 106228 77760 106236 77824
rect 105916 77200 106236 77760
rect 106652 136032 106972 136592
rect 106652 135968 106660 136032
rect 106724 135968 106740 136032
rect 106804 135968 106820 136032
rect 106884 135968 106900 136032
rect 106964 135968 106972 136032
rect 106652 134944 106972 135968
rect 106652 134880 106660 134944
rect 106724 134880 106740 134944
rect 106804 134880 106820 134944
rect 106884 134880 106900 134944
rect 106964 134880 106972 134944
rect 106652 133856 106972 134880
rect 106652 133792 106660 133856
rect 106724 133792 106740 133856
rect 106804 133792 106820 133856
rect 106884 133792 106900 133856
rect 106964 133792 106972 133856
rect 106652 132768 106972 133792
rect 106652 132704 106660 132768
rect 106724 132704 106740 132768
rect 106804 132704 106820 132768
rect 106884 132704 106900 132768
rect 106964 132704 106972 132768
rect 106652 131680 106972 132704
rect 106652 131616 106660 131680
rect 106724 131616 106740 131680
rect 106804 131616 106820 131680
rect 106884 131616 106900 131680
rect 106964 131616 106972 131680
rect 106652 130592 106972 131616
rect 106652 130528 106660 130592
rect 106724 130528 106740 130592
rect 106804 130528 106820 130592
rect 106884 130528 106900 130592
rect 106964 130528 106972 130592
rect 106652 129504 106972 130528
rect 106652 129440 106660 129504
rect 106724 129440 106740 129504
rect 106804 129440 106820 129504
rect 106884 129440 106900 129504
rect 106964 129440 106972 129504
rect 106652 128828 106972 129440
rect 106652 128592 106694 128828
rect 106930 128592 106972 128828
rect 106652 128416 106972 128592
rect 106652 128352 106660 128416
rect 106724 128352 106740 128416
rect 106804 128352 106820 128416
rect 106884 128352 106900 128416
rect 106964 128352 106972 128416
rect 106652 127328 106972 128352
rect 106652 127264 106660 127328
rect 106724 127264 106740 127328
rect 106804 127264 106820 127328
rect 106884 127264 106900 127328
rect 106964 127264 106972 127328
rect 106652 126240 106972 127264
rect 106652 126176 106660 126240
rect 106724 126176 106740 126240
rect 106804 126176 106820 126240
rect 106884 126176 106900 126240
rect 106964 126176 106972 126240
rect 106652 125152 106972 126176
rect 106652 125088 106660 125152
rect 106724 125088 106740 125152
rect 106804 125088 106820 125152
rect 106884 125088 106900 125152
rect 106964 125088 106972 125152
rect 106652 124064 106972 125088
rect 106652 124000 106660 124064
rect 106724 124000 106740 124064
rect 106804 124000 106820 124064
rect 106884 124000 106900 124064
rect 106964 124000 106972 124064
rect 106652 122976 106972 124000
rect 106652 122912 106660 122976
rect 106724 122912 106740 122976
rect 106804 122912 106820 122976
rect 106884 122912 106900 122976
rect 106964 122912 106972 122976
rect 106652 121888 106972 122912
rect 106652 121824 106660 121888
rect 106724 121824 106740 121888
rect 106804 121824 106820 121888
rect 106884 121824 106900 121888
rect 106964 121824 106972 121888
rect 106652 120800 106972 121824
rect 106652 120736 106660 120800
rect 106724 120736 106740 120800
rect 106804 120736 106820 120800
rect 106884 120736 106900 120800
rect 106964 120736 106972 120800
rect 106652 119712 106972 120736
rect 106652 119648 106660 119712
rect 106724 119648 106740 119712
rect 106804 119648 106820 119712
rect 106884 119648 106900 119712
rect 106964 119648 106972 119712
rect 106652 118624 106972 119648
rect 106652 118560 106660 118624
rect 106724 118560 106740 118624
rect 106804 118560 106820 118624
rect 106884 118560 106900 118624
rect 106964 118560 106972 118624
rect 106652 117536 106972 118560
rect 106652 117472 106660 117536
rect 106724 117472 106740 117536
rect 106804 117472 106820 117536
rect 106884 117472 106900 117536
rect 106964 117472 106972 117536
rect 106652 116448 106972 117472
rect 106652 116384 106660 116448
rect 106724 116384 106740 116448
rect 106804 116384 106820 116448
rect 106884 116384 106900 116448
rect 106964 116384 106972 116448
rect 106652 115360 106972 116384
rect 106652 115296 106660 115360
rect 106724 115296 106740 115360
rect 106804 115296 106820 115360
rect 106884 115296 106900 115360
rect 106964 115296 106972 115360
rect 106652 114272 106972 115296
rect 106652 114208 106660 114272
rect 106724 114208 106740 114272
rect 106804 114208 106820 114272
rect 106884 114208 106900 114272
rect 106964 114208 106972 114272
rect 106652 113184 106972 114208
rect 106652 113120 106660 113184
rect 106724 113120 106740 113184
rect 106804 113120 106820 113184
rect 106884 113120 106900 113184
rect 106964 113120 106972 113184
rect 106652 112096 106972 113120
rect 106652 112032 106660 112096
rect 106724 112032 106740 112096
rect 106804 112032 106820 112096
rect 106884 112032 106900 112096
rect 106964 112032 106972 112096
rect 106652 111008 106972 112032
rect 106652 110944 106660 111008
rect 106724 110944 106740 111008
rect 106804 110944 106820 111008
rect 106884 110944 106900 111008
rect 106964 110944 106972 111008
rect 106652 109920 106972 110944
rect 106652 109856 106660 109920
rect 106724 109856 106740 109920
rect 106804 109856 106820 109920
rect 106884 109856 106900 109920
rect 106964 109856 106972 109920
rect 106652 108832 106972 109856
rect 106652 108768 106660 108832
rect 106724 108768 106740 108832
rect 106804 108768 106820 108832
rect 106884 108768 106900 108832
rect 106964 108768 106972 108832
rect 106652 107744 106972 108768
rect 106652 107680 106660 107744
rect 106724 107680 106740 107744
rect 106804 107680 106820 107744
rect 106884 107680 106900 107744
rect 106964 107680 106972 107744
rect 106652 106656 106972 107680
rect 106652 106592 106660 106656
rect 106724 106592 106740 106656
rect 106804 106592 106820 106656
rect 106884 106592 106900 106656
rect 106964 106592 106972 106656
rect 106652 105568 106972 106592
rect 106652 105504 106660 105568
rect 106724 105504 106740 105568
rect 106804 105504 106820 105568
rect 106884 105504 106900 105568
rect 106964 105504 106972 105568
rect 106652 104480 106972 105504
rect 106652 104416 106660 104480
rect 106724 104416 106740 104480
rect 106804 104416 106820 104480
rect 106884 104416 106900 104480
rect 106964 104416 106972 104480
rect 106652 103392 106972 104416
rect 106652 103328 106660 103392
rect 106724 103328 106740 103392
rect 106804 103328 106820 103392
rect 106884 103328 106900 103392
rect 106964 103328 106972 103392
rect 106652 102304 106972 103328
rect 106652 102240 106660 102304
rect 106724 102240 106740 102304
rect 106804 102240 106820 102304
rect 106884 102240 106900 102304
rect 106964 102240 106972 102304
rect 106652 101216 106972 102240
rect 106652 101152 106660 101216
rect 106724 101152 106740 101216
rect 106804 101152 106820 101216
rect 106884 101152 106900 101216
rect 106964 101152 106972 101216
rect 106652 100128 106972 101152
rect 106652 100064 106660 100128
rect 106724 100064 106740 100128
rect 106804 100064 106820 100128
rect 106884 100064 106900 100128
rect 106964 100064 106972 100128
rect 106652 99040 106972 100064
rect 106652 98976 106660 99040
rect 106724 98976 106740 99040
rect 106804 98976 106820 99040
rect 106884 98976 106900 99040
rect 106964 98976 106972 99040
rect 106652 98192 106972 98976
rect 106652 97956 106694 98192
rect 106930 97956 106972 98192
rect 106652 97952 106972 97956
rect 106652 97888 106660 97952
rect 106724 97888 106740 97952
rect 106804 97888 106820 97952
rect 106884 97888 106900 97952
rect 106964 97888 106972 97952
rect 106652 96864 106972 97888
rect 106652 96800 106660 96864
rect 106724 96800 106740 96864
rect 106804 96800 106820 96864
rect 106884 96800 106900 96864
rect 106964 96800 106972 96864
rect 106652 95776 106972 96800
rect 106652 95712 106660 95776
rect 106724 95712 106740 95776
rect 106804 95712 106820 95776
rect 106884 95712 106900 95776
rect 106964 95712 106972 95776
rect 106652 94688 106972 95712
rect 106652 94624 106660 94688
rect 106724 94624 106740 94688
rect 106804 94624 106820 94688
rect 106884 94624 106900 94688
rect 106964 94624 106972 94688
rect 106652 93600 106972 94624
rect 106652 93536 106660 93600
rect 106724 93536 106740 93600
rect 106804 93536 106820 93600
rect 106884 93536 106900 93600
rect 106964 93536 106972 93600
rect 106652 92512 106972 93536
rect 106652 92448 106660 92512
rect 106724 92448 106740 92512
rect 106804 92448 106820 92512
rect 106884 92448 106900 92512
rect 106964 92448 106972 92512
rect 106652 91424 106972 92448
rect 106652 91360 106660 91424
rect 106724 91360 106740 91424
rect 106804 91360 106820 91424
rect 106884 91360 106900 91424
rect 106964 91360 106972 91424
rect 106652 90336 106972 91360
rect 106652 90272 106660 90336
rect 106724 90272 106740 90336
rect 106804 90272 106820 90336
rect 106884 90272 106900 90336
rect 106964 90272 106972 90336
rect 106652 89248 106972 90272
rect 106652 89184 106660 89248
rect 106724 89184 106740 89248
rect 106804 89184 106820 89248
rect 106884 89184 106900 89248
rect 106964 89184 106972 89248
rect 106652 88160 106972 89184
rect 106652 88096 106660 88160
rect 106724 88096 106740 88160
rect 106804 88096 106820 88160
rect 106884 88096 106900 88160
rect 106964 88096 106972 88160
rect 106652 87072 106972 88096
rect 106652 87008 106660 87072
rect 106724 87008 106740 87072
rect 106804 87008 106820 87072
rect 106884 87008 106900 87072
rect 106964 87008 106972 87072
rect 106652 85984 106972 87008
rect 106652 85920 106660 85984
rect 106724 85920 106740 85984
rect 106804 85920 106820 85984
rect 106884 85920 106900 85984
rect 106964 85920 106972 85984
rect 106652 84896 106972 85920
rect 106652 84832 106660 84896
rect 106724 84832 106740 84896
rect 106804 84832 106820 84896
rect 106884 84832 106900 84896
rect 106964 84832 106972 84896
rect 106652 83808 106972 84832
rect 106652 83744 106660 83808
rect 106724 83744 106740 83808
rect 106804 83744 106820 83808
rect 106884 83744 106900 83808
rect 106964 83744 106972 83808
rect 106652 82720 106972 83744
rect 106652 82656 106660 82720
rect 106724 82656 106740 82720
rect 106804 82656 106820 82720
rect 106884 82656 106900 82720
rect 106964 82656 106972 82720
rect 106652 81632 106972 82656
rect 106652 81568 106660 81632
rect 106724 81568 106740 81632
rect 106804 81568 106820 81632
rect 106884 81568 106900 81632
rect 106964 81568 106972 81632
rect 106652 80544 106972 81568
rect 106652 80480 106660 80544
rect 106724 80480 106740 80544
rect 106804 80480 106820 80544
rect 106884 80480 106900 80544
rect 106964 80480 106972 80544
rect 106652 79456 106972 80480
rect 106652 79392 106660 79456
rect 106724 79392 106740 79456
rect 106804 79392 106820 79456
rect 106884 79392 106900 79456
rect 106964 79392 106972 79456
rect 106652 78368 106972 79392
rect 106652 78304 106660 78368
rect 106724 78304 106740 78368
rect 106804 78304 106820 78368
rect 106884 78304 106900 78368
rect 106964 78304 106972 78368
rect 106652 77280 106972 78304
rect 106652 77216 106660 77280
rect 106724 77216 106740 77280
rect 106804 77216 106820 77280
rect 106884 77216 106900 77280
rect 106964 77216 106972 77280
rect 106652 77200 106972 77216
rect 102182 70350 102794 70410
rect 97028 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97348 69664
rect 97028 68576 97348 69600
rect 102734 68917 102794 70350
rect 102731 68916 102797 68917
rect 102731 68852 102732 68916
rect 102796 68852 102797 68916
rect 102731 68851 102797 68852
rect 97028 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97348 68576
rect 97028 67556 97348 68512
rect 97028 67488 97070 67556
rect 97306 67488 97348 67556
rect 97028 67424 97036 67488
rect 97340 67424 97348 67488
rect 97028 67320 97070 67424
rect 97306 67320 97348 67424
rect 97028 66400 97348 67320
rect 97028 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97348 66400
rect 97028 65650 97348 66336
rect 87278 64230 87372 64290
rect 71018 63884 71084 63885
rect 71018 63820 71019 63884
rect 71083 63820 71084 63884
rect 71018 63819 71084 63820
rect 71021 63676 71081 63819
rect 73517 63676 73577 64230
rect 86144 63676 86204 64230
rect 87312 63676 87372 64230
rect 95857 64156 95923 64157
rect 95857 64092 95858 64156
rect 95922 64092 95923 64156
rect 95857 64091 95923 64092
rect 95860 63676 95920 64091
rect 4868 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5188 63136
rect 4868 62048 5188 63072
rect 4868 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5188 62048
rect 4868 60960 5188 61984
rect 4868 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5188 60960
rect 4868 59872 5188 60896
rect 4868 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5188 59872
rect 4868 58784 5188 59808
rect 4868 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5188 58784
rect 4868 57696 5188 58720
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 10696 36920 11044 36962
rect 10696 36684 10752 36920
rect 10988 36684 11044 36920
rect 10696 36642 11044 36684
rect 100936 36920 101284 36962
rect 100936 36684 100992 36920
rect 101228 36684 101284 36920
rect 100936 36642 101284 36684
rect 10000 36260 10348 36302
rect 10000 36024 10056 36260
rect 10292 36024 10348 36260
rect 10000 35982 10348 36024
rect 101632 36260 101980 36302
rect 101632 36024 101688 36260
rect 101924 36024 101980 36260
rect 101632 35982 101980 36024
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 102734 23493 102794 68851
rect 105916 65856 106236 66416
rect 105916 65792 105924 65856
rect 105988 65792 106004 65856
rect 106068 65792 106084 65856
rect 106148 65792 106164 65856
rect 106228 65792 106236 65856
rect 105916 64768 106236 65792
rect 105916 64704 105924 64768
rect 105988 64704 106004 64768
rect 106068 64704 106084 64768
rect 106148 64704 106164 64768
rect 106228 64704 106236 64768
rect 105916 63680 106236 64704
rect 105916 63616 105924 63680
rect 105988 63616 106004 63680
rect 106068 63616 106084 63680
rect 106148 63616 106164 63680
rect 106228 63616 106236 63680
rect 105916 62592 106236 63616
rect 105916 62528 105924 62592
rect 105988 62528 106004 62592
rect 106068 62528 106084 62592
rect 106148 62528 106164 62592
rect 106228 62528 106236 62592
rect 105916 61504 106236 62528
rect 105916 61440 105924 61504
rect 105988 61440 106004 61504
rect 106068 61440 106084 61504
rect 106148 61440 106164 61504
rect 106228 61440 106236 61504
rect 105916 60416 106236 61440
rect 105916 60352 105924 60416
rect 105988 60352 106004 60416
rect 106068 60352 106084 60416
rect 106148 60352 106164 60416
rect 106228 60352 106236 60416
rect 105916 59328 106236 60352
rect 105916 59264 105924 59328
rect 105988 59264 106004 59328
rect 106068 59264 106084 59328
rect 106148 59264 106164 59328
rect 106228 59264 106236 59328
rect 105916 58240 106236 59264
rect 105916 58176 105924 58240
rect 105988 58176 106004 58240
rect 106068 58176 106084 58240
rect 106148 58176 106164 58240
rect 106228 58176 106236 58240
rect 105916 57152 106236 58176
rect 105916 57088 105924 57152
rect 105988 57088 106004 57152
rect 106068 57088 106084 57152
rect 106148 57088 106164 57152
rect 106228 57088 106236 57152
rect 105916 56064 106236 57088
rect 105916 56000 105924 56064
rect 105988 56000 106004 56064
rect 106068 56000 106084 56064
rect 106148 56000 106164 56064
rect 106228 56000 106236 56064
rect 105916 54976 106236 56000
rect 105916 54912 105924 54976
rect 105988 54912 106004 54976
rect 106068 54912 106084 54976
rect 106148 54912 106164 54976
rect 106228 54912 106236 54976
rect 105916 53888 106236 54912
rect 105916 53824 105924 53888
rect 105988 53824 106004 53888
rect 106068 53824 106084 53888
rect 106148 53824 106164 53888
rect 106228 53824 106236 53888
rect 105916 52800 106236 53824
rect 105916 52736 105924 52800
rect 105988 52736 106004 52800
rect 106068 52736 106084 52800
rect 106148 52736 106164 52800
rect 106228 52736 106236 52800
rect 105916 51712 106236 52736
rect 105916 51648 105924 51712
rect 105988 51648 106004 51712
rect 106068 51648 106084 51712
rect 106148 51648 106164 51712
rect 106228 51648 106236 51712
rect 105916 50624 106236 51648
rect 105916 50560 105924 50624
rect 105988 50560 106004 50624
rect 106068 50560 106084 50624
rect 106148 50560 106164 50624
rect 106228 50560 106236 50624
rect 105916 49536 106236 50560
rect 105916 49472 105924 49536
rect 105988 49472 106004 49536
rect 106068 49472 106084 49536
rect 106148 49472 106164 49536
rect 106228 49472 106236 49536
rect 105916 48448 106236 49472
rect 105916 48384 105924 48448
rect 105988 48384 106004 48448
rect 106068 48384 106084 48448
rect 106148 48384 106164 48448
rect 106228 48384 106236 48448
rect 105916 47360 106236 48384
rect 105916 47296 105924 47360
rect 105988 47296 106004 47360
rect 106068 47296 106084 47360
rect 106148 47296 106164 47360
rect 106228 47296 106236 47360
rect 105916 46272 106236 47296
rect 105916 46208 105924 46272
rect 105988 46208 106004 46272
rect 106068 46208 106084 46272
rect 106148 46208 106164 46272
rect 106228 46208 106236 46272
rect 105916 45184 106236 46208
rect 105916 45120 105924 45184
rect 105988 45120 106004 45184
rect 106068 45120 106084 45184
rect 106148 45120 106164 45184
rect 106228 45120 106236 45184
rect 105916 44096 106236 45120
rect 105916 44032 105924 44096
rect 105988 44032 106004 44096
rect 106068 44032 106084 44096
rect 106148 44032 106164 44096
rect 106228 44032 106236 44096
rect 105916 43008 106236 44032
rect 105916 42944 105924 43008
rect 105988 42944 106004 43008
rect 106068 42944 106084 43008
rect 106148 42944 106164 43008
rect 106228 42944 106236 43008
rect 105916 41920 106236 42944
rect 105916 41856 105924 41920
rect 105988 41856 106004 41920
rect 106068 41856 106084 41920
rect 106148 41856 106164 41920
rect 106228 41856 106236 41920
rect 105916 40832 106236 41856
rect 105916 40768 105924 40832
rect 105988 40768 106004 40832
rect 106068 40768 106084 40832
rect 106148 40768 106164 40832
rect 106228 40768 106236 40832
rect 105916 39744 106236 40768
rect 105916 39680 105924 39744
rect 105988 39680 106004 39744
rect 106068 39680 106084 39744
rect 106148 39680 106164 39744
rect 106228 39680 106236 39744
rect 105916 38656 106236 39680
rect 105916 38592 105924 38656
rect 105988 38592 106004 38656
rect 106068 38592 106084 38656
rect 106148 38592 106164 38656
rect 106228 38592 106236 38656
rect 105916 37568 106236 38592
rect 105916 37504 105924 37568
rect 105988 37504 106004 37568
rect 106068 37504 106084 37568
rect 106148 37504 106164 37568
rect 106228 37504 106236 37568
rect 105916 36480 106236 37504
rect 105916 36416 105924 36480
rect 105988 36416 106004 36480
rect 106068 36416 106084 36480
rect 106148 36416 106164 36480
rect 106228 36416 106236 36480
rect 105916 36260 106236 36416
rect 105916 36024 105958 36260
rect 106194 36024 106236 36260
rect 105916 35392 106236 36024
rect 105916 35328 105924 35392
rect 105988 35328 106004 35392
rect 106068 35328 106084 35392
rect 106148 35328 106164 35392
rect 106228 35328 106236 35392
rect 105916 34304 106236 35328
rect 105916 34240 105924 34304
rect 105988 34240 106004 34304
rect 106068 34240 106084 34304
rect 106148 34240 106164 34304
rect 106228 34240 106236 34304
rect 105916 33216 106236 34240
rect 105916 33152 105924 33216
rect 105988 33152 106004 33216
rect 106068 33152 106084 33216
rect 106148 33152 106164 33216
rect 106228 33152 106236 33216
rect 105916 32128 106236 33152
rect 105916 32064 105924 32128
rect 105988 32064 106004 32128
rect 106068 32064 106084 32128
rect 106148 32064 106164 32128
rect 106228 32064 106236 32128
rect 105916 31040 106236 32064
rect 105916 30976 105924 31040
rect 105988 30976 106004 31040
rect 106068 30976 106084 31040
rect 106148 30976 106164 31040
rect 106228 30976 106236 31040
rect 105916 29952 106236 30976
rect 105916 29888 105924 29952
rect 105988 29888 106004 29952
rect 106068 29888 106084 29952
rect 106148 29888 106164 29952
rect 106228 29888 106236 29952
rect 105916 28864 106236 29888
rect 105916 28800 105924 28864
rect 105988 28800 106004 28864
rect 106068 28800 106084 28864
rect 106148 28800 106164 28864
rect 106228 28800 106236 28864
rect 105916 27776 106236 28800
rect 105916 27712 105924 27776
rect 105988 27712 106004 27776
rect 106068 27712 106084 27776
rect 106148 27712 106164 27776
rect 106228 27712 106236 27776
rect 105916 26688 106236 27712
rect 105916 26624 105924 26688
rect 105988 26624 106004 26688
rect 106068 26624 106084 26688
rect 106148 26624 106164 26688
rect 106228 26624 106236 26688
rect 105916 25600 106236 26624
rect 105916 25536 105924 25600
rect 105988 25536 106004 25600
rect 106068 25536 106084 25600
rect 106148 25536 106164 25600
rect 106228 25536 106236 25600
rect 105916 24512 106236 25536
rect 105916 24448 105924 24512
rect 105988 24448 106004 24512
rect 106068 24448 106084 24512
rect 106148 24448 106164 24512
rect 106228 24448 106236 24512
rect 102731 23492 102797 23493
rect 102731 23428 102732 23492
rect 102796 23428 102797 23492
rect 102731 23427 102797 23428
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 105916 23424 106236 24448
rect 105916 23360 105924 23424
rect 105988 23360 106004 23424
rect 106068 23360 106084 23424
rect 106148 23360 106164 23424
rect 106228 23360 106236 23424
rect 105916 22336 106236 23360
rect 105916 22272 105924 22336
rect 105988 22272 106004 22336
rect 106068 22272 106084 22336
rect 106148 22272 106164 22336
rect 106228 22272 106236 22336
rect 105916 21248 106236 22272
rect 105916 21184 105924 21248
rect 105988 21184 106004 21248
rect 106068 21184 106084 21248
rect 106148 21184 106164 21248
rect 106228 21184 106236 21248
rect 105916 20160 106236 21184
rect 105916 20096 105924 20160
rect 105988 20096 106004 20160
rect 106068 20096 106084 20160
rect 106148 20096 106164 20160
rect 106228 20096 106236 20160
rect 105916 19072 106236 20096
rect 105916 19008 105924 19072
rect 105988 19008 106004 19072
rect 106068 19008 106084 19072
rect 106148 19008 106164 19072
rect 106228 19008 106236 19072
rect 105916 17984 106236 19008
rect 105916 17920 105924 17984
rect 105988 17920 106004 17984
rect 106068 17920 106084 17984
rect 106148 17920 106164 17984
rect 106228 17920 106236 17984
rect 105916 16896 106236 17920
rect 105916 16832 105924 16896
rect 105988 16832 106004 16896
rect 106068 16832 106084 16896
rect 106148 16832 106164 16896
rect 106228 16832 106236 16896
rect 105916 15808 106236 16832
rect 105916 15744 105924 15808
rect 105988 15744 106004 15808
rect 106068 15744 106084 15808
rect 106148 15744 106164 15808
rect 106228 15744 106236 15808
rect 105916 14720 106236 15744
rect 105916 14656 105924 14720
rect 105988 14656 106004 14720
rect 106068 14656 106084 14720
rect 106148 14656 106164 14720
rect 106228 14656 106236 14720
rect 105916 13632 106236 14656
rect 105916 13568 105924 13632
rect 105988 13568 106004 13632
rect 106068 13568 106084 13632
rect 106148 13568 106164 13632
rect 106228 13568 106236 13632
rect 105916 12544 106236 13568
rect 105916 12480 105924 12544
rect 105988 12480 106004 12544
rect 106068 12480 106084 12544
rect 106148 12480 106164 12544
rect 106228 12480 106236 12544
rect 105916 11456 106236 12480
rect 105916 11392 105924 11456
rect 105988 11392 106004 11456
rect 106068 11392 106084 11456
rect 106148 11392 106164 11456
rect 106228 11392 106236 11456
rect 105916 10368 106236 11392
rect 105916 10304 105924 10368
rect 105988 10304 106004 10368
rect 106068 10304 106084 10368
rect 106148 10304 106164 10368
rect 106228 10304 106236 10368
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 16060 9621 16120 10038
rect 23440 9757 23500 10038
rect 23437 9756 23503 9757
rect 23437 9692 23438 9756
rect 23502 9692 23503 9756
rect 23437 9691 23503 9692
rect 24626 9621 24686 10038
rect 25776 9757 25836 10038
rect 25773 9756 25839 9757
rect 25773 9692 25774 9756
rect 25838 9692 25839 9756
rect 25773 9691 25839 9692
rect 16057 9620 16123 9621
rect 16057 9556 16058 9620
rect 16122 9556 16123 9620
rect 16057 9555 16123 9556
rect 24623 9620 24689 9621
rect 24623 9556 24624 9620
rect 24688 9556 24689 9620
rect 24623 9555 24689 9556
rect 26926 8941 26986 10038
rect 28122 9757 28182 10038
rect 29280 9757 29340 10038
rect 30448 9757 30508 10038
rect 28119 9756 28185 9757
rect 28119 9692 28120 9756
rect 28184 9692 28185 9756
rect 28119 9691 28185 9692
rect 29277 9756 29343 9757
rect 29277 9692 29278 9756
rect 29342 9692 29343 9756
rect 29277 9691 29343 9692
rect 30445 9756 30511 9757
rect 30445 9692 30446 9756
rect 30510 9692 30511 9756
rect 31618 9754 31678 10038
rect 32784 9754 32844 10038
rect 33952 9754 34012 10038
rect 35120 9890 35180 10038
rect 36288 9890 36348 10038
rect 37456 9890 37516 10038
rect 35120 9830 35266 9890
rect 36288 9830 36370 9890
rect 31618 9694 31770 9754
rect 32784 9694 32874 9754
rect 30445 9691 30511 9692
rect 26923 8940 26989 8941
rect 26923 8876 26924 8940
rect 26988 8876 26989 8940
rect 26923 8875 26989 8876
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 31710 8261 31770 9694
rect 32814 8261 32874 9694
rect 33918 9694 34012 9754
rect 33918 8261 33978 9694
rect 35206 8261 35266 9830
rect 36310 8261 36370 9830
rect 37414 9830 37516 9890
rect 38624 9890 38684 10038
rect 38624 9830 38762 9890
rect 37414 8261 37474 9830
rect 38702 8261 38762 9830
rect 31707 8260 31773 8261
rect 31707 8196 31708 8260
rect 31772 8196 31773 8260
rect 31707 8195 31773 8196
rect 32811 8260 32877 8261
rect 32811 8196 32812 8260
rect 32876 8196 32877 8260
rect 32811 8195 32877 8196
rect 33915 8260 33981 8261
rect 33915 8196 33916 8260
rect 33980 8196 33981 8260
rect 33915 8195 33981 8196
rect 35203 8260 35269 8261
rect 35203 8196 35204 8260
rect 35268 8196 35269 8260
rect 35203 8195 35269 8196
rect 36307 8260 36373 8261
rect 36307 8196 36308 8260
rect 36372 8196 36373 8260
rect 36307 8195 36373 8196
rect 37411 8260 37477 8261
rect 37411 8196 37412 8260
rect 37476 8196 37477 8260
rect 37411 8195 37477 8196
rect 38699 8260 38765 8261
rect 38699 8196 38700 8260
rect 38764 8196 38765 8260
rect 38699 8195 38765 8196
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 7104 35248 7880
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 7648 35908 8064
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 39806 4589 39866 10038
rect 40960 9890 41020 10038
rect 40910 9830 41020 9890
rect 42128 9890 42188 10038
rect 42128 9830 42258 9890
rect 40910 8261 40970 9830
rect 42198 8261 42258 9830
rect 43302 8261 43362 10038
rect 90529 9890 90589 10038
rect 90406 9830 90589 9890
rect 90406 8397 90466 9830
rect 90667 9621 90727 10038
rect 90816 9621 90876 10038
rect 90664 9620 90730 9621
rect 90664 9556 90665 9620
rect 90729 9556 90730 9620
rect 90664 9555 90730 9556
rect 90813 9620 90879 9621
rect 90813 9556 90814 9620
rect 90878 9556 90879 9620
rect 90813 9555 90879 9556
rect 105916 9280 106236 10304
rect 105916 9216 105924 9280
rect 105988 9216 106004 9280
rect 106068 9216 106084 9280
rect 106148 9216 106164 9280
rect 106228 9216 106236 9280
rect 90403 8396 90469 8397
rect 90403 8332 90404 8396
rect 90468 8332 90469 8396
rect 90403 8331 90469 8332
rect 40907 8260 40973 8261
rect 40907 8196 40908 8260
rect 40972 8196 40973 8260
rect 40907 8195 40973 8196
rect 42195 8260 42261 8261
rect 42195 8196 42196 8260
rect 42260 8196 42261 8260
rect 42195 8195 42261 8196
rect 43299 8260 43365 8261
rect 43299 8196 43300 8260
rect 43364 8196 43365 8260
rect 43299 8195 43365 8196
rect 105916 8192 106236 9216
rect 105916 8128 105924 8192
rect 105988 8128 106004 8192
rect 106068 8128 106084 8192
rect 106148 8128 106164 8192
rect 106228 8128 106236 8192
rect 65648 7104 65968 8064
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5624 65968 5952
rect 65648 5388 65690 5624
rect 65926 5388 65968 5624
rect 65648 4928 65968 5388
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 39803 4588 39869 4589
rect 39803 4524 39804 4588
rect 39868 4524 39869 4588
rect 39803 4523 39869 4524
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 66308 7648 66628 8064
rect 66308 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66628 7648
rect 66308 6560 66628 7584
rect 66308 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66628 6560
rect 66308 6284 66628 6496
rect 66308 6048 66350 6284
rect 66586 6048 66628 6284
rect 66308 5472 66628 6048
rect 66308 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66628 5472
rect 66308 4384 66628 5408
rect 66308 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66628 4384
rect 66308 3296 66628 4320
rect 66308 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66628 3296
rect 66308 2208 66628 3232
rect 66308 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66628 2208
rect 66308 2128 66628 2144
rect 96368 7104 96688 8064
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 5624 96688 5952
rect 96368 5388 96410 5624
rect 96646 5388 96688 5624
rect 96368 4928 96688 5388
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2128 96688 2688
rect 97028 7648 97348 8064
rect 97028 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97348 7648
rect 97028 6560 97348 7584
rect 105916 7104 106236 8128
rect 105916 7040 105924 7104
rect 105988 7040 106004 7104
rect 106068 7040 106084 7104
rect 106148 7040 106164 7104
rect 106228 7040 106236 7104
rect 105916 7024 106236 7040
rect 106652 66400 106972 66416
rect 106652 66336 106660 66400
rect 106724 66336 106740 66400
rect 106804 66336 106820 66400
rect 106884 66336 106900 66400
rect 106964 66336 106972 66400
rect 106652 65312 106972 66336
rect 106652 65248 106660 65312
rect 106724 65248 106740 65312
rect 106804 65248 106820 65312
rect 106884 65248 106900 65312
rect 106964 65248 106972 65312
rect 106652 64224 106972 65248
rect 106652 64160 106660 64224
rect 106724 64160 106740 64224
rect 106804 64160 106820 64224
rect 106884 64160 106900 64224
rect 106964 64160 106972 64224
rect 106652 63136 106972 64160
rect 106652 63072 106660 63136
rect 106724 63072 106740 63136
rect 106804 63072 106820 63136
rect 106884 63072 106900 63136
rect 106964 63072 106972 63136
rect 106652 62048 106972 63072
rect 106652 61984 106660 62048
rect 106724 61984 106740 62048
rect 106804 61984 106820 62048
rect 106884 61984 106900 62048
rect 106964 61984 106972 62048
rect 106652 60960 106972 61984
rect 106652 60896 106660 60960
rect 106724 60896 106740 60960
rect 106804 60896 106820 60960
rect 106884 60896 106900 60960
rect 106964 60896 106972 60960
rect 106652 59872 106972 60896
rect 106652 59808 106660 59872
rect 106724 59808 106740 59872
rect 106804 59808 106820 59872
rect 106884 59808 106900 59872
rect 106964 59808 106972 59872
rect 106652 58784 106972 59808
rect 106652 58720 106660 58784
rect 106724 58720 106740 58784
rect 106804 58720 106820 58784
rect 106884 58720 106900 58784
rect 106964 58720 106972 58784
rect 106652 57696 106972 58720
rect 106652 57632 106660 57696
rect 106724 57632 106740 57696
rect 106804 57632 106820 57696
rect 106884 57632 106900 57696
rect 106964 57632 106972 57696
rect 106652 56608 106972 57632
rect 106652 56544 106660 56608
rect 106724 56544 106740 56608
rect 106804 56544 106820 56608
rect 106884 56544 106900 56608
rect 106964 56544 106972 56608
rect 106652 55520 106972 56544
rect 106652 55456 106660 55520
rect 106724 55456 106740 55520
rect 106804 55456 106820 55520
rect 106884 55456 106900 55520
rect 106964 55456 106972 55520
rect 106652 54432 106972 55456
rect 106652 54368 106660 54432
rect 106724 54368 106740 54432
rect 106804 54368 106820 54432
rect 106884 54368 106900 54432
rect 106964 54368 106972 54432
rect 106652 53344 106972 54368
rect 106652 53280 106660 53344
rect 106724 53280 106740 53344
rect 106804 53280 106820 53344
rect 106884 53280 106900 53344
rect 106964 53280 106972 53344
rect 106652 52256 106972 53280
rect 106652 52192 106660 52256
rect 106724 52192 106740 52256
rect 106804 52192 106820 52256
rect 106884 52192 106900 52256
rect 106964 52192 106972 52256
rect 106652 51168 106972 52192
rect 106652 51104 106660 51168
rect 106724 51104 106740 51168
rect 106804 51104 106820 51168
rect 106884 51104 106900 51168
rect 106964 51104 106972 51168
rect 106652 50080 106972 51104
rect 106652 50016 106660 50080
rect 106724 50016 106740 50080
rect 106804 50016 106820 50080
rect 106884 50016 106900 50080
rect 106964 50016 106972 50080
rect 106652 48992 106972 50016
rect 106652 48928 106660 48992
rect 106724 48928 106740 48992
rect 106804 48928 106820 48992
rect 106884 48928 106900 48992
rect 106964 48928 106972 48992
rect 106652 47904 106972 48928
rect 106652 47840 106660 47904
rect 106724 47840 106740 47904
rect 106804 47840 106820 47904
rect 106884 47840 106900 47904
rect 106964 47840 106972 47904
rect 106652 46816 106972 47840
rect 106652 46752 106660 46816
rect 106724 46752 106740 46816
rect 106804 46752 106820 46816
rect 106884 46752 106900 46816
rect 106964 46752 106972 46816
rect 106652 45728 106972 46752
rect 106652 45664 106660 45728
rect 106724 45664 106740 45728
rect 106804 45664 106820 45728
rect 106884 45664 106900 45728
rect 106964 45664 106972 45728
rect 106652 44640 106972 45664
rect 106652 44576 106660 44640
rect 106724 44576 106740 44640
rect 106804 44576 106820 44640
rect 106884 44576 106900 44640
rect 106964 44576 106972 44640
rect 106652 43552 106972 44576
rect 106652 43488 106660 43552
rect 106724 43488 106740 43552
rect 106804 43488 106820 43552
rect 106884 43488 106900 43552
rect 106964 43488 106972 43552
rect 106652 42464 106972 43488
rect 106652 42400 106660 42464
rect 106724 42400 106740 42464
rect 106804 42400 106820 42464
rect 106884 42400 106900 42464
rect 106964 42400 106972 42464
rect 106652 41376 106972 42400
rect 106652 41312 106660 41376
rect 106724 41312 106740 41376
rect 106804 41312 106820 41376
rect 106884 41312 106900 41376
rect 106964 41312 106972 41376
rect 106652 40288 106972 41312
rect 106652 40224 106660 40288
rect 106724 40224 106740 40288
rect 106804 40224 106820 40288
rect 106884 40224 106900 40288
rect 106964 40224 106972 40288
rect 106652 39200 106972 40224
rect 106652 39136 106660 39200
rect 106724 39136 106740 39200
rect 106804 39136 106820 39200
rect 106884 39136 106900 39200
rect 106964 39136 106972 39200
rect 106652 38112 106972 39136
rect 106652 38048 106660 38112
rect 106724 38048 106740 38112
rect 106804 38048 106820 38112
rect 106884 38048 106900 38112
rect 106964 38048 106972 38112
rect 106652 37024 106972 38048
rect 106652 36960 106660 37024
rect 106724 36960 106740 37024
rect 106804 36960 106820 37024
rect 106884 36960 106900 37024
rect 106964 36960 106972 37024
rect 106652 36920 106972 36960
rect 106652 36684 106694 36920
rect 106930 36684 106972 36920
rect 106652 35936 106972 36684
rect 106652 35872 106660 35936
rect 106724 35872 106740 35936
rect 106804 35872 106820 35936
rect 106884 35872 106900 35936
rect 106964 35872 106972 35936
rect 106652 34848 106972 35872
rect 106652 34784 106660 34848
rect 106724 34784 106740 34848
rect 106804 34784 106820 34848
rect 106884 34784 106900 34848
rect 106964 34784 106972 34848
rect 106652 33760 106972 34784
rect 106652 33696 106660 33760
rect 106724 33696 106740 33760
rect 106804 33696 106820 33760
rect 106884 33696 106900 33760
rect 106964 33696 106972 33760
rect 106652 32672 106972 33696
rect 106652 32608 106660 32672
rect 106724 32608 106740 32672
rect 106804 32608 106820 32672
rect 106884 32608 106900 32672
rect 106964 32608 106972 32672
rect 106652 31584 106972 32608
rect 106652 31520 106660 31584
rect 106724 31520 106740 31584
rect 106804 31520 106820 31584
rect 106884 31520 106900 31584
rect 106964 31520 106972 31584
rect 106652 30496 106972 31520
rect 106652 30432 106660 30496
rect 106724 30432 106740 30496
rect 106804 30432 106820 30496
rect 106884 30432 106900 30496
rect 106964 30432 106972 30496
rect 106652 29408 106972 30432
rect 106652 29344 106660 29408
rect 106724 29344 106740 29408
rect 106804 29344 106820 29408
rect 106884 29344 106900 29408
rect 106964 29344 106972 29408
rect 106652 28320 106972 29344
rect 106652 28256 106660 28320
rect 106724 28256 106740 28320
rect 106804 28256 106820 28320
rect 106884 28256 106900 28320
rect 106964 28256 106972 28320
rect 106652 27232 106972 28256
rect 106652 27168 106660 27232
rect 106724 27168 106740 27232
rect 106804 27168 106820 27232
rect 106884 27168 106900 27232
rect 106964 27168 106972 27232
rect 106652 26144 106972 27168
rect 106652 26080 106660 26144
rect 106724 26080 106740 26144
rect 106804 26080 106820 26144
rect 106884 26080 106900 26144
rect 106964 26080 106972 26144
rect 106652 25056 106972 26080
rect 106652 24992 106660 25056
rect 106724 24992 106740 25056
rect 106804 24992 106820 25056
rect 106884 24992 106900 25056
rect 106964 24992 106972 25056
rect 106652 23968 106972 24992
rect 106652 23904 106660 23968
rect 106724 23904 106740 23968
rect 106804 23904 106820 23968
rect 106884 23904 106900 23968
rect 106964 23904 106972 23968
rect 106652 22880 106972 23904
rect 106652 22816 106660 22880
rect 106724 22816 106740 22880
rect 106804 22816 106820 22880
rect 106884 22816 106900 22880
rect 106964 22816 106972 22880
rect 106652 21792 106972 22816
rect 106652 21728 106660 21792
rect 106724 21728 106740 21792
rect 106804 21728 106820 21792
rect 106884 21728 106900 21792
rect 106964 21728 106972 21792
rect 106652 20704 106972 21728
rect 106652 20640 106660 20704
rect 106724 20640 106740 20704
rect 106804 20640 106820 20704
rect 106884 20640 106900 20704
rect 106964 20640 106972 20704
rect 106652 19616 106972 20640
rect 106652 19552 106660 19616
rect 106724 19552 106740 19616
rect 106804 19552 106820 19616
rect 106884 19552 106900 19616
rect 106964 19552 106972 19616
rect 106652 18528 106972 19552
rect 106652 18464 106660 18528
rect 106724 18464 106740 18528
rect 106804 18464 106820 18528
rect 106884 18464 106900 18528
rect 106964 18464 106972 18528
rect 106652 17440 106972 18464
rect 106652 17376 106660 17440
rect 106724 17376 106740 17440
rect 106804 17376 106820 17440
rect 106884 17376 106900 17440
rect 106964 17376 106972 17440
rect 106652 16352 106972 17376
rect 106652 16288 106660 16352
rect 106724 16288 106740 16352
rect 106804 16288 106820 16352
rect 106884 16288 106900 16352
rect 106964 16288 106972 16352
rect 106652 15264 106972 16288
rect 106652 15200 106660 15264
rect 106724 15200 106740 15264
rect 106804 15200 106820 15264
rect 106884 15200 106900 15264
rect 106964 15200 106972 15264
rect 106652 14176 106972 15200
rect 106652 14112 106660 14176
rect 106724 14112 106740 14176
rect 106804 14112 106820 14176
rect 106884 14112 106900 14176
rect 106964 14112 106972 14176
rect 106652 13088 106972 14112
rect 106652 13024 106660 13088
rect 106724 13024 106740 13088
rect 106804 13024 106820 13088
rect 106884 13024 106900 13088
rect 106964 13024 106972 13088
rect 106652 12000 106972 13024
rect 106652 11936 106660 12000
rect 106724 11936 106740 12000
rect 106804 11936 106820 12000
rect 106884 11936 106900 12000
rect 106964 11936 106972 12000
rect 106652 10912 106972 11936
rect 106652 10848 106660 10912
rect 106724 10848 106740 10912
rect 106804 10848 106820 10912
rect 106884 10848 106900 10912
rect 106964 10848 106972 10912
rect 106652 9824 106972 10848
rect 106652 9760 106660 9824
rect 106724 9760 106740 9824
rect 106804 9760 106820 9824
rect 106884 9760 106900 9824
rect 106964 9760 106972 9824
rect 106652 8736 106972 9760
rect 106652 8672 106660 8736
rect 106724 8672 106740 8736
rect 106804 8672 106820 8736
rect 106884 8672 106900 8736
rect 106964 8672 106972 8736
rect 106652 7648 106972 8672
rect 106652 7584 106660 7648
rect 106724 7584 106740 7648
rect 106804 7584 106820 7648
rect 106884 7584 106900 7648
rect 106964 7584 106972 7648
rect 106652 7024 106972 7584
rect 97028 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97348 6560
rect 97028 6284 97348 6496
rect 97028 6048 97070 6284
rect 97306 6048 97348 6284
rect 97028 5472 97348 6048
rect 97028 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97348 5472
rect 97028 4384 97348 5408
rect 97028 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97348 4384
rect 97028 3296 97348 4320
rect 97028 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97348 3296
rect 97028 2208 97348 3232
rect 97028 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97348 2208
rect 97028 2128 97348 2144
<< via4 >>
rect 4250 140982 4486 141218
rect 4250 127932 4486 128168
rect 4250 97408 4486 97532
rect 4250 97344 4280 97408
rect 4280 97344 4296 97408
rect 4296 97344 4360 97408
rect 4360 97344 4376 97408
rect 4376 97344 4440 97408
rect 4440 97344 4456 97408
rect 4456 97344 4486 97408
rect 4250 97296 4486 97344
rect 4250 66880 4280 66896
rect 4280 66880 4296 66896
rect 4296 66880 4360 66896
rect 4360 66880 4376 66896
rect 4376 66880 4440 66896
rect 4440 66880 4456 66896
rect 4456 66880 4486 66896
rect 4250 66660 4486 66880
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 141662 5146 141898
rect 34970 140982 35206 141218
rect 35630 141662 35866 141898
rect 65690 140982 65926 141218
rect 66350 141662 66586 141898
rect 96410 140982 96646 141218
rect 97070 141662 97306 141898
rect 4910 128592 5146 128828
rect 10752 128592 10988 128828
rect 100992 128592 101228 128828
rect 10056 127932 10292 128168
rect 101688 127932 101924 128168
rect 105958 127932 106194 128168
rect 4910 97956 5146 98192
rect 10752 97956 10988 98192
rect 100992 97956 101228 98192
rect 10056 97296 10292 97532
rect 101688 97296 101924 97532
rect 105958 97408 106194 97532
rect 105958 97344 105988 97408
rect 105988 97344 106004 97408
rect 106004 97344 106068 97408
rect 106068 97344 106084 97408
rect 106084 97344 106148 97408
rect 106148 97344 106164 97408
rect 106164 97344 106194 97408
rect 105958 97296 106194 97344
rect 4910 67488 5146 67556
rect 4910 67424 4940 67488
rect 4940 67424 4956 67488
rect 4956 67424 5020 67488
rect 5020 67424 5036 67488
rect 5036 67424 5100 67488
rect 5100 67424 5116 67488
rect 5116 67424 5146 67488
rect 4910 67320 5146 67424
rect 34970 66880 35000 66896
rect 35000 66880 35016 66896
rect 35016 66880 35080 66896
rect 35080 66880 35096 66896
rect 35096 66880 35160 66896
rect 35160 66880 35176 66896
rect 35176 66880 35206 66896
rect 34970 66660 35206 66880
rect 35630 67488 35866 67556
rect 35630 67424 35660 67488
rect 35660 67424 35676 67488
rect 35676 67424 35740 67488
rect 35740 67424 35756 67488
rect 35756 67424 35820 67488
rect 35820 67424 35836 67488
rect 35836 67424 35866 67488
rect 35630 67320 35866 67424
rect 65690 66880 65720 66896
rect 65720 66880 65736 66896
rect 65736 66880 65800 66896
rect 65800 66880 65816 66896
rect 65816 66880 65880 66896
rect 65880 66880 65896 66896
rect 65896 66880 65926 66896
rect 65690 66660 65926 66880
rect 66350 67488 66586 67556
rect 66350 67424 66380 67488
rect 66380 67424 66396 67488
rect 66396 67424 66460 67488
rect 66460 67424 66476 67488
rect 66476 67424 66540 67488
rect 66540 67424 66556 67488
rect 66556 67424 66586 67488
rect 66350 67320 66586 67424
rect 96410 66880 96440 66896
rect 96440 66880 96456 66896
rect 96456 66880 96520 66896
rect 96520 66880 96536 66896
rect 96536 66880 96600 66896
rect 96600 66880 96616 66896
rect 96616 66880 96646 66896
rect 96410 66660 96646 66880
rect 106694 128592 106930 128828
rect 106694 97956 106930 98192
rect 97070 67488 97306 67556
rect 97070 67424 97100 67488
rect 97100 67424 97116 67488
rect 97116 67424 97180 67488
rect 97180 67424 97196 67488
rect 97196 67424 97260 67488
rect 97260 67424 97276 67488
rect 97276 67424 97306 67488
rect 97070 67320 97306 67424
rect 4910 36684 5146 36920
rect 10752 36684 10988 36920
rect 100992 36684 101228 36920
rect 10056 36024 10292 36260
rect 101688 36024 101924 36260
rect 105958 36024 106194 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 6048 35866 6284
rect 65690 5388 65926 5624
rect 66350 6048 66586 6284
rect 96410 5388 96646 5624
rect 106694 36684 106930 36920
rect 97070 6048 97306 6284
<< metal5 >>
rect 4208 141898 108884 141940
rect 4208 141662 4910 141898
rect 5146 141662 35630 141898
rect 35866 141662 66350 141898
rect 66586 141662 97070 141898
rect 97306 141662 108884 141898
rect 4208 141620 108884 141662
rect 4208 141218 108884 141260
rect 4208 140982 4250 141218
rect 4486 140982 34970 141218
rect 35206 140982 65690 141218
rect 65926 140982 96410 141218
rect 96646 140982 108884 141218
rect 4208 140940 108884 140982
rect 1056 128828 108884 128870
rect 1056 128592 4910 128828
rect 5146 128592 10752 128828
rect 10988 128592 100992 128828
rect 101228 128592 106694 128828
rect 106930 128592 108884 128828
rect 1056 128550 108884 128592
rect 1056 128168 108884 128210
rect 1056 127932 4250 128168
rect 4486 127932 10056 128168
rect 10292 127932 101688 128168
rect 101924 127932 105958 128168
rect 106194 127932 108884 128168
rect 1056 127890 108884 127932
rect 1056 98192 108884 98234
rect 1056 97956 4910 98192
rect 5146 97956 10752 98192
rect 10988 97956 100992 98192
rect 101228 97956 106694 98192
rect 106930 97956 108884 98192
rect 1056 97914 108884 97956
rect 1056 97532 108884 97574
rect 1056 97296 4250 97532
rect 4486 97296 10056 97532
rect 10292 97296 101688 97532
rect 101924 97296 105958 97532
rect 106194 97296 108884 97532
rect 1056 97254 108884 97296
rect 1056 67556 108884 67598
rect 1056 67320 4910 67556
rect 5146 67320 35630 67556
rect 35866 67320 66350 67556
rect 66586 67320 97070 67556
rect 97306 67320 108884 67556
rect 1056 67278 108884 67320
rect 1056 66896 108884 66938
rect 1056 66660 4250 66896
rect 4486 66660 34970 66896
rect 35206 66660 65690 66896
rect 65926 66660 96410 66896
rect 96646 66660 108884 66896
rect 1056 66618 108884 66660
rect 1056 36920 108884 36962
rect 1056 36684 4910 36920
rect 5146 36684 10752 36920
rect 10988 36684 100992 36920
rect 101228 36684 106694 36920
rect 106930 36684 108884 36920
rect 1056 36642 108884 36684
rect 1056 36260 108884 36302
rect 1056 36024 4250 36260
rect 4486 36024 10056 36260
rect 10292 36024 101688 36260
rect 101924 36024 105958 36260
rect 106194 36024 108884 36260
rect 1056 35982 108884 36024
rect 1056 6284 108884 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 66350 6284
rect 66586 6048 97070 6284
rect 97306 6048 108884 6284
rect 1056 6006 108884 6048
rect 1056 5624 108884 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 65690 5624
rect 65926 5388 96410 5624
rect 96646 5388 108884 5624
rect 1056 5346 108884 5388
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1
transform -1 0 106352 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1
transform -1 0 105156 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1
transform -1 0 107824 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1
transform 1 0 102212 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1
transform 1 0 101292 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1
transform 1 0 101844 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _299_
timestamp 1
transform 1 0 100924 0 1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1
transform -1 0 24656 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _301_
timestamp 1
transform 1 0 102304 0 -1 73984
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _302_
timestamp 1
transform 1 0 102488 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _303_
timestamp 1
transform -1 0 103960 0 1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _304_
timestamp 1
transform 1 0 102764 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _305_
timestamp 1
transform 1 0 103040 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _306_
timestamp 1
transform -1 0 103500 0 1 75072
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _307_
timestamp 1
transform 1 0 104236 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _308_
timestamp 1
transform -1 0 104604 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _309_
timestamp 1
transform 1 0 103500 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _310_
timestamp 1
transform -1 0 103684 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _311_
timestamp 1
transform -1 0 104788 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _312_
timestamp 1
transform -1 0 104144 0 -1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _313_
timestamp 1
transform 1 0 105156 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _314_
timestamp 1
transform -1 0 104880 0 1 75072
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _315_
timestamp 1
transform -1 0 104420 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _316_
timestamp 1
transform 1 0 104420 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _317_
timestamp 1
transform -1 0 105892 0 -1 73984
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _318_
timestamp 1
transform 1 0 104420 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _319_
timestamp 1
transform -1 0 103776 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _320_
timestamp 1
transform -1 0 103040 0 -1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _321_
timestamp 1
transform 1 0 102856 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _322_
timestamp 1
transform 1 0 102764 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _323_
timestamp 1
transform -1 0 104880 0 -1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _324_
timestamp 1
transform -1 0 105432 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _325_
timestamp 1
transform -1 0 105432 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _326_
timestamp 1
transform 1 0 104972 0 -1 75072
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _327_
timestamp 1
transform 1 0 104880 0 1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _328_
timestamp 1
transform 1 0 104236 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _329_
timestamp 1
transform 1 0 101568 0 -1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _330_
timestamp 1
transform 1 0 105432 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _331_
timestamp 1
transform 1 0 105984 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _332_
timestamp 1
transform -1 0 105616 0 -1 71808
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _333_
timestamp 1
transform 1 0 105064 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _334_
timestamp 1
transform -1 0 105984 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _335_
timestamp 1
transform 1 0 106076 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _336_
timestamp 1
transform -1 0 106076 0 1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _337_
timestamp 1
transform -1 0 105616 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _338_
timestamp 1
transform -1 0 104052 0 -1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _339_
timestamp 1
transform -1 0 104052 0 -1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1
transform -1 0 98164 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _341_
timestamp 1
transform -1 0 104604 0 1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1
transform 1 0 103132 0 1 70720
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _343_
timestamp 1
transform 1 0 101752 0 -1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _344_
timestamp 1
transform -1 0 106444 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _345_
timestamp 1
transform -1 0 106076 0 -1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1
transform 1 0 104052 0 1 69632
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _347_
timestamp 1
transform -1 0 104052 0 -1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _348_
timestamp 1
transform -1 0 103592 0 -1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _349_
timestamp 1
transform 1 0 104972 0 -1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _350_
timestamp 1
transform -1 0 105432 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _351_
timestamp 1
transform -1 0 104144 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _352_
timestamp 1
transform 1 0 104880 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _353_
timestamp 1
transform -1 0 105524 0 1 68544
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _354_
timestamp 1
transform -1 0 105064 0 -1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _355_
timestamp 1
transform 1 0 104328 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _356_
timestamp 1
transform 1 0 102948 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _357_
timestamp 1
transform -1 0 104052 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _358_
timestamp 1
transform -1 0 102948 0 1 73984
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_2  _359_
timestamp 1
transform 1 0 101844 0 1 70720
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _360_
timestamp 1
transform -1 0 101384 0 1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _361_
timestamp 1
transform -1 0 102672 0 -1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _362_
timestamp 1
transform 1 0 102580 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _363_
timestamp 1
transform 1 0 102396 0 -1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _364_
timestamp 1
transform 1 0 103132 0 1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _365_
timestamp 1
transform 1 0 103868 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _366_
timestamp 1
transform 1 0 104420 0 1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _367_
timestamp 1
transform -1 0 103132 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _368_
timestamp 1
transform -1 0 104420 0 1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _369_
timestamp 1
transform -1 0 103960 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _370_
timestamp 1
transform 1 0 102948 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _371_
timestamp 1
transform -1 0 101568 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _372_
timestamp 1
transform -1 0 103500 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _373_
timestamp 1
transform -1 0 104880 0 -1 68544
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _374_
timestamp 1
transform 1 0 102488 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _375_
timestamp 1
transform 1 0 101660 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1
transform -1 0 101476 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _377_
timestamp 1
transform -1 0 102212 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _378_
timestamp 1
transform 1 0 102304 0 1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _379_
timestamp 1
transform -1 0 102212 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _380_
timestamp 1
transform -1 0 101384 0 -1 68544
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _381_
timestamp 1
transform -1 0 102212 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _382_
timestamp 1
transform 1 0 101660 0 1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _383_
timestamp 1
transform -1 0 100556 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1
transform -1 0 98440 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _385_
timestamp 1
transform 1 0 100188 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1
transform 1 0 100188 0 1 66368
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _387_
timestamp 1
transform -1 0 100556 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _388_
timestamp 1
transform -1 0 100832 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _389_
timestamp 1
transform 1 0 100372 0 1 68544
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _390_
timestamp 1
transform 1 0 101384 0 -1 68544
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _391_
timestamp 1
transform 1 0 99360 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _392_
timestamp 1
transform 1 0 98808 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _393_
timestamp 1
transform -1 0 99360 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _394_
timestamp 1
transform -1 0 98808 0 1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _395_
timestamp 1
transform 1 0 98348 0 -1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _396_
timestamp 1
transform 1 0 99636 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _397_
timestamp 1
transform 1 0 100556 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _398_
timestamp 1
transform 1 0 101660 0 1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _399_
timestamp 1
transform 1 0 101660 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1
transform 1 0 101660 0 1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _401_
timestamp 1
transform 1 0 99452 0 -1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _402_
timestamp 1
transform 1 0 98072 0 1 66368
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _403_
timestamp 1
transform -1 0 100188 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _404_
timestamp 1
transform 1 0 99084 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1
transform -1 0 100372 0 1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _406_
timestamp 1
transform 1 0 100188 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _407_
timestamp 1
transform -1 0 101200 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _408_
timestamp 1
transform -1 0 100280 0 1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _409_
timestamp 1
transform -1 0 97796 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _410_
timestamp 1
transform 1 0 97060 0 1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1
transform -1 0 98256 0 -1 68544
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _412_
timestamp 1
transform 1 0 97704 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _413_
timestamp 1
transform 1 0 98440 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_2  _414_
timestamp 1
transform 1 0 99084 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _415_
timestamp 1
transform -1 0 99728 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _416_
timestamp 1
transform -1 0 98992 0 -1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _417_
timestamp 1
transform 1 0 97796 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _418_
timestamp 1
transform 1 0 97612 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _419_
timestamp 1
transform 1 0 96508 0 1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _420_
timestamp 1
transform 1 0 98440 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _421_
timestamp 1
transform 1 0 96508 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _422_
timestamp 1
transform -1 0 98808 0 -1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _423_
timestamp 1
transform -1 0 98992 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _424_
timestamp 1
transform 1 0 95864 0 -1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1
transform -1 0 98164 0 -1 70720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1
transform 1 0 98624 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _427_
timestamp 1
transform 1 0 97796 0 -1 71808
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _428_
timestamp 1
transform 1 0 96232 0 -1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _429_
timestamp 1
transform 1 0 99268 0 -1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _430_
timestamp 1
transform 1 0 98900 0 1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _431_
timestamp 1
transform 1 0 99360 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _432_
timestamp 1
transform -1 0 99636 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _433_
timestamp 1
transform -1 0 99544 0 -1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _434_
timestamp 1
transform -1 0 101292 0 -1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _435_
timestamp 1
transform 1 0 99544 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _436_
timestamp 1
transform -1 0 98808 0 -1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _437_
timestamp 1
transform -1 0 97336 0 -1 71808
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _438_
timestamp 1
transform 1 0 96508 0 1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _439_
timestamp 1
transform -1 0 98072 0 1 71808
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _440_
timestamp 1
transform -1 0 98808 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _441_
timestamp 1
transform 1 0 99820 0 1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _442_
timestamp 1
transform -1 0 101108 0 -1 71808
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1
transform 1 0 100004 0 -1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _444_
timestamp 1
transform 1 0 100372 0 -1 76160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _445_
timestamp 1
transform 1 0 100280 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _446_
timestamp 1
transform 1 0 101108 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _447_
timestamp 1
transform -1 0 100556 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _448_
timestamp 1
transform 1 0 101016 0 1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp 1
transform 1 0 101660 0 1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _450_
timestamp 1
transform 1 0 102120 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _451_
timestamp 1
transform -1 0 102304 0 1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _452_
timestamp 1
transform 1 0 101568 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _453_
timestamp 1
transform 1 0 101568 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _454_
timestamp 1
transform -1 0 100188 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _455_
timestamp 1
transform 1 0 100464 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _456_
timestamp 1
transform 1 0 97612 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _457_
timestamp 1
transform -1 0 98624 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _458_
timestamp 1
transform -1 0 99268 0 1 71808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _459_
timestamp 1
transform -1 0 99912 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _460_
timestamp 1
transform 1 0 100832 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _461_
timestamp 1
transform -1 0 102304 0 1 75072
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1
transform 1 0 100740 0 1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _463_
timestamp 1
transform -1 0 99360 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _464_
timestamp 1
transform -1 0 100832 0 -1 75072
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _465_
timestamp 1
transform -1 0 101016 0 1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _466_
timestamp 1
transform 1 0 99912 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _467_
timestamp 1
transform -1 0 99176 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _468_
timestamp 1
transform -1 0 100372 0 1 73984
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_2  _469_
timestamp 1
transform 1 0 97980 0 -1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _470_
timestamp 1
transform -1 0 101384 0 1 76160
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _471_
timestamp 1
transform 1 0 99912 0 1 76160
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1
transform -1 0 99636 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _473_
timestamp 1
transform -1 0 99912 0 1 76160
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _474_
timestamp 1
transform -1 0 99268 0 1 76160
box -38 -48 1602 592
use sky130_fd_sc_hd__a311o_1  _475_
timestamp 1
transform 1 0 99084 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _476_
timestamp 1
transform -1 0 99820 0 1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _477_
timestamp 1
transform 1 0 100372 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _478_
timestamp 1
transform 1 0 99084 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _479_
timestamp 1
transform -1 0 97244 0 1 73984
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _480_
timestamp 1
transform 1 0 96416 0 -1 75072
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 1
transform -1 0 97888 0 1 75072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _482_
timestamp 1
transform 1 0 98624 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _483_
timestamp 1
transform -1 0 98440 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _484_
timestamp 1
transform -1 0 98348 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _485_
timestamp 1
transform -1 0 98992 0 -1 76160
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _486_
timestamp 1
transform 1 0 98072 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _487_
timestamp 1
transform 1 0 97060 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _488_
timestamp 1
transform -1 0 95956 0 1 72896
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _489_
timestamp 1
transform -1 0 97428 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _490_
timestamp 1
transform -1 0 96048 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _491_
timestamp 1
transform -1 0 97520 0 1 68544
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _492_
timestamp 1
transform 1 0 96140 0 -1 68544
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _493_
timestamp 1
transform -1 0 97152 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _494_
timestamp 1
transform 1 0 94576 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _495_
timestamp 1
transform 1 0 96600 0 -1 68544
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _496_
timestamp 1
transform 1 0 95220 0 -1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _497_
timestamp 1
transform -1 0 96048 0 1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _498_
timestamp 1
transform 1 0 93932 0 -1 66368
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _499_
timestamp 1
transform -1 0 96048 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _500_
timestamp 1
transform -1 0 96140 0 1 68544
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _501_
timestamp 1
transform -1 0 96048 0 -1 67456
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _502_
timestamp 1
transform -1 0 96416 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _503_
timestamp 1
transform 1 0 94576 0 1 68544
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _504_
timestamp 1
transform 1 0 97428 0 1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _505_
timestamp 1
transform -1 0 96232 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _506_
timestamp 1
transform -1 0 94668 0 -1 75072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _507_
timestamp 1
transform -1 0 93748 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _508_
timestamp 1
transform 1 0 93932 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _509_
timestamp 1
transform 1 0 93380 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _510_
timestamp 1
transform -1 0 95404 0 1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _511_
timestamp 1
transform 1 0 94944 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _512_
timestamp 1
transform 1 0 94024 0 1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _513_
timestamp 1
transform -1 0 97060 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _514_
timestamp 1
transform 1 0 97060 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _515_
timestamp 1
transform -1 0 96324 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _516_
timestamp 1
transform -1 0 95404 0 1 67456
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _517_
timestamp 1
transform -1 0 88044 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _518_
timestamp 1
transform 1 0 89516 0 1 77248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _519_
timestamp 1
transform -1 0 90620 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _520_
timestamp 1
transform -1 0 90344 0 -1 76160
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _521_
timestamp 1
transform -1 0 92184 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _522_
timestamp 1
transform 1 0 91264 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _523_
timestamp 1
transform -1 0 91080 0 -1 73984
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _524_
timestamp 1
transform -1 0 94208 0 1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _525_
timestamp 1
transform -1 0 92644 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _526_
timestamp 1
transform 1 0 92920 0 1 70720
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _527_
timestamp 1
transform -1 0 92368 0 -1 69632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _528_
timestamp 1
transform -1 0 93656 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _529_
timestamp 1
transform -1 0 93380 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _530_
timestamp 1
transform -1 0 92000 0 -1 68544
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _531_
timestamp 1
transform -1 0 92828 0 1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _532_
timestamp 1
transform -1 0 90528 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _533_
timestamp 1
transform 1 0 91632 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _534_
timestamp 1
transform -1 0 90068 0 1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _535_
timestamp 1
transform -1 0 91448 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _536_
timestamp 1
transform -1 0 90988 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _537_
timestamp 1
transform -1 0 90712 0 -1 66368
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _538_
timestamp 1
transform -1 0 89976 0 1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _539_
timestamp 1
transform -1 0 89608 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _540_
timestamp 1
transform -1 0 89976 0 -1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _541_
timestamp 1
transform -1 0 89516 0 1 67456
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _542_
timestamp 1
transform -1 0 89424 0 -1 69632
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _543_
timestamp 1
transform -1 0 88412 0 -1 70720
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _544_
timestamp 1
transform 1 0 26680 0 1 76160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _545_
timestamp 1
transform 1 0 23184 0 1 76160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _546_
timestamp 1
transform 1 0 28520 0 1 76160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _547_
timestamp 1
transform 1 0 35052 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _548_
timestamp 1
transform 1 0 25392 0 -1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _549_
timestamp 1
transform 1 0 37352 0 1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _550_
timestamp 1
transform 1 0 39836 0 1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _551_
timestamp 1
transform -1 0 69000 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _552_
timestamp 1
transform -1 0 70656 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _553_
timestamp 1
transform -1 0 73140 0 1 72896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _554_
timestamp 1
transform -1 0 74980 0 -1 73984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _555_
timestamp 1
transform -1 0 84456 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _556_
timestamp 1
transform -1 0 83536 0 1 76160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _557_
timestamp 1
transform -1 0 91816 0 -1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _558_
timestamp 1
transform -1 0 87124 0 1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _559_
timestamp 1
transform -1 0 89608 0 -1 77248
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _560_
timestamp 1
transform -1 0 22448 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _561_
timestamp 1
transform -1 0 25668 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _562_
timestamp 1
transform -1 0 28060 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _563_
timestamp 1
transform -1 0 22540 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _564_
timestamp 1
transform -1 0 28336 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _565_
timestamp 1
transform -1 0 29808 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _566_
timestamp 1
transform -1 0 85008 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _567_
timestamp 1
transform 1 0 85376 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _568_
timestamp 1
transform 1 0 87768 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp 1
transform 1 0 87124 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _570_
timestamp 1
transform 1 0 90712 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _571_
timestamp 1
transform 1 0 91448 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _572_
timestamp 1
transform 1 0 94852 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _573_
timestamp 1
transform 1 0 93932 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _574_
timestamp 1
transform 1 0 94024 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1
transform 1 0 85560 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _576_
timestamp 1
transform 1 0 89516 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1
transform 1 0 88412 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _578_
timestamp 1
transform 1 0 89792 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _579_
timestamp 1
transform 1 0 89424 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _580_
timestamp 1
transform 1 0 86664 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _581_
timestamp 1
transform 1 0 86664 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _582_
timestamp 1
transform 1 0 84916 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _583_
timestamp 1
transform 1 0 85376 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _584_
timestamp 1
transform -1 0 19044 0 -1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _585_
timestamp 1
transform -1 0 16560 0 -1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _586_
timestamp 1
transform -1 0 19964 0 -1 75072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _587_
timestamp 1
transform -1 0 23276 0 1 72896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _588_
timestamp 1
transform -1 0 16560 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _589_
timestamp 1
transform -1 0 23644 0 1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _590_
timestamp 1
transform -1 0 25116 0 -1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _591_
timestamp 1
transform 1 0 85652 0 -1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _592_
timestamp 1
transform 1 0 86388 0 -1 72896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _593_
timestamp 1
transform 1 0 88780 0 -1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _594_
timestamp 1
transform 1 0 88320 0 1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _595_
timestamp 1
transform 1 0 92736 0 1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _596_
timestamp 1
transform 1 0 93104 0 1 75072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _597_
timestamp 1
transform 1 0 97152 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _598_
timestamp 1
transform 1 0 95128 0 -1 76160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _599_
timestamp 1
transform 1 0 95772 0 -1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _600_
timestamp 1
transform -1 0 88136 0 -1 75072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _601_
timestamp 1
transform 1 0 88688 0 1 75072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _602_
timestamp 1
transform 1 0 89332 0 -1 71808
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _603_
timestamp 1
transform 1 0 91356 0 1 68544
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _604_
timestamp 1
transform -1 0 91908 0 -1 69632
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _605_
timestamp 1
transform -1 0 89332 0 1 66368
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _606_
timestamp 1
transform -1 0 89056 0 1 67456
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _607_
timestamp 1
transform -1 0 88320 0 -1 66368
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _608_
timestamp 1
transform -1 0 88136 0 1 70720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _609_
timestamp 1
transform -1 0 33580 0 -1 70720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _610_
timestamp 1
transform -1 0 32016 0 -1 70720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _611_
timestamp 1
transform -1 0 35972 0 -1 70720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _612_
timestamp 1
transform -1 0 40296 0 -1 68544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _613_
timestamp 1
transform -1 0 37168 0 1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _614_
timestamp 1
transform -1 0 43884 0 -1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _615_
timestamp 1
transform -1 0 46460 0 1 68544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _616_
timestamp 1
transform 1 0 58880 0 1 68544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _617_
timestamp 1
transform 1 0 61456 0 -1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _618_
timestamp 1
transform 1 0 65596 0 1 68544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _619_
timestamp 1
transform 1 0 66608 0 -1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _620_
timestamp 1
transform 1 0 72864 0 1 70720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _621_
timestamp 1
transform 1 0 73692 0 1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _622_
timestamp 1
transform 1 0 79396 0 1 70720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _623_
timestamp 1
transform 1 0 77556 0 1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _624_
timestamp 1
transform 1 0 79488 0 1 69632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _625_
timestamp 1
transform 1 0 6164 0 1 93568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _626_
timestamp 1
transform 1 0 6164 0 1 100096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _627_
timestamp 1
transform 1 0 24380 0 1 77248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _628_
timestamp 1
transform -1 0 41308 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _629_
timestamp 1
transform 1 0 6164 0 1 117504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _630_
timestamp 1
transform -1 0 44344 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _631_
timestamp 1
transform -1 0 46920 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _632_
timestamp 1
transform 1 0 60720 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _633_
timestamp 1
transform 1 0 62836 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _634_
timestamp 1
transform 1 0 65596 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _635_
timestamp 1
transform 1 0 67620 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _636_
timestamp 1
transform -1 0 85376 0 -1 137088
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _637_
timestamp 1
transform -1 0 85192 0 1 76160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _638_
timestamp 1
transform 1 0 104328 0 1 113152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _639_
timestamp 1
transform 1 0 104328 0 -1 101184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _640_
timestamp 1
transform 1 0 104328 0 -1 96832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _641_
timestamp 1
transform -1 0 80224 0 1 72896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _642_
timestamp 1
transform -1 0 83444 0 1 71808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform -1 0 21804 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 66424 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform -1 0 66792 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 72864 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform -1 0 73692 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform -1 0 77556 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform -1 0 79488 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform 1 0 79488 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform -1 0 30728 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform -1 0 42596 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform -1 0 46644 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform -1 0 58880 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform 1 0 61272 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform 1 0 61456 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform -1 0 67252 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform 1 0 86204 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform -1 0 1932 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform 1 0 83536 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1
transform 1 0 24656 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1
transform 1 0 94392 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__A
timestamp 1
transform 1 0 95036 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__A
timestamp 1
transform 1 0 93656 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__B1
timestamp 1
transform -1 0 96232 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__A
timestamp 1
transform 1 0 95220 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__A
timestamp 1
transform 1 0 94392 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__A
timestamp 1
transform 1 0 93288 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__A1
timestamp 1
transform 1 0 93748 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__A
timestamp 1
transform 1 0 94576 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__A_N
timestamp 1
transform 1 0 88044 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__A
timestamp 1
transform -1 0 89516 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__A
timestamp 1
transform 1 0 90160 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__A
timestamp 1
transform 1 0 92184 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__C
timestamp 1
transform 1 0 92368 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A1
timestamp 1
transform 1 0 90896 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__B1
timestamp 1
transform -1 0 91264 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1
transform 1 0 93012 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__C
timestamp 1
transform 1 0 94208 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__D
timestamp 1
transform 1 0 93196 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A1
timestamp 1
transform 1 0 92552 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A3
timestamp 1
transform 1 0 92736 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__B1
timestamp 1
transform 1 0 94392 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__A
timestamp 1
transform 1 0 93656 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__A
timestamp 1
transform 1 0 92736 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__531__A
timestamp 1
transform 1 0 92184 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__531__B
timestamp 1
transform 1 0 92000 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__A1
timestamp 1
transform 1 0 92184 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__B1
timestamp 1
transform 1 0 91356 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__A
timestamp 1
transform 1 0 90804 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__536__A
timestamp 1
transform 1 0 90988 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__A
timestamp 1
transform 1 0 90068 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A
timestamp 1
transform 1 0 89148 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__A
timestamp 1
transform 1 0 89332 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A1
timestamp 1
transform 1 0 26496 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__S
timestamp 1
transform 1 0 27508 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__A1
timestamp 1
transform 1 0 23000 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__S
timestamp 1
transform 1 0 24012 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__S
timestamp 1
transform 1 0 29532 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__S
timestamp 1
transform 1 0 35880 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A1
timestamp 1
transform -1 0 25392 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__S
timestamp 1
transform -1 0 26404 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__S
timestamp 1
transform -1 0 38364 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__S
timestamp 1
transform -1 0 40848 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__S
timestamp 1
transform 1 0 69000 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__S
timestamp 1
transform 1 0 70656 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__553__S
timestamp 1
transform -1 0 73324 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__S
timestamp 1
transform 1 0 74980 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A1
timestamp 1
transform 1 0 84456 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__S
timestamp 1
transform 1 0 83352 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__S
timestamp 1
transform 1 0 82524 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A1
timestamp 1
transform -1 0 92184 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__S
timestamp 1
transform 1 0 90804 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A1
timestamp 1
transform 1 0 87124 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__S
timestamp 1
transform 1 0 85928 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__A1
timestamp 1
transform -1 0 89792 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__S
timestamp 1
transform 1 0 88504 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1
transform 1 0 22448 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A
timestamp 1
transform 1 0 25668 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A
timestamp 1
transform 1 0 28060 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__563__A
timestamp 1
transform 1 0 22540 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1
transform 1 0 28336 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1
transform 1 0 29808 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1
transform 1 0 85008 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A
timestamp 1
transform 1 0 85652 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A
timestamp 1
transform 1 0 88044 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__A
timestamp 1
transform 1 0 87400 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__A
timestamp 1
transform 1 0 90988 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__A
timestamp 1
transform 1 0 91724 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1
transform -1 0 95312 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1
transform 1 0 94208 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1
transform -1 0 94484 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A
timestamp 1
transform 1 0 85836 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__A
timestamp 1
transform 1 0 89792 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__A
timestamp 1
transform 1 0 88688 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A
timestamp 1
transform 1 0 90068 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__A
timestamp 1
transform 1 0 89700 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__A
timestamp 1
transform -1 0 87124 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__581__A
timestamp 1
transform 1 0 86940 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__A
timestamp 1
transform 1 0 85192 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A
timestamp 1
transform 1 0 85652 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__CLK
timestamp 1
transform 1 0 17020 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__585__CLK
timestamp 1
transform 1 0 14536 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__CLK
timestamp 1
transform 1 0 17940 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__587__CLK
timestamp 1
transform 1 0 23460 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__587__Q
timestamp 1
transform -1 0 23460 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__CLK
timestamp 1
transform -1 0 14720 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__CLK
timestamp 1
transform -1 0 24012 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__Q
timestamp 1
transform -1 0 23828 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__CLK
timestamp 1
transform 1 0 25300 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__Q
timestamp 1
transform -1 0 25300 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__CLK
timestamp 1
transform 1 0 85468 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__Q
timestamp 1
transform -1 0 87676 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__592__CLK
timestamp 1
transform 1 0 86020 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__592__Q
timestamp 1
transform -1 0 88412 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__CLK
timestamp 1
transform 1 0 91264 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__Q
timestamp 1
transform -1 0 91264 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__594__CLK
timestamp 1
transform 1 0 90344 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__594__Q
timestamp 1
transform 1 0 90160 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__595__CLK
timestamp 1
transform 1 0 92552 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__596__CLK
timestamp 1
transform 1 0 92920 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__597__CLK
timestamp 1
transform 1 0 99084 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__CLK
timestamp 1
transform 1 0 94944 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__CLK
timestamp 1
transform -1 0 97796 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__CLK
timestamp 1
transform 1 0 88320 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__Q
timestamp 1
transform -1 0 88320 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__CLK
timestamp 1
transform 1 0 90804 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__CLK
timestamp 1
transform 1 0 89148 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__Q
timestamp 1
transform 1 0 91448 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__CLK
timestamp 1
transform 1 0 91080 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__Q
timestamp 1
transform 1 0 93472 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__CLK
timestamp 1
transform -1 0 93012 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__Q
timestamp 1
transform 1 0 92644 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__CLK
timestamp 1
transform 1 0 87032 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__Q
timestamp 1
transform 1 0 90068 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__CLK
timestamp 1
transform 1 0 86756 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__Q
timestamp 1
transform 1 0 89056 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__CLK
timestamp 1
transform 1 0 85928 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__Q
timestamp 1
transform 1 0 88504 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__608__CLK
timestamp 1
transform 1 0 85928 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__CLK
timestamp 1
transform 1 0 32200 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__CLK
timestamp 1
transform 1 0 32016 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__CLK
timestamp 1
transform 1 0 34316 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__CLK
timestamp 1
transform -1 0 38824 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__CLK
timestamp 1
transform 1 0 35512 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__614__CLK
timestamp 1
transform 1 0 42136 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__615__CLK
timestamp 1
transform 1 0 44712 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__CLK
timestamp 1
transform 1 0 58512 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__617__CLK
timestamp 1
transform 1 0 63020 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__CLK
timestamp 1
transform 1 0 67252 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__CLK
timestamp 1
transform 1 0 68172 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__CLK
timestamp 1
transform 1 0 72496 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__CLK
timestamp 1
transform 1 0 73324 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__CLK
timestamp 1
transform 1 0 81052 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__D
timestamp 1
transform -1 0 79396 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__CLK
timestamp 1
transform 1 0 79028 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__CLK
timestamp 1
transform 1 0 81052 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__CLK
timestamp 1
transform 1 0 7452 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__D
timestamp 1
transform -1 0 7452 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__Q
timestamp 1
transform -1 0 7268 0 -1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__CLK
timestamp 1
transform 1 0 7452 0 -1 100096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__D
timestamp 1
transform 1 0 7452 0 -1 101184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__Q
timestamp 1
transform -1 0 7452 0 -1 100096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__CLK
timestamp 1
transform -1 0 24288 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__D
timestamp 1
transform 1 0 25852 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__CLK
timestamp 1
transform 1 0 41492 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__D
timestamp 1
transform 1 0 41308 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__CLK
timestamp 1
transform 1 0 7452 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__D
timestamp 1
transform 1 0 7452 0 -1 118592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__Q
timestamp 1
transform -1 0 7452 0 -1 117504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__CLK
timestamp 1
transform 1 0 44528 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__D
timestamp 1
transform 1 0 44344 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__CLK
timestamp 1
transform 1 0 47104 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__D
timestamp 1
transform 1 0 46920 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__632__CLK
timestamp 1
transform 1 0 60444 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__632__D
timestamp 1
transform 1 0 60168 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__CLK
timestamp 1
transform -1 0 64492 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__D
timestamp 1
transform 1 0 62652 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__634__CLK
timestamp 1
transform -1 0 67252 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__634__D
timestamp 1
transform 1 0 65320 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__CLK
timestamp 1
transform -1 0 69276 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__D
timestamp 1
transform 1 0 67436 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__CLK
timestamp 1
transform 1 0 85560 0 -1 137088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__D
timestamp 1
transform 1 0 83628 0 -1 137088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__Q
timestamp 1
transform -1 0 85560 0 -1 137088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__637__CLK
timestamp 1
transform 1 0 85192 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__637__D
timestamp 1
transform -1 0 83812 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__CLK
timestamp 1
transform 1 0 105984 0 1 113152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__D
timestamp 1
transform -1 0 104512 0 -1 113152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__Q
timestamp 1
transform -1 0 105984 0 1 113152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__CLK
timestamp 1
transform 1 0 105984 0 -1 101184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__D
timestamp 1
transform -1 0 104512 0 1 100096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__Q
timestamp 1
transform -1 0 105984 0 -1 101184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__CLK
timestamp 1
transform 1 0 105984 0 -1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__D
timestamp 1
transform -1 0 104512 0 1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__Q
timestamp 1
transform -1 0 105984 0 -1 96832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__CLK
timestamp 1
transform 1 0 78568 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__CLK
timestamp 1
transform 1 0 83444 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1
transform 1 0 55108 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 1
transform 1 0 57132 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_A
timestamp 1
transform -1 0 73232 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_X
timestamp 1
transform -1 0 74520 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_A
timestamp 1
transform -1 0 104512 0 -1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_X
timestamp 1
transform 1 0 105340 0 1 91392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_A
timestamp 1
transform 1 0 5060 0 -1 82688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_X
timestamp 1
transform 1 0 5244 0 -1 82688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_A
timestamp 1
transform 1 0 48300 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_X
timestamp 1
transform 1 0 48484 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_clk_A
timestamp 1
transform -1 0 70380 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_clk_X
timestamp 1
transform 1 0 70380 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_clk_A
timestamp 1
transform 1 0 82800 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_clk_X
timestamp 1
transform 1 0 84824 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_clk_A
timestamp 1
transform 1 0 94484 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_clk_X
timestamp 1
transform -1 0 94852 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_clk_A
timestamp 1
transform -1 0 106352 0 1 106624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_clk_X
timestamp 1
transform -1 0 106536 0 1 106624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_clk_A
timestamp 1
transform -1 0 11408 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_clk_X
timestamp 1
transform 1 0 13432 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_clk_A
timestamp 1
transform -1 0 5796 0 1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_clk_X
timestamp 1
transform 1 0 7452 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_clk_A
timestamp 1
transform 1 0 32936 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_clk_X
timestamp 1
transform 1 0 33120 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_clk_A
timestamp 1
transform -1 0 55200 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_clk_X
timestamp 1
transform -1 0 57316 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 1
transform 1 0 69000 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload1_A
timestamp 1
transform 1 0 93104 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload2_A
timestamp 1
transform 1 0 6440 0 -1 94656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload3_A
timestamp 1
transform 1 0 55016 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout100_X
timestamp 1
transform -1 0 74060 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout101_X
timestamp 1
transform 1 0 74980 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_A
timestamp 1
transform 1 0 87860 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_X
timestamp 1
transform 1 0 88780 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1
transform 1 0 90988 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_X
timestamp 1
transform 1 0 91540 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1
transform -1 0 91540 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_X
timestamp 1
transform 1 0 89516 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1
transform 1 0 90988 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_X
timestamp 1
transform 1 0 91172 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1
transform -1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_X
timestamp 1
transform -1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1
transform -1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_X
timestamp 1
transform 1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1
transform -1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_X
timestamp 1
transform -1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1
transform -1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_X
timestamp 1
transform -1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1
transform -1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_X
timestamp 1
transform -1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1
transform -1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_X
timestamp 1
transform 1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1
transform -1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_X
timestamp 1
transform 1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1
transform -1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_X
timestamp 1
transform -1 0 1932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1
transform -1 0 2116 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_X
timestamp 1
transform -1 0 1932 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1
transform -1 0 1564 0 -1 80512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_X
timestamp 1
transform -1 0 2484 0 1 80512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1
transform -1 0 1840 0 -1 104448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1
transform -1 0 1840 0 1 105536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1
transform -1 0 1840 0 1 106624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1
transform -1 0 1840 0 -1 108800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1
transform -1 0 1840 0 -1 109888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1
transform -1 0 1840 0 1 110976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1
transform -1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_X
timestamp 1
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1
transform -1 0 1840 0 1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1
transform -1 0 108284 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1
transform -1 0 108284 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1
transform -1 0 108560 0 -1 80512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1
transform -1 0 108284 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1
transform -1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_X
timestamp 1
transform -1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1
transform -1 0 37444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1
transform -1 0 38732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1
transform -1 0 40020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1
transform -1 0 41308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1
transform -1 0 43240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1
transform -1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_X
timestamp 1
transform 1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1
transform -1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_X
timestamp 1
transform -1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1
transform -1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_X
timestamp 1
transform -1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1
transform -1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_X
timestamp 1
transform 1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1
transform -1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1
transform -1 0 35512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1
transform -1 0 36156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1
transform -1 0 2116 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_X
timestamp 1
transform 1 0 1748 0 -1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1
transform -1 0 2116 0 1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_X
timestamp 1
transform 1 0 1748 0 1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1
transform -1 0 2116 0 1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_X
timestamp 1
transform -1 0 1932 0 1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1
transform -1 0 2116 0 -1 82688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_X
timestamp 1
transform 1 0 1748 0 -1 82688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1
transform -1 0 2116 0 -1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_X
timestamp 1
transform 1 0 1748 0 -1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1
transform -1 0 2116 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_X
timestamp 1
transform 1 0 1748 0 -1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1
transform -1 0 2116 0 1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_X
timestamp 1
transform -1 0 1932 0 1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1
transform -1 0 2116 0 -1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_X
timestamp 1
transform 1 0 1748 0 -1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1
transform -1 0 2116 0 1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_X
timestamp 1
transform -1 0 1932 0 1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1
transform -1 0 2116 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_X
timestamp 1
transform 1 0 1748 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1
transform -1 0 2116 0 -1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_X
timestamp 1
transform 1 0 1748 0 -1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1
transform -1 0 2116 0 1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_X
timestamp 1
transform -1 0 1932 0 1 87040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1
transform -1 0 2116 0 -1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_X
timestamp 1
transform 1 0 1748 0 -1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1
transform -1 0 2116 0 -1 88128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_X
timestamp 1
transform 1 0 1748 0 -1 88128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1
transform -1 0 2116 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_X
timestamp 1
transform -1 0 1932 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1
transform -1 0 2116 0 -1 89216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_X
timestamp 1
transform 1 0 1748 0 -1 89216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1
transform -1 0 108284 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1
transform -1 0 108284 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1
transform -1 0 108284 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1
transform -1 0 108284 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1
transform -1 0 108284 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_X
timestamp 1
transform 1 0 107916 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[0]
timestamp 1
transform -1 0 23644 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[1]
timestamp 1
transform -1 0 24840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[2]
timestamp 1
transform -1 0 7636 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[3]
timestamp 1
transform -1 0 7636 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[4]
timestamp 1
transform -1 0 7636 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[5]
timestamp 1
transform -1 0 7636 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[6]
timestamp 1
transform -1 0 7636 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr0[7]
timestamp 1
transform -1 0 7636 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[0]
timestamp 1
transform 1 0 88320 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[2]
timestamp 1
transform -1 0 104512 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[3]
timestamp 1
transform -1 0 104512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[4]
timestamp 1
transform -1 0 104512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[5]
timestamp 1
transform -1 0 90712 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[6]
timestamp 1
transform -1 0 90896 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_addr1[7]
timestamp 1
transform -1 0 91080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_clk0
timestamp 1
transform -1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_clk1
timestamp 1
transform -1 0 96416 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_csb0
timestamp 1
transform -1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[0]
timestamp 1
transform -1 0 26036 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[1]
timestamp 1
transform -1 0 27140 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[2]
timestamp 1
transform -1 0 28336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[3]
timestamp 1
transform -1 0 29716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_din0[4]
timestamp 1
transform -1 0 30636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i0_dout1[13]
timestamp 1
transform 1 0 68540 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr0[0]
timestamp 1
transform -1 0 23644 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr0[1]
timestamp 1
transform -1 0 24840 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[0]
timestamp 1
transform -1 0 87492 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[1]
timestamp 1
transform -1 0 86388 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[2]
timestamp 1
transform -1 0 104512 0 -1 95744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[3]
timestamp 1
transform -1 0 104512 0 1 93568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[4]
timestamp 1
transform -1 0 104512 0 1 92480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[5]
timestamp 1
transform 1 0 91356 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[6]
timestamp 1
transform 1 0 91540 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_addr1[7]
timestamp 1
transform 1 0 91724 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_clk0
timestamp 1
transform -1 0 16836 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_clk1
timestamp 1
transform 1 0 95864 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[0]
timestamp 1
transform -1 0 26220 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[1]
timestamp 1
transform -1 0 27140 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[2]
timestamp 1
transform -1 0 28336 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[3]
timestamp 1
transform -1 0 29716 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[4]
timestamp 1
transform -1 0 30636 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[5]
timestamp 1
transform -1 0 31832 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[6]
timestamp 1
transform -1 0 33028 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[7]
timestamp 1
transform -1 0 34132 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[8]
timestamp 1
transform -1 0 35328 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[9]
timestamp 1
transform -1 0 36524 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[10]
timestamp 1
transform -1 0 37628 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[11]
timestamp 1
transform -1 0 38824 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[12]
timestamp 1
transform -1 0 40020 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[13]
timestamp 1
transform -1 0 41216 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[14]
timestamp 1
transform -1 0 42320 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_din0[15]
timestamp 1
transform -1 0 43516 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_dout1[4]
timestamp 1
transform -1 0 46276 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_dout1[11]
timestamp 1
transform 1 0 63572 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i1_dout1[13]
timestamp 1
transform -1 0 68724 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1
transform -1 0 108192 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output69_A
timestamp 1
transform 1 0 1748 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1
transform -1 0 1932 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1
transform 1 0 1748 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1
transform -1 0 108192 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1
transform -1 0 108192 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1
transform 1 0 108008 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_rebuffer3_X
timestamp 1
transform -1 0 92000 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire87_X
timestamp 1
transform -1 0 60996 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire88_X
timestamp 1
transform -1 0 58420 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire89_X
timestamp 1
transform -1 0 55844 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire90_X
timestamp 1
transform -1 0 50692 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire91_X
timestamp 1
transform -1 0 48116 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire92_X
timestamp 1
transform -1 0 43516 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire93_X
timestamp 1
transform -1 0 36524 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire94_X
timestamp 1
transform -1 0 35512 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire95_X
timestamp 1
transform -1 0 77832 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire96_X
timestamp 1
transform -1 0 73876 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire97_X
timestamp 1
transform -1 0 72956 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire98_X
timestamp 1
transform -1 0 63572 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wire99_X
timestamp 1
transform -1 0 34868 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform 1 0 55292 0 -1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_2_0_0_clk
timestamp 1
transform 1 0 73324 0 -1 66368
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_2_1_0_clk
timestamp 1
transform 1 0 104328 0 1 91392
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_2_2_0_clk
timestamp 1
transform -1 0 5060 0 -1 82688
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_2_3_0_clk
timestamp 1
transform 1 0 47288 0 1 70720
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1
transform -1 0 70196 0 1 72896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1
transform 1 0 82984 0 1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1
transform -1 0 93840 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1
transform 1 0 104328 0 1 106624
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1
transform 1 0 11592 0 -1 73984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1
transform 1 0 5796 0 1 94656
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1
transform -1 0 32936 0 1 70720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1
transform 1 0 55292 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_6  clkload0
timestamp 1
transform 1 0 68356 0 -1 72896
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp 1
transform 1 0 92552 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp 1
transform 1 0 6624 0 -1 94656
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinvlp_4  clkload3
timestamp 1
transform 1 0 54464 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 1
transform -1 0 98348 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout100
timestamp 1
transform -1 0 73876 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout101
timestamp 1
transform -1 0 74980 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout102
timestamp 1
transform 1 0 88044 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout103
timestamp 1
transform 1 0 90436 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout104
timestamp 1
transform -1 0 90436 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout105
timestamp 1
transform -1 0 90988 0 -1 70720
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp 1
transform -1 0 103316 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout107
timestamp 1
transform -1 0 102764 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  fanout108
timestamp 1
transform -1 0 104604 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 1
transform 1 0 103776 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout110
timestamp 1
transform -1 0 104328 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp 1
transform -1 0 105708 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout112
timestamp 1
transform -1 0 106076 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 1
transform 1 0 105616 0 -1 71808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636968456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_321
timestamp 1
transform 1 0 30636 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_329
timestamp 1
transform 1 0 31372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_343
timestamp 1
transform 1 0 32660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 1
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_357
timestamp 1
transform 1 0 33948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_365
timestamp 1
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_371
timestamp 1
transform 1 0 35236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_377
timestamp 1
transform 1 0 35788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_398
timestamp 1
transform 1 0 37720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_406
timestamp 1
transform 1 0 38456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_426
timestamp 1
transform 1 0 40296 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_434
timestamp 1
transform 1 0 41032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_440
timestamp 1
transform 1 0 41584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_449
timestamp 1
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_455
timestamp 1
transform 1 0 42964 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1636968456
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636968456
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636968456
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636968456
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1636968456
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1636968456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1636968456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1636968456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1636968456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1636968456
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1636968456
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1636968456
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1636968456
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1636968456
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1636968456
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1636968456
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1636968456
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1636968456
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1636968456
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1636968456
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1636968456
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1636968456
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1636968456
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1636968456
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1636968456
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1636968456
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1636968456
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1636968456
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1636968456
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1636968456
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1636968456
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1636968456
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1636968456
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1636968456
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1636968456
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1636968456
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1636968456
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1636968456
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1636968456
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1636968456
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1636968456
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1636968456
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1636968456
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1636968456
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1636968456
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1636968456
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1636968456
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1636968456
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1636968456
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1636968456
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1161
timestamp 1
transform 1 0 107916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1167
timestamp 1
transform 1 0 108468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636968456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636968456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636968456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636968456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636968456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636968456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636968456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636968456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636968456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636968456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636968456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636968456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636968456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636968456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636968456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636968456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636968456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636968456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636968456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636968456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636968456
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636968456
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636968456
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636968456
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636968456
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636968456
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636968456
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636968456
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636968456
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636968456
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636968456
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636968456
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636968456
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636968456
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636968456
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636968456
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636968456
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636968456
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636968456
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636968456
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1636968456
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1636968456
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1636968456
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1636968456
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1636968456
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1636968456
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1636968456
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1636968456
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1636968456
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1636968456
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1636968456
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1636968456
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1636968456
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1636968456
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1636968456
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1636968456
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1636968456
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1636968456
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1636968456
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1157
timestamp 1
transform 1 0 107548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1165
timestamp 1
transform 1 0 108284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636968456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636968456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636968456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636968456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636968456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636968456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636968456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636968456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636968456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636968456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636968456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636968456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636968456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636968456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636968456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636968456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636968456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636968456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636968456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636968456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636968456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636968456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636968456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636968456
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636968456
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636968456
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636968456
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636968456
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636968456
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636968456
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636968456
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636968456
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636968456
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636968456
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636968456
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636968456
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636968456
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636968456
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636968456
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636968456
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636968456
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636968456
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636968456
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1636968456
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1636968456
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1636968456
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1636968456
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1636968456
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1636968456
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1636968456
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1636968456
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1636968456
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1636968456
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1636968456
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1636968456
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1636968456
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1636968456
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1636968456
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1636968456
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1636968456
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1636968456
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1161
timestamp 1
transform 1 0 107916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1167
timestamp 1
transform 1 0 108468 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636968456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636968456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636968456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636968456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636968456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636968456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636968456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636968456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636968456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636968456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636968456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636968456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636968456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636968456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636968456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636968456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636968456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636968456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636968456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636968456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636968456
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636968456
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636968456
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636968456
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636968456
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636968456
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636968456
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636968456
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636968456
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636968456
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636968456
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636968456
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636968456
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636968456
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636968456
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636968456
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636968456
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636968456
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636968456
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636968456
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1636968456
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1636968456
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1636968456
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1636968456
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1636968456
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1636968456
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1636968456
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1636968456
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1636968456
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1636968456
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1636968456
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1636968456
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1636968456
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1636968456
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1636968456
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1636968456
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1636968456
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1636968456
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1636968456
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1157
timestamp 1
transform 1 0 107548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1165
timestamp 1
transform 1 0 108284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636968456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636968456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636968456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636968456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636968456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636968456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636968456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636968456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636968456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636968456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636968456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636968456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636968456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636968456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636968456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636968456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636968456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636968456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636968456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636968456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636968456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636968456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636968456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636968456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636968456
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636968456
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636968456
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636968456
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636968456
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636968456
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636968456
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636968456
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636968456
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636968456
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636968456
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636968456
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636968456
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636968456
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636968456
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1636968456
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1636968456
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636968456
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636968456
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1636968456
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1636968456
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1636968456
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1636968456
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1636968456
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1636968456
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1636968456
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1636968456
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1636968456
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1636968456
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1636968456
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1636968456
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1636968456
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1636968456
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1636968456
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1636968456
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1636968456
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1636968456
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1636968456
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1161
timestamp 1
transform 1 0 107916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1167
timestamp 1
transform 1 0 108468 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1636968456
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1636968456
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1636968456
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636968456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636968456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636968456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636968456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636968456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636968456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636968456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636968456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636968456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636968456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636968456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636968456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636968456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636968456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636968456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636968456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636968456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636968456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636968456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636968456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636968456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636968456
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636968456
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636968456
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636968456
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636968456
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636968456
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636968456
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636968456
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636968456
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636968456
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636968456
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636968456
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636968456
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636968456
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1636968456
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1636968456
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1636968456
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1636968456
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1636968456
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636968456
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1636968456
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1636968456
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1636968456
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1636968456
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1636968456
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1636968456
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1636968456
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1636968456
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1636968456
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1636968456
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1636968456
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1636968456
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1636968456
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1636968456
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1636968456
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1636968456
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1636968456
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1636968456
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1636968456
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1157
timestamp 1
transform 1 0 107548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1165
timestamp 1
transform 1 0 108284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_10
timestamp 1636968456
transform 1 0 2024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636968456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636968456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636968456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636968456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636968456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636968456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636968456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636968456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636968456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636968456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636968456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636968456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636968456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636968456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636968456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1636968456
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1636968456
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636968456
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636968456
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1636968456
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1636968456
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636968456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636968456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1636968456
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1636968456
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636968456
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636968456
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1636968456
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1636968456
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636968456
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636968456
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1636968456
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1636968456
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636968456
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636968456
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1636968456
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1636968456
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1636968456
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1636968456
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1636968456
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1636968456
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1636968456
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1636968456
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1636968456
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1636968456
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1636968456
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1636968456
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1636968456
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1636968456
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1636968456
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1636968456
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1636968456
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1636968456
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1636968456
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1636968456
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1636968456
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1636968456
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1636968456
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1636968456
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1636968456
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1636968456
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1636968456
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1161
timestamp 1
transform 1 0 107916 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1167
timestamp 1
transform 1 0 108468 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_11
timestamp 1636968456
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1636968456
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1636968456
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636968456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636968456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636968456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636968456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636968456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636968456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636968456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636968456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636968456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636968456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636968456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636968456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636968456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636968456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636968456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636968456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1636968456
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1636968456
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1636968456
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636968456
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636968456
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636968456
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636968456
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1636968456
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1636968456
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1636968456
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1636968456
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1636968456
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1636968456
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1636968456
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1636968456
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1636968456
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1636968456
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1636968456
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1636968456
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1636968456
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1636968456
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1636968456
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1636968456
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1636968456
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1636968456
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1636968456
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1636968456
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1636968456
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1636968456
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1636968456
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1636968456
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1636968456
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1636968456
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1636968456
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1636968456
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1636968456
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1636968456
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1636968456
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1636968456
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1636968456
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1636968456
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1636968456
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1636968456
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1636968456
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1636968456
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1636968456
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1636968456
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1636968456
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1636968456
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1636968456
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1157
timestamp 1
transform 1 0 107548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_1165
timestamp 1
transform 1 0 108284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636968456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636968456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636968456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636968456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636968456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636968456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636968456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636968456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636968456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636968456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636968456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636968456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636968456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636968456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636968456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636968456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636968456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636968456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636968456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636968456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636968456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636968456
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636968456
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636968456
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636968456
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636968456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636968456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1636968456
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1636968456
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1636968456
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1636968456
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1636968456
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1636968456
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1636968456
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1636968456
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1636968456
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1636968456
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1636968456
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1636968456
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1636968456
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1636968456
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1636968456
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1636968456
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1636968456
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1636968456
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1636968456
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1636968456
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1636968456
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1636968456
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1636968456
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1636968456
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1636968456
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1636968456
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1636968456
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1636968456
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1636968456
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1636968456
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1636968456
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1636968456
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1636968456
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1636968456
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1636968456
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1636968456
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1636968456
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1636968456
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1636968456
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1636968456
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1636968456
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1636968456
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1636968456
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1161
timestamp 1
transform 1 0 107916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1167
timestamp 1
transform 1 0 108468 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_11
timestamp 1636968456
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1636968456
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1636968456
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1636968456
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1636968456
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1636968456
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_153
timestamp 1
transform 1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636968456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1636968456
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1636968456
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1
transform 1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_245
timestamp 1
transform 1 0 23644 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_251
timestamp 1
transform 1 0 24196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_253
timestamp 1
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_258
timestamp 1
transform 1 0 24840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_266
timestamp 1
transform 1 0 25576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_283
timestamp 1
transform 1 0 27140 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_291
timestamp 1
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_296
timestamp 1636968456
transform 1 0 28336 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_311
timestamp 1
transform 1 0 29716 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1636968456
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636968456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636968456
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_365
timestamp 1636968456
transform 1 0 34684 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_377
timestamp 1636968456
transform 1 0 35788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636968456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636968456
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_417
timestamp 1
transform 1 0 39468 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_421
timestamp 1636968456
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1636968456
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636968456
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636968456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_473
timestamp 1
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1636968456
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1636968456
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636968456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636968456
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_529
timestamp 1
transform 1 0 49772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1636968456
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1636968456
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1636968456
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1636968456
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_585
timestamp 1
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_589
timestamp 1636968456
transform 1 0 55292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_601
timestamp 1636968456
transform 1 0 56396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_613
timestamp 1
transform 1 0 57500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1636968456
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1636968456
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_641
timestamp 1
transform 1 0 60076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_645
timestamp 1636968456
transform 1 0 60444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_657
timestamp 1636968456
transform 1 0 61548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_669
timestamp 1
transform 1 0 62652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1636968456
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1636968456
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_697
timestamp 1
transform 1 0 65228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_701
timestamp 1636968456
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_713
timestamp 1636968456
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_725
timestamp 1
transform 1 0 67804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1636968456
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1636968456
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_753
timestamp 1
transform 1 0 70380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_757
timestamp 1636968456
transform 1 0 70748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_769
timestamp 1636968456
transform 1 0 71852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_781
timestamp 1
transform 1 0 72956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1636968456
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1636968456
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_809
timestamp 1
transform 1 0 75532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_813
timestamp 1636968456
transform 1 0 75900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_825
timestamp 1636968456
transform 1 0 77004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_837
timestamp 1
transform 1 0 78108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1636968456
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1636968456
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_865
timestamp 1
transform 1 0 80684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_869
timestamp 1636968456
transform 1 0 81052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_881
timestamp 1636968456
transform 1 0 82156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_893
timestamp 1
transform 1 0 83260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1636968456
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1636968456
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_925
timestamp 1636968456
transform 1 0 86204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_937
timestamp 1636968456
transform 1 0 87308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_949
timestamp 1
transform 1 0 88412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1636968456
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_965
timestamp 1
transform 1 0 89884 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_971
timestamp 1
transform 1 0 90436 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_978
timestamp 1
transform 1 0 91080 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_981
timestamp 1636968456
transform 1 0 91356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_993
timestamp 1636968456
transform 1 0 92460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1005
timestamp 1
transform 1 0 93564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1636968456
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1636968456
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1033
timestamp 1
transform 1 0 96140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1636968456
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1049
timestamp 1636968456
transform 1 0 97612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1061
timestamp 1
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1636968456
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1636968456
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1089
timestamp 1
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1093
timestamp 1636968456
transform 1 0 101660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1105
timestamp 1636968456
transform 1 0 102764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1117
timestamp 1
transform 1 0 103868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1636968456
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1636968456
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1145
timestamp 1
transform 1 0 106444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1149
timestamp 1636968456
transform 1 0 106812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1161
timestamp 1
transform 1 0 107916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1167
timestamp 1
transform 1 0 108468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1636968456
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636968456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1122
timestamp 1636968456
transform 1 0 104328 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1134
timestamp 1636968456
transform 1 0 105432 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1146
timestamp 1
transform 1 0 106536 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1148
timestamp 1636968456
transform 1 0 106720 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_1160
timestamp 1
transform 1 0 107824 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636968456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1122
timestamp 1636968456
transform 1 0 104328 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1134
timestamp 1636968456
transform 1 0 105432 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1146
timestamp 1636968456
transform 1 0 106536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1158
timestamp 1
transform 1 0 107640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1166
timestamp 1
transform 1 0 108376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1636968456
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636968456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_65
timestamp 1
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1122
timestamp 1636968456
transform 1 0 104328 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1134
timestamp 1636968456
transform 1 0 105432 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1146
timestamp 1
transform 1 0 106536 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1148
timestamp 1636968456
transform 1 0 106720 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_1160
timestamp 1
transform 1 0 107824 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp 1
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1122
timestamp 1636968456
transform 1 0 104328 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1134
timestamp 1636968456
transform 1 0 105432 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1146
timestamp 1636968456
transform 1 0 106536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1158
timestamp 1
transform 1 0 107640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1166
timestamp 1
transform 1 0 108376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_11
timestamp 1636968456
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636968456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1122
timestamp 1636968456
transform 1 0 104328 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1134
timestamp 1636968456
transform 1 0 105432 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1146
timestamp 1
transform 1 0 106536 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1148
timestamp 1636968456
transform 1 0 106720 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_1160
timestamp 1
transform 1 0 107824 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1636968456
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1636968456
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1636968456
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1122
timestamp 1636968456
transform 1 0 104328 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1134
timestamp 1636968456
transform 1 0 105432 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1146
timestamp 1636968456
transform 1 0 106536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1158
timestamp 1
transform 1 0 107640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1166
timestamp 1
transform 1 0 108376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_11
timestamp 1636968456
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636968456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636968456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_65
timestamp 1
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1122
timestamp 1636968456
transform 1 0 104328 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1134
timestamp 1636968456
transform 1 0 105432 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1146
timestamp 1
transform 1 0 106536 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1148
timestamp 1636968456
transform 1 0 106720 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_1160
timestamp 1
transform 1 0 107824 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1636968456
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1636968456
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1636968456
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1122
timestamp 1636968456
transform 1 0 104328 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1134
timestamp 1636968456
transform 1 0 105432 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1146
timestamp 1636968456
transform 1 0 106536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1158
timestamp 1
transform 1 0 107640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1166
timestamp 1
transform 1 0 108376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636968456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636968456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_65
timestamp 1
transform 1 0 7084 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1122
timestamp 1636968456
transform 1 0 104328 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1134
timestamp 1636968456
transform 1 0 105432 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1146
timestamp 1
transform 1 0 106536 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1148
timestamp 1636968456
transform 1 0 106720 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_1160
timestamp 1
transform 1 0 107824 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_11
timestamp 1636968456
transform 1 0 2116 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_23
timestamp 1636968456
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1636968456
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636968456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1122
timestamp 1636968456
transform 1 0 104328 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1134
timestamp 1636968456
transform 1 0 105432 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1146
timestamp 1636968456
transform 1 0 106536 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1158
timestamp 1
transform 1 0 107640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1166
timestamp 1
transform 1 0 108376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1636968456
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636968456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636968456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_65
timestamp 1
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1122
timestamp 1636968456
transform 1 0 104328 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1134
timestamp 1636968456
transform 1 0 105432 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1146
timestamp 1
transform 1 0 106536 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1148
timestamp 1636968456
transform 1 0 106720 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_1160
timestamp 1
transform 1 0 107824 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_11
timestamp 1636968456
transform 1 0 2116 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1636968456
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_35
timestamp 1636968456
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636968456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1122
timestamp 1636968456
transform 1 0 104328 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1134
timestamp 1636968456
transform 1 0 105432 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1146
timestamp 1636968456
transform 1 0 106536 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1158
timestamp 1
transform 1 0 107640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_1166
timestamp 1
transform 1 0 108376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636968456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1122
timestamp 1636968456
transform 1 0 104328 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1134
timestamp 1636968456
transform 1 0 105432 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1146
timestamp 1
transform 1 0 106536 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1148
timestamp 1636968456
transform 1 0 106720 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_1160
timestamp 1
transform 1 0 107824 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636968456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636968456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1122
timestamp 1636968456
transform 1 0 104328 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1134
timestamp 1636968456
transform 1 0 105432 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1146
timestamp 1636968456
transform 1 0 106536 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1158
timestamp 1
transform 1 0 107640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_1166
timestamp 1
transform 1 0 108376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636968456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1122
timestamp 1636968456
transform 1 0 104328 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1134
timestamp 1636968456
transform 1 0 105432 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1146
timestamp 1
transform 1 0 106536 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1148
timestamp 1636968456
transform 1 0 106720 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_1160
timestamp 1
transform 1 0 107824 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636968456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636968456
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636968456
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1122
timestamp 1636968456
transform 1 0 104328 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1134
timestamp 1636968456
transform 1 0 105432 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1146
timestamp 1636968456
transform 1 0 106536 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1158
timestamp 1
transform 1 0 107640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_1166
timestamp 1
transform 1 0 108376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1122
timestamp 1636968456
transform 1 0 104328 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1134
timestamp 1636968456
transform 1 0 105432 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1146
timestamp 1
transform 1 0 106536 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1148
timestamp 1636968456
transform 1 0 106720 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_1160
timestamp 1
transform 1 0 107824 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636968456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636968456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1122
timestamp 1636968456
transform 1 0 104328 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1134
timestamp 1636968456
transform 1 0 105432 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1146
timestamp 1636968456
transform 1 0 106536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1158
timestamp 1
transform 1 0 107640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_1166
timestamp 1
transform 1 0 108376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636968456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_65
timestamp 1
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1122
timestamp 1636968456
transform 1 0 104328 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1134
timestamp 1636968456
transform 1 0 105432 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1146
timestamp 1
transform 1 0 106536 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1148
timestamp 1636968456
transform 1 0 106720 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_1160
timestamp 1
transform 1 0 107824 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636968456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636968456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636968456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1122
timestamp 1636968456
transform 1 0 104328 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1134
timestamp 1636968456
transform 1 0 105432 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1146
timestamp 1636968456
transform 1 0 106536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_1158
timestamp 1
transform 1 0 107640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_1166
timestamp 1
transform 1 0 108376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636968456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636968456
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1122
timestamp 1636968456
transform 1 0 104328 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1134
timestamp 1636968456
transform 1 0 105432 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1146
timestamp 1
transform 1 0 106536 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1148
timestamp 1636968456
transform 1 0 106720 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_1160
timestamp 1
transform 1 0 107824 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636968456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636968456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636968456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636968456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_69
timestamp 1
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1122
timestamp 1636968456
transform 1 0 104328 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1134
timestamp 1636968456
transform 1 0 105432 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1146
timestamp 1636968456
transform 1 0 106536 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1158
timestamp 1
transform 1 0 107640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1166
timestamp 1
transform 1 0 108376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636968456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636968456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636968456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636968456
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 1
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1122
timestamp 1636968456
transform 1 0 104328 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1134
timestamp 1636968456
transform 1 0 105432 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1146
timestamp 1
transform 1 0 106536 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1148
timestamp 1636968456
transform 1 0 106720 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_1160
timestamp 1
transform 1 0 107824 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636968456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636968456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636968456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636968456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1122
timestamp 1636968456
transform 1 0 104328 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1134
timestamp 1636968456
transform 1 0 105432 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1146
timestamp 1636968456
transform 1 0 106536 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_1158
timestamp 1
transform 1 0 107640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_1166
timestamp 1
transform 1 0 108376 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636968456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636968456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636968456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636968456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636968456
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_65
timestamp 1
transform 1 0 7084 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1122
timestamp 1636968456
transform 1 0 104328 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1134
timestamp 1636968456
transform 1 0 105432 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1146
timestamp 1
transform 1 0 106536 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1148
timestamp 1636968456
transform 1 0 106720 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_1160
timestamp 1
transform 1 0 107824 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636968456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636968456
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636968456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636968456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1122
timestamp 1636968456
transform 1 0 104328 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1134
timestamp 1636968456
transform 1 0 105432 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1146
timestamp 1636968456
transform 1 0 106536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1158
timestamp 1
transform 1 0 107640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_1166
timestamp 1
transform 1 0 108376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636968456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636968456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636968456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636968456
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_65
timestamp 1
transform 1 0 7084 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1122
timestamp 1636968456
transform 1 0 104328 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1134
timestamp 1636968456
transform 1 0 105432 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1146
timestamp 1
transform 1 0 106536 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1148
timestamp 1636968456
transform 1 0 106720 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_1160
timestamp 1
transform 1 0 107824 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636968456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636968456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636968456
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636968456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1124
timestamp 1636968456
transform 1 0 104512 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1136
timestamp 1636968456
transform 1 0 105616 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1148
timestamp 1636968456
transform 1 0 106720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1160
timestamp 1
transform 1 0 107824 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636968456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636968456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636968456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636968456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1122
timestamp 1636968456
transform 1 0 104328 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1134
timestamp 1636968456
transform 1 0 105432 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1146
timestamp 1
transform 1 0 106536 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1148
timestamp 1636968456
transform 1 0 106720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_1160
timestamp 1
transform 1 0 107824 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636968456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636968456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636968456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636968456
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636968456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_69
timestamp 1
transform 1 0 7452 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1124
timestamp 1636968456
transform 1 0 104512 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1136
timestamp 1636968456
transform 1 0 105616 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1148
timestamp 1636968456
transform 1 0 106720 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_1160
timestamp 1
transform 1 0 107824 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636968456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636968456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636968456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_65
timestamp 1
transform 1 0 7084 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1122
timestamp 1636968456
transform 1 0 104328 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1134
timestamp 1636968456
transform 1 0 105432 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1146
timestamp 1
transform 1 0 106536 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1148
timestamp 1636968456
transform 1 0 106720 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_1160
timestamp 1
transform 1 0 107824 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636968456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636968456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636968456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636968456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1122
timestamp 1636968456
transform 1 0 104328 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1134
timestamp 1636968456
transform 1 0 105432 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1146
timestamp 1636968456
transform 1 0 106536 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1158
timestamp 1
transform 1 0 107640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_1166
timestamp 1
transform 1 0 108376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636968456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636968456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636968456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636968456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1124
timestamp 1636968456
transform 1 0 104512 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1136
timestamp 1
transform 1 0 105616 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_1144
timestamp 1
transform 1 0 106352 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1148
timestamp 1636968456
transform 1 0 106720 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_1160
timestamp 1
transform 1 0 107824 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636968456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636968456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1122
timestamp 1636968456
transform 1 0 104328 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1134
timestamp 1636968456
transform 1 0 105432 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1146
timestamp 1636968456
transform 1 0 106536 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1158
timestamp 1
transform 1 0 107640 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_1166
timestamp 1
transform 1 0 108376 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636968456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636968456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_65
timestamp 1
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1122
timestamp 1636968456
transform 1 0 104328 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1134
timestamp 1636968456
transform 1 0 105432 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1146
timestamp 1
transform 1 0 106536 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1148
timestamp 1636968456
transform 1 0 106720 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_1160
timestamp 1
transform 1 0 107824 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636968456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636968456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636968456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1122
timestamp 1636968456
transform 1 0 104328 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1134
timestamp 1636968456
transform 1 0 105432 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1146
timestamp 1636968456
transform 1 0 106536 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1158
timestamp 1
transform 1 0 107640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1166
timestamp 1
transform 1 0 108376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_65
timestamp 1
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1122
timestamp 1636968456
transform 1 0 104328 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1134
timestamp 1636968456
transform 1 0 105432 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1146
timestamp 1
transform 1 0 106536 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1148
timestamp 1636968456
transform 1 0 106720 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1160
timestamp 1
transform 1 0 107824 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_69
timestamp 1
transform 1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1122
timestamp 1636968456
transform 1 0 104328 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1134
timestamp 1636968456
transform 1 0 105432 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1146
timestamp 1636968456
transform 1 0 106536 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1158
timestamp 1
transform 1 0 107640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_1166
timestamp 1
transform 1 0 108376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_65
timestamp 1
transform 1 0 7084 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1122
timestamp 1636968456
transform 1 0 104328 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1134
timestamp 1636968456
transform 1 0 105432 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1146
timestamp 1
transform 1 0 106536 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1148
timestamp 1636968456
transform 1 0 106720 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_1160
timestamp 1
transform 1 0 107824 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636968456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636968456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636968456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1636968456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636968456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1
transform 1 0 7452 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1122
timestamp 1636968456
transform 1 0 104328 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1134
timestamp 1636968456
transform 1 0 105432 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1146
timestamp 1636968456
transform 1 0 106536 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_1158
timestamp 1
transform 1 0 107640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_1166
timestamp 1
transform 1 0 108376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636968456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_65
timestamp 1
transform 1 0 7084 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1122
timestamp 1636968456
transform 1 0 104328 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1134
timestamp 1636968456
transform 1 0 105432 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1146
timestamp 1
transform 1 0 106536 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1148
timestamp 1636968456
transform 1 0 106720 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1160
timestamp 1
transform 1 0 107824 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636968456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636968456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_69
timestamp 1
transform 1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1122
timestamp 1636968456
transform 1 0 104328 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1134
timestamp 1636968456
transform 1 0 105432 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1146
timestamp 1636968456
transform 1 0 106536 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1158
timestamp 1
transform 1 0 107640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1166
timestamp 1
transform 1 0 108376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636968456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636968456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_65
timestamp 1
transform 1 0 7084 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1122
timestamp 1636968456
transform 1 0 104328 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1134
timestamp 1636968456
transform 1 0 105432 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1146
timestamp 1
transform 1 0 106536 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1148
timestamp 1636968456
transform 1 0 106720 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_1160
timestamp 1
transform 1 0 107824 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636968456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636968456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636968456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1636968456
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_69
timestamp 1
transform 1 0 7452 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1122
timestamp 1636968456
transform 1 0 104328 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1134
timestamp 1636968456
transform 1 0 105432 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1146
timestamp 1636968456
transform 1 0 106536 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_1158
timestamp 1
transform 1 0 107640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_1166
timestamp 1
transform 1 0 108376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636968456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636968456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636968456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1636968456
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1636968456
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_65
timestamp 1
transform 1 0 7084 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1122
timestamp 1636968456
transform 1 0 104328 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1134
timestamp 1636968456
transform 1 0 105432 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1146
timestamp 1
transform 1 0 106536 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1148
timestamp 1636968456
transform 1 0 106720 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_1160
timestamp 1
transform 1 0 107824 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636968456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636968456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1636968456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1636968456
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1636968456
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_69
timestamp 1
transform 1 0 7452 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1122
timestamp 1636968456
transform 1 0 104328 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1134
timestamp 1636968456
transform 1 0 105432 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1146
timestamp 1636968456
transform 1 0 106536 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_1158
timestamp 1
transform 1 0 107640 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1166
timestamp 1
transform 1 0 108376 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636968456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636968456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636968456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636968456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1636968456
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_65
timestamp 1
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1122
timestamp 1636968456
transform 1 0 104328 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1134
timestamp 1636968456
transform 1 0 105432 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1146
timestamp 1
transform 1 0 106536 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1148
timestamp 1636968456
transform 1 0 106720 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_1160
timestamp 1
transform 1 0 107824 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636968456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636968456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636968456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636968456
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636968456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_69
timestamp 1
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1122
timestamp 1636968456
transform 1 0 104328 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1134
timestamp 1636968456
transform 1 0 105432 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1146
timestamp 1636968456
transform 1 0 106536 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_1158
timestamp 1
transform 1 0 107640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_1166
timestamp 1
transform 1 0 108376 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636968456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636968456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636968456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636968456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636968456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_65
timestamp 1
transform 1 0 7084 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1122
timestamp 1636968456
transform 1 0 104328 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1134
timestamp 1636968456
transform 1 0 105432 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1146
timestamp 1
transform 1 0 106536 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1148
timestamp 1636968456
transform 1 0 106720 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_1160
timestamp 1
transform 1 0 107824 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636968456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636968456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636968456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636968456
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636968456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_69
timestamp 1
transform 1 0 7452 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1122
timestamp 1636968456
transform 1 0 104328 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1134
timestamp 1636968456
transform 1 0 105432 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1146
timestamp 1636968456
transform 1 0 106536 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1158
timestamp 1
transform 1 0 107640 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1166
timestamp 1
transform 1 0 108376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636968456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636968456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636968456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636968456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636968456
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_65
timestamp 1
transform 1 0 7084 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1122
timestamp 1636968456
transform 1 0 104328 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1134
timestamp 1636968456
transform 1 0 105432 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1146
timestamp 1
transform 1 0 106536 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1148
timestamp 1636968456
transform 1 0 106720 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_1160
timestamp 1
transform 1 0 107824 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636968456
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636968456
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1636968456
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1636968456
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636968456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1122
timestamp 1636968456
transform 1 0 104328 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1134
timestamp 1636968456
transform 1 0 105432 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1146
timestamp 1636968456
transform 1 0 106536 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1158
timestamp 1
transform 1 0 107640 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1166
timestamp 1
transform 1 0 108376 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636968456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636968456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636968456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636968456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1636968456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_65
timestamp 1
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1122
timestamp 1636968456
transform 1 0 104328 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1134
timestamp 1636968456
transform 1 0 105432 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1146
timestamp 1
transform 1 0 106536 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1148
timestamp 1636968456
transform 1 0 106720 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1160
timestamp 1
transform 1 0 107824 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636968456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636968456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1636968456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1636968456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1636968456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1122
timestamp 1636968456
transform 1 0 104328 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1134
timestamp 1636968456
transform 1 0 105432 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1146
timestamp 1636968456
transform 1 0 106536 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1158
timestamp 1
transform 1 0 107640 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1166
timestamp 1
transform 1 0 108376 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636968456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636968456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636968456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1636968456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1636968456
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_65
timestamp 1
transform 1 0 7084 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1122
timestamp 1636968456
transform 1 0 104328 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1134
timestamp 1636968456
transform 1 0 105432 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1146
timestamp 1
transform 1 0 106536 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1148
timestamp 1636968456
transform 1 0 106720 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_1160
timestamp 1
transform 1 0 107824 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1636968456
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1636968456
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1636968456
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1636968456
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1636968456
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_69
timestamp 1
transform 1 0 7452 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1122
timestamp 1636968456
transform 1 0 104328 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1134
timestamp 1636968456
transform 1 0 105432 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1146
timestamp 1636968456
transform 1 0 106536 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_1158
timestamp 1
transform 1 0 107640 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_1166
timestamp 1
transform 1 0 108376 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636968456
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636968456
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636968456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1636968456
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1636968456
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_65
timestamp 1
transform 1 0 7084 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1122
timestamp 1636968456
transform 1 0 104328 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1134
timestamp 1636968456
transform 1 0 105432 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1146
timestamp 1
transform 1 0 106536 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1148
timestamp 1636968456
transform 1 0 106720 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_1160
timestamp 1
transform 1 0 107824 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636968456
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636968456
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1636968456
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1636968456
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636968456
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1122
timestamp 1636968456
transform 1 0 104328 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1134
timestamp 1636968456
transform 1 0 105432 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1146
timestamp 1636968456
transform 1 0 106536 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1158
timestamp 1
transform 1 0 107640 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_1166
timestamp 1
transform 1 0 108376 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636968456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636968456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636968456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636968456
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636968456
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_65
timestamp 1
transform 1 0 7084 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1122
timestamp 1636968456
transform 1 0 104328 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1134
timestamp 1636968456
transform 1 0 105432 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1146
timestamp 1
transform 1 0 106536 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1148
timestamp 1636968456
transform 1 0 106720 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_1160
timestamp 1
transform 1 0 107824 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636968456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636968456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636968456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636968456
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636968456
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1122
timestamp 1636968456
transform 1 0 104328 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1134
timestamp 1636968456
transform 1 0 105432 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1146
timestamp 1636968456
transform 1 0 106536 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_1158
timestamp 1
transform 1 0 107640 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_1166
timestamp 1
transform 1 0 108376 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636968456
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636968456
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636968456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636968456
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636968456
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_65
timestamp 1
transform 1 0 7084 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1122
timestamp 1636968456
transform 1 0 104328 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1134
timestamp 1636968456
transform 1 0 105432 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1146
timestamp 1
transform 1 0 106536 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1148
timestamp 1636968456
transform 1 0 106720 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_1160
timestamp 1
transform 1 0 107824 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636968456
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636968456
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636968456
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636968456
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636968456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_69
timestamp 1
transform 1 0 7452 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1122
timestamp 1636968456
transform 1 0 104328 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1134
timestamp 1636968456
transform 1 0 105432 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1146
timestamp 1636968456
transform 1 0 106536 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_1158
timestamp 1
transform 1 0 107640 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1166
timestamp 1
transform 1 0 108376 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636968456
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636968456
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636968456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636968456
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636968456
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_65
timestamp 1
transform 1 0 7084 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1122
timestamp 1636968456
transform 1 0 104328 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1134
timestamp 1636968456
transform 1 0 105432 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_1146
timestamp 1
transform 1 0 106536 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1148
timestamp 1636968456
transform 1 0 106720 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_1160
timestamp 1
transform 1 0 107824 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636968456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636968456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636968456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636968456
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636968456
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_69
timestamp 1
transform 1 0 7452 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1122
timestamp 1636968456
transform 1 0 104328 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1134
timestamp 1636968456
transform 1 0 105432 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1146
timestamp 1636968456
transform 1 0 106536 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_1158
timestamp 1
transform 1 0 107640 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_1166
timestamp 1
transform 1 0 108376 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636968456
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636968456
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636968456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636968456
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636968456
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_65
timestamp 1
transform 1 0 7084 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1122
timestamp 1636968456
transform 1 0 104328 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1134
timestamp 1636968456
transform 1 0 105432 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1146
timestamp 1
transform 1 0 106536 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1148
timestamp 1636968456
transform 1 0 106720 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_1160
timestamp 1
transform 1 0 107824 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636968456
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636968456
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1636968456
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1636968456
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636968456
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_69
timestamp 1
transform 1 0 7452 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1122
timestamp 1636968456
transform 1 0 104328 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1134
timestamp 1636968456
transform 1 0 105432 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1146
timestamp 1636968456
transform 1 0 106536 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_1158
timestamp 1
transform 1 0 107640 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_1166
timestamp 1
transform 1 0 108376 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636968456
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636968456
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636968456
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1636968456
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1636968456
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_65
timestamp 1
transform 1 0 7084 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1122
timestamp 1636968456
transform 1 0 104328 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1134
timestamp 1636968456
transform 1 0 105432 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1146
timestamp 1
transform 1 0 106536 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1148
timestamp 1636968456
transform 1 0 106720 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_1160
timestamp 1
transform 1 0 107824 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636968456
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636968456
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1636968456
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1636968456
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1636968456
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_69
timestamp 1
transform 1 0 7452 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1122
timestamp 1636968456
transform 1 0 104328 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1134
timestamp 1636968456
transform 1 0 105432 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1146
timestamp 1636968456
transform 1 0 106536 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_1158
timestamp 1
transform 1 0 107640 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_1166
timestamp 1
transform 1 0 108376 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636968456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636968456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636968456
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1636968456
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1636968456
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_65
timestamp 1
transform 1 0 7084 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1122
timestamp 1636968456
transform 1 0 104328 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1134
timestamp 1636968456
transform 1 0 105432 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_1146
timestamp 1
transform 1 0 106536 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1148
timestamp 1636968456
transform 1 0 106720 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_1160
timestamp 1
transform 1 0 107824 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636968456
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636968456
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636968456
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1636968456
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1636968456
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_69
timestamp 1
transform 1 0 7452 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1122
timestamp 1636968456
transform 1 0 104328 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1134
timestamp 1636968456
transform 1 0 105432 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1146
timestamp 1636968456
transform 1 0 106536 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_1158
timestamp 1
transform 1 0 107640 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_1166
timestamp 1
transform 1 0 108376 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636968456
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636968456
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636968456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1636968456
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1636968456
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_65
timestamp 1
transform 1 0 7084 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1122
timestamp 1636968456
transform 1 0 104328 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1134
timestamp 1636968456
transform 1 0 105432 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1146
timestamp 1
transform 1 0 106536 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1148
timestamp 1636968456
transform 1 0 106720 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_1160
timestamp 1
transform 1 0 107824 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636968456
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636968456
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1636968456
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1636968456
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1636968456
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_69
timestamp 1
transform 1 0 7452 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1122
timestamp 1636968456
transform 1 0 104328 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1134
timestamp 1636968456
transform 1 0 105432 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1146
timestamp 1636968456
transform 1 0 106536 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_1158
timestamp 1
transform 1 0 107640 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_1166
timestamp 1
transform 1 0 108376 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636968456
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636968456
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636968456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1636968456
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1636968456
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_65
timestamp 1
transform 1 0 7084 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1122
timestamp 1636968456
transform 1 0 104328 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1134
timestamp 1636968456
transform 1 0 105432 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1146
timestamp 1
transform 1 0 106536 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1148
timestamp 1636968456
transform 1 0 106720 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_1160
timestamp 1
transform 1 0 107824 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636968456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636968456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636968456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1636968456
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1636968456
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_69
timestamp 1
transform 1 0 7452 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1122
timestamp 1636968456
transform 1 0 104328 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1134
timestamp 1636968456
transform 1 0 105432 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1146
timestamp 1636968456
transform 1 0 106536 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_1158
timestamp 1
transform 1 0 107640 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_1166
timestamp 1
transform 1 0 108376 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636968456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636968456
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636968456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1636968456
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1636968456
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_65
timestamp 1
transform 1 0 7084 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1122
timestamp 1636968456
transform 1 0 104328 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1134
timestamp 1636968456
transform 1 0 105432 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_1146
timestamp 1
transform 1 0 106536 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1148
timestamp 1636968456
transform 1 0 106720 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_1160
timestamp 1
transform 1 0 107824 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1636968456
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1636968456
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1636968456
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1636968456
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1636968456
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_69
timestamp 1
transform 1 0 7452 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1122
timestamp 1636968456
transform 1 0 104328 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1134
timestamp 1636968456
transform 1 0 105432 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1146
timestamp 1636968456
transform 1 0 106536 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_1158
timestamp 1
transform 1 0 107640 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_1166
timestamp 1
transform 1 0 108376 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636968456
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636968456
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636968456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1636968456
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1636968456
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_65
timestamp 1
transform 1 0 7084 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1122
timestamp 1636968456
transform 1 0 104328 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1134
timestamp 1636968456
transform 1 0 105432 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_1146
timestamp 1
transform 1 0 106536 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1148
timestamp 1636968456
transform 1 0 106720 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_1160
timestamp 1
transform 1 0 107824 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636968456
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636968456
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1636968456
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1636968456
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1636968456
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_69
timestamp 1
transform 1 0 7452 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1122
timestamp 1636968456
transform 1 0 104328 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1134
timestamp 1636968456
transform 1 0 105432 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1146
timestamp 1636968456
transform 1 0 106536 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_1158
timestamp 1
transform 1 0 107640 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_1166
timestamp 1
transform 1 0 108376 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636968456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636968456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636968456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1636968456
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1636968456
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_65
timestamp 1
transform 1 0 7084 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1122
timestamp 1636968456
transform 1 0 104328 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1134
timestamp 1636968456
transform 1 0 105432 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_1146
timestamp 1
transform 1 0 106536 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1148
timestamp 1636968456
transform 1 0 106720 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_1160
timestamp 1
transform 1 0 107824 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636968456
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636968456
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1636968456
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1636968456
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1636968456
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_69
timestamp 1
transform 1 0 7452 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1122
timestamp 1636968456
transform 1 0 104328 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1134
timestamp 1636968456
transform 1 0 105432 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1146
timestamp 1636968456
transform 1 0 106536 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_1158
timestamp 1
transform 1 0 107640 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_1166
timestamp 1
transform 1 0 108376 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1636968456
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1636968456
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636968456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1636968456
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1636968456
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_65
timestamp 1
transform 1 0 7084 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1122
timestamp 1636968456
transform 1 0 104328 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1134
timestamp 1636968456
transform 1 0 105432 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_1146
timestamp 1
transform 1 0 106536 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1148
timestamp 1636968456
transform 1 0 106720 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_1160
timestamp 1
transform 1 0 107824 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636968456
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636968456
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1636968456
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1636968456
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1636968456
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_69
timestamp 1
transform 1 0 7452 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1122
timestamp 1636968456
transform 1 0 104328 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1134
timestamp 1636968456
transform 1 0 105432 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1146
timestamp 1636968456
transform 1 0 106536 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_1158
timestamp 1
transform 1 0 107640 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_1166
timestamp 1
transform 1 0 108376 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1636968456
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1636968456
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636968456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1636968456
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1636968456
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_65
timestamp 1
transform 1 0 7084 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1122
timestamp 1636968456
transform 1 0 104328 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1134
timestamp 1636968456
transform 1 0 105432 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_1146
timestamp 1
transform 1 0 106536 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1148
timestamp 1636968456
transform 1 0 106720 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_1160
timestamp 1
transform 1 0 107824 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636968456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636968456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636968456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1636968456
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1636968456
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_69
timestamp 1
transform 1 0 7452 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1122
timestamp 1636968456
transform 1 0 104328 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1134
timestamp 1636968456
transform 1 0 105432 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1146
timestamp 1636968456
transform 1 0 106536 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_1158
timestamp 1
transform 1 0 107640 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_1166
timestamp 1
transform 1 0 108376 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636968456
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636968456
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636968456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1636968456
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1636968456
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_65
timestamp 1
transform 1 0 7084 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1122
timestamp 1636968456
transform 1 0 104328 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1134
timestamp 1636968456
transform 1 0 105432 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_1146
timestamp 1
transform 1 0 106536 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1148
timestamp 1636968456
transform 1 0 106720 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_1160
timestamp 1
transform 1 0 107824 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1636968456
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1636968456
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1636968456
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1636968456
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1636968456
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_69
timestamp 1
transform 1 0 7452 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1122
timestamp 1636968456
transform 1 0 104328 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1134
timestamp 1636968456
transform 1 0 105432 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1146
timestamp 1636968456
transform 1 0 106536 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_1158
timestamp 1
transform 1 0 107640 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_1166
timestamp 1
transform 1 0 108376 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636968456
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636968456
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636968456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1636968456
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1636968456
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_65
timestamp 1
transform 1 0 7084 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1122
timestamp 1636968456
transform 1 0 104328 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1134
timestamp 1636968456
transform 1 0 105432 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_1146
timestamp 1
transform 1 0 106536 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1148
timestamp 1636968456
transform 1 0 106720 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_1160
timestamp 1
transform 1 0 107824 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636968456
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636968456
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1636968456
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1636968456
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1636968456
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_69
timestamp 1
transform 1 0 7452 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1122
timestamp 1636968456
transform 1 0 104328 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1134
timestamp 1636968456
transform 1 0 105432 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1146
timestamp 1636968456
transform 1 0 106536 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_1158
timestamp 1
transform 1 0 107640 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_1166
timestamp 1
transform 1 0 108376 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636968456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636968456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636968456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1636968456
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1636968456
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_65
timestamp 1
transform 1 0 7084 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1122
timestamp 1636968456
transform 1 0 104328 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1134
timestamp 1636968456
transform 1 0 105432 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_1146
timestamp 1
transform 1 0 106536 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1148
timestamp 1636968456
transform 1 0 106720 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_1160
timestamp 1
transform 1 0 107824 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636968456
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636968456
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1636968456
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1636968456
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1636968456
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_69
timestamp 1
transform 1 0 7452 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1122
timestamp 1636968456
transform 1 0 104328 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1134
timestamp 1636968456
transform 1 0 105432 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1146
timestamp 1636968456
transform 1 0 106536 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_1158
timestamp 1
transform 1 0 107640 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_1166
timestamp 1
transform 1 0 108376 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1636968456
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1636968456
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1636968456
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1636968456
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1636968456
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_65
timestamp 1
transform 1 0 7084 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1122
timestamp 1636968456
transform 1 0 104328 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1134
timestamp 1636968456
transform 1 0 105432 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_1146
timestamp 1
transform 1 0 106536 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1148
timestamp 1636968456
transform 1 0 106720 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_1160
timestamp 1
transform 1 0 107824 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636968456
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636968456
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_27
timestamp 1636968456
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1636968456
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1636968456
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_69
timestamp 1
transform 1 0 7452 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1122
timestamp 1636968456
transform 1 0 104328 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1134
timestamp 1636968456
transform 1 0 105432 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1146
timestamp 1636968456
transform 1 0 106536 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_1158
timestamp 1
transform 1 0 107640 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_1166
timestamp 1
transform 1 0 108376 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1636968456
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1636968456
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1636968456
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1636968456
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1636968456
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_65
timestamp 1
transform 1 0 7084 0 1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1122
timestamp 1636968456
transform 1 0 104328 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1134
timestamp 1636968456
transform 1 0 105432 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_1146
timestamp 1
transform 1 0 106536 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1148
timestamp 1636968456
transform 1 0 106720 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_1160
timestamp 1
transform 1 0 107824 0 1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636968456
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636968456
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1636968456
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_39
timestamp 1636968456
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1636968456
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_69
timestamp 1
transform 1 0 7452 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1122
timestamp 1636968456
transform 1 0 104328 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1134
timestamp 1636968456
transform 1 0 105432 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1146
timestamp 1636968456
transform 1 0 106536 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_1158
timestamp 1
transform 1 0 107640 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_1166
timestamp 1
transform 1 0 108376 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1636968456
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1636968456
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1636968456
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1636968456
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1636968456
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_65
timestamp 1
transform 1 0 7084 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1122
timestamp 1636968456
transform 1 0 104328 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1134
timestamp 1636968456
transform 1 0 105432 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_1146
timestamp 1
transform 1 0 106536 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1148
timestamp 1636968456
transform 1 0 106720 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_1160
timestamp 1
transform 1 0 107824 0 1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_105_3
timestamp 1636968456
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_15
timestamp 1636968456
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_27
timestamp 1636968456
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_39
timestamp 1636968456
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1636968456
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_69
timestamp 1
transform 1 0 7452 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1122
timestamp 1636968456
transform 1 0 104328 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1134
timestamp 1636968456
transform 1 0 105432 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1146
timestamp 1636968456
transform 1 0 106536 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_1158
timestamp 1
transform 1 0 107640 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_1166
timestamp 1
transform 1 0 108376 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636968456
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636968456
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636968456
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1636968456
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1636968456
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_65
timestamp 1
transform 1 0 7084 0 1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1125
timestamp 1636968456
transform 1 0 104604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_1137
timestamp 1
transform 1 0 105708 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_1145
timestamp 1
transform 1 0 106444 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1148
timestamp 1636968456
transform 1 0 106720 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_1160
timestamp 1
transform 1 0 107824 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636968456
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636968456
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1636968456
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_39
timestamp 1636968456
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1636968456
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_69
timestamp 1
transform 1 0 7452 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1122
timestamp 1636968456
transform 1 0 104328 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1134
timestamp 1636968456
transform 1 0 105432 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1146
timestamp 1636968456
transform 1 0 106536 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_1158
timestamp 1
transform 1 0 107640 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_1166
timestamp 1
transform 1 0 108376 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636968456
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636968456
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636968456
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1636968456
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1636968456
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_65
timestamp 1
transform 1 0 7084 0 1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1122
timestamp 1636968456
transform 1 0 104328 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1134
timestamp 1636968456
transform 1 0 105432 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_1146
timestamp 1
transform 1 0 106536 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1148
timestamp 1636968456
transform 1 0 106720 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_1160
timestamp 1
transform 1 0 107824 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1636968456
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1636968456
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_27
timestamp 1636968456
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_39
timestamp 1636968456
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1636968456
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_69
timestamp 1
transform 1 0 7452 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1122
timestamp 1636968456
transform 1 0 104328 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1134
timestamp 1636968456
transform 1 0 105432 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1146
timestamp 1636968456
transform 1 0 106536 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_1158
timestamp 1
transform 1 0 107640 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_1166
timestamp 1
transform 1 0 108376 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_110_3
timestamp 1636968456
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_15
timestamp 1636968456
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636968456
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1636968456
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1636968456
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_65
timestamp 1
transform 1 0 7084 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1122
timestamp 1636968456
transform 1 0 104328 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1134
timestamp 1636968456
transform 1 0 105432 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_1146
timestamp 1
transform 1 0 106536 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1148
timestamp 1636968456
transform 1 0 106720 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_1160
timestamp 1
transform 1 0 107824 0 1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636968456
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636968456
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1636968456
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_39
timestamp 1636968456
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1636968456
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_69
timestamp 1
transform 1 0 7452 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1122
timestamp 1636968456
transform 1 0 104328 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1134
timestamp 1636968456
transform 1 0 105432 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1146
timestamp 1636968456
transform 1 0 106536 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_1158
timestamp 1
transform 1 0 107640 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_111_1166
timestamp 1
transform 1 0 108376 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1636968456
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1636968456
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636968456
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1636968456
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1636968456
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_65
timestamp 1
transform 1 0 7084 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1122
timestamp 1636968456
transform 1 0 104328 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1134
timestamp 1636968456
transform 1 0 105432 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_1146
timestamp 1
transform 1 0 106536 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1148
timestamp 1636968456
transform 1 0 106720 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_1160
timestamp 1
transform 1 0 107824 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636968456
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636968456
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636968456
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1636968456
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1636968456
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_69
timestamp 1
transform 1 0 7452 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1122
timestamp 1636968456
transform 1 0 104328 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1134
timestamp 1636968456
transform 1 0 105432 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1146
timestamp 1636968456
transform 1 0 106536 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_1158
timestamp 1
transform 1 0 107640 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_113_1166
timestamp 1
transform 1 0 108376 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636968456
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636968456
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636968456
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1636968456
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1636968456
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_65
timestamp 1
transform 1 0 7084 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1122
timestamp 1636968456
transform 1 0 104328 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1134
timestamp 1636968456
transform 1 0 105432 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_1146
timestamp 1
transform 1 0 106536 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1148
timestamp 1636968456
transform 1 0 106720 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_1160
timestamp 1
transform 1 0 107824 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_115_3
timestamp 1636968456
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_15
timestamp 1636968456
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_27
timestamp 1636968456
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_39
timestamp 1636968456
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1636968456
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_115_69
timestamp 1
transform 1 0 7452 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1122
timestamp 1636968456
transform 1 0 104328 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1134
timestamp 1636968456
transform 1 0 105432 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1146
timestamp 1636968456
transform 1 0 106536 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_1158
timestamp 1
transform 1 0 107640 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_115_1166
timestamp 1
transform 1 0 108376 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636968456
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636968456
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636968456
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1636968456
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_53
timestamp 1636968456
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_65
timestamp 1
transform 1 0 7084 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1122
timestamp 1636968456
transform 1 0 104328 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1134
timestamp 1636968456
transform 1 0 105432 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_1146
timestamp 1
transform 1 0 106536 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1148
timestamp 1636968456
transform 1 0 106720 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_1160
timestamp 1
transform 1 0 107824 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636968456
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636968456
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_27
timestamp 1
transform 1 0 3588 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_29
timestamp 1636968456
transform 1 0 3772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_41
timestamp 1636968456
transform 1 0 4876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_53
timestamp 1
transform 1 0 5980 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1636968456
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1636968456
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_81
timestamp 1
transform 1 0 8556 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_85
timestamp 1636968456
transform 1 0 8924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_97
timestamp 1636968456
transform 1 0 10028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_109
timestamp 1
transform 1 0 11132 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1636968456
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_125
timestamp 1636968456
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_137
timestamp 1
transform 1 0 13708 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_141
timestamp 1636968456
transform 1 0 14076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_153
timestamp 1636968456
transform 1 0 15180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_165
timestamp 1
transform 1 0 16284 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_169
timestamp 1636968456
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_181
timestamp 1636968456
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_193
timestamp 1
transform 1 0 18860 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_197
timestamp 1636968456
transform 1 0 19228 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_209
timestamp 1636968456
transform 1 0 20332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_221
timestamp 1
transform 1 0 21436 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_225
timestamp 1636968456
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_237
timestamp 1636968456
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_249
timestamp 1
transform 1 0 24012 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_253
timestamp 1636968456
transform 1 0 24380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_265
timestamp 1636968456
transform 1 0 25484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_277
timestamp 1
transform 1 0 26588 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_281
timestamp 1636968456
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_293
timestamp 1636968456
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_305
timestamp 1
transform 1 0 29164 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_309
timestamp 1636968456
transform 1 0 29532 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_321
timestamp 1636968456
transform 1 0 30636 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_333
timestamp 1
transform 1 0 31740 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_337
timestamp 1636968456
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_349
timestamp 1636968456
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_361
timestamp 1
transform 1 0 34316 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_365
timestamp 1636968456
transform 1 0 34684 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_377
timestamp 1636968456
transform 1 0 35788 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_389
timestamp 1
transform 1 0 36892 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_393
timestamp 1636968456
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_405
timestamp 1636968456
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_417
timestamp 1
transform 1 0 39468 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_421
timestamp 1636968456
transform 1 0 39836 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_433
timestamp 1636968456
transform 1 0 40940 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_445
timestamp 1
transform 1 0 42044 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_449
timestamp 1636968456
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_461
timestamp 1636968456
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_473
timestamp 1
transform 1 0 44620 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_477
timestamp 1636968456
transform 1 0 44988 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_489
timestamp 1636968456
transform 1 0 46092 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_501
timestamp 1
transform 1 0 47196 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_505
timestamp 1636968456
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_517
timestamp 1636968456
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_529
timestamp 1
transform 1 0 49772 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_533
timestamp 1636968456
transform 1 0 50140 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_545
timestamp 1636968456
transform 1 0 51244 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_557
timestamp 1
transform 1 0 52348 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_561
timestamp 1636968456
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_573
timestamp 1636968456
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_585
timestamp 1
transform 1 0 54924 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_589
timestamp 1636968456
transform 1 0 55292 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_601
timestamp 1636968456
transform 1 0 56396 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_613
timestamp 1
transform 1 0 57500 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_617
timestamp 1636968456
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_629
timestamp 1636968456
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_641
timestamp 1
transform 1 0 60076 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_645
timestamp 1636968456
transform 1 0 60444 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_657
timestamp 1636968456
transform 1 0 61548 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_669
timestamp 1
transform 1 0 62652 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_673
timestamp 1636968456
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_685
timestamp 1636968456
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_697
timestamp 1
transform 1 0 65228 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_701
timestamp 1636968456
transform 1 0 65596 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_713
timestamp 1636968456
transform 1 0 66700 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_725
timestamp 1
transform 1 0 67804 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_729
timestamp 1
transform 1 0 68172 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_735
timestamp 1636968456
transform 1 0 68724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_747
timestamp 1
transform 1 0 69828 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_755
timestamp 1
transform 1 0 70564 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_757
timestamp 1636968456
transform 1 0 70748 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_769
timestamp 1636968456
transform 1 0 71852 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_781
timestamp 1
transform 1 0 72956 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_798
timestamp 1636968456
transform 1 0 74520 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_810
timestamp 1
transform 1 0 75624 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_813
timestamp 1636968456
transform 1 0 75900 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_825
timestamp 1636968456
transform 1 0 77004 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_837
timestamp 1
transform 1 0 78108 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_841
timestamp 1636968456
transform 1 0 78476 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_853
timestamp 1636968456
transform 1 0 79580 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_865
timestamp 1
transform 1 0 80684 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_869
timestamp 1636968456
transform 1 0 81052 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_881
timestamp 1636968456
transform 1 0 82156 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_893
timestamp 1
transform 1 0 83260 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_897
timestamp 1636968456
transform 1 0 83628 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_909
timestamp 1636968456
transform 1 0 84732 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_921
timestamp 1
transform 1 0 85836 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_953
timestamp 1
transform 1 0 88780 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_117_959
timestamp 1
transform 1 0 89332 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_979
timestamp 1
transform 1 0 91172 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_117_983
timestamp 1
transform 1 0 91540 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_992
timestamp 1636968456
transform 1 0 92368 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_1004
timestamp 1
transform 1 0 93472 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_117_1051
timestamp 1
transform 1 0 97796 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_117_1062
timestamp 1
transform 1 0 98808 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_117_1072
timestamp 1
transform 1 0 99728 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1076
timestamp 1
transform 1 0 100096 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_1084
timestamp 1
transform 1 0 100832 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1091
timestamp 1
transform 1 0 101476 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1104
timestamp 1636968456
transform 1 0 102672 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1116
timestamp 1
transform 1 0 103776 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1121
timestamp 1636968456
transform 1 0 104236 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1133
timestamp 1636968456
transform 1 0 105340 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1145
timestamp 1
transform 1 0 106444 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1149
timestamp 1636968456
transform 1 0 106812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_1161
timestamp 1
transform 1 0 107916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1167
timestamp 1
transform 1 0 108468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636968456
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636968456
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636968456
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1636968456
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1636968456
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1636968456
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1636968456
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1636968456
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1636968456
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1636968456
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1636968456
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1636968456
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_165
timestamp 1636968456
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_177
timestamp 1636968456
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_197
timestamp 1636968456
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_209
timestamp 1636968456
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_221
timestamp 1636968456
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_233
timestamp 1636968456
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_253
timestamp 1636968456
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_265
timestamp 1636968456
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_277
timestamp 1636968456
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_289
timestamp 1636968456
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_309
timestamp 1636968456
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_321
timestamp 1636968456
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_333
timestamp 1636968456
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_345
timestamp 1636968456
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_365
timestamp 1636968456
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_377
timestamp 1636968456
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_389
timestamp 1636968456
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_401
timestamp 1636968456
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_421
timestamp 1636968456
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_433
timestamp 1636968456
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_445
timestamp 1636968456
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_457
timestamp 1636968456
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_477
timestamp 1636968456
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_489
timestamp 1636968456
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_501
timestamp 1636968456
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_513
timestamp 1636968456
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_533
timestamp 1636968456
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_545
timestamp 1636968456
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_557
timestamp 1636968456
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_569
timestamp 1636968456
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_589
timestamp 1636968456
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_601
timestamp 1636968456
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_613
timestamp 1636968456
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_625
timestamp 1636968456
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_645
timestamp 1636968456
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_657
timestamp 1636968456
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_669
timestamp 1636968456
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_681
timestamp 1636968456
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_701
timestamp 1636968456
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_713
timestamp 1636968456
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_725
timestamp 1636968456
transform 1 0 67804 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_737
timestamp 1636968456
transform 1 0 68908 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_749
timestamp 1
transform 1 0 70012 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_755
timestamp 1
transform 1 0 70564 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_757
timestamp 1636968456
transform 1 0 70748 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_769
timestamp 1636968456
transform 1 0 71852 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_781
timestamp 1636968456
transform 1 0 72956 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_793
timestamp 1636968456
transform 1 0 74060 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_805
timestamp 1
transform 1 0 75164 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_811
timestamp 1
transform 1 0 75716 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_813
timestamp 1636968456
transform 1 0 75900 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_825
timestamp 1636968456
transform 1 0 77004 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_837
timestamp 1636968456
transform 1 0 78108 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_849
timestamp 1636968456
transform 1 0 79212 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_861
timestamp 1
transform 1 0 80316 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_867
timestamp 1
transform 1 0 80868 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_869
timestamp 1636968456
transform 1 0 81052 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_881
timestamp 1636968456
transform 1 0 82156 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_893
timestamp 1636968456
transform 1 0 83260 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_905
timestamp 1
transform 1 0 84364 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_118_916
timestamp 1
transform 1 0 85376 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_118_925
timestamp 1
transform 1 0 86204 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_933
timestamp 1
transform 1 0 86940 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_969
timestamp 1
transform 1 0 90252 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_977
timestamp 1
transform 1 0 90988 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_118_981
timestamp 1
transform 1 0 91356 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_987
timestamp 1
transform 1 0 91908 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_997
timestamp 1636968456
transform 1 0 92828 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_1009
timestamp 1
transform 1 0 93932 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1013
timestamp 1
transform 1 0 94300 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_1016
timestamp 1
transform 1 0 94576 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1020
timestamp 1
transform 1 0 94944 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1023
timestamp 1
transform 1 0 95220 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1035
timestamp 1
transform 1 0 96324 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1037
timestamp 1
transform 1 0 96508 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_118_1050
timestamp 1
transform 1 0 97704 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1086
timestamp 1
transform 1 0 101016 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_118_1099
timestamp 1
transform 1 0 102212 0 1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1128
timestamp 1636968456
transform 1 0 104880 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_1140
timestamp 1
transform 1 0 105984 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1149
timestamp 1636968456
transform 1 0 106812 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1161
timestamp 1
transform 1 0 107916 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1167
timestamp 1
transform 1 0 108468 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636968456
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636968456
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1636968456
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_39
timestamp 1636968456
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1636968456
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_69
timestamp 1636968456
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_81
timestamp 1636968456
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_93
timestamp 1636968456
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1636968456
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1636968456
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1636968456
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1636968456
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_169
timestamp 1636968456
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_181
timestamp 1636968456
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_193
timestamp 1636968456
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_205
timestamp 1636968456
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_225
timestamp 1636968456
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_237
timestamp 1636968456
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_249
timestamp 1636968456
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_261
timestamp 1636968456
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_281
timestamp 1636968456
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_293
timestamp 1636968456
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_305
timestamp 1636968456
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_317
timestamp 1636968456
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_337
timestamp 1636968456
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_349
timestamp 1636968456
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_361
timestamp 1636968456
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_373
timestamp 1636968456
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_393
timestamp 1636968456
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_405
timestamp 1636968456
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_417
timestamp 1636968456
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_429
timestamp 1636968456
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_449
timestamp 1636968456
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_461
timestamp 1636968456
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_473
timestamp 1636968456
transform 1 0 44620 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_485
timestamp 1636968456
transform 1 0 45724 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1
transform 1 0 46828 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_505
timestamp 1636968456
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_517
timestamp 1636968456
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_529
timestamp 1636968456
transform 1 0 49772 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_541
timestamp 1636968456
transform 1 0 50876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1
transform 1 0 51980 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_561
timestamp 1636968456
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_573
timestamp 1636968456
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_585
timestamp 1636968456
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_597
timestamp 1636968456
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_617
timestamp 1636968456
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_629
timestamp 1636968456
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_641
timestamp 1636968456
transform 1 0 60076 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_653
timestamp 1636968456
transform 1 0 61180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_665
timestamp 1
transform 1 0 62284 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1
transform 1 0 62836 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_673
timestamp 1636968456
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_685
timestamp 1636968456
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_697
timestamp 1636968456
transform 1 0 65228 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_709
timestamp 1636968456
transform 1 0 66332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_721
timestamp 1
transform 1 0 67436 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1
transform 1 0 67988 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_729
timestamp 1636968456
transform 1 0 68172 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_741
timestamp 1636968456
transform 1 0 69276 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_753
timestamp 1636968456
transform 1 0 70380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_765
timestamp 1636968456
transform 1 0 71484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_777
timestamp 1
transform 1 0 72588 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_783
timestamp 1
transform 1 0 73140 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_785
timestamp 1636968456
transform 1 0 73324 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_797
timestamp 1636968456
transform 1 0 74428 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_809
timestamp 1636968456
transform 1 0 75532 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_821
timestamp 1636968456
transform 1 0 76636 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_833
timestamp 1
transform 1 0 77740 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_839
timestamp 1
transform 1 0 78292 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_841
timestamp 1636968456
transform 1 0 78476 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_853
timestamp 1636968456
transform 1 0 79580 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_865
timestamp 1636968456
transform 1 0 80684 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_877
timestamp 1636968456
transform 1 0 81788 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_889
timestamp 1
transform 1 0 82892 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_895
timestamp 1
transform 1 0 83444 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_897
timestamp 1636968456
transform 1 0 83628 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_909
timestamp 1636968456
transform 1 0 84732 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_921
timestamp 1
transform 1 0 85836 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_929
timestamp 1
transform 1 0 86572 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_935
timestamp 1636968456
transform 1 0 87124 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_947
timestamp 1
transform 1 0 88228 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_951
timestamp 1
transform 1 0 88596 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_119_953
timestamp 1
transform 1 0 88780 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_119_958
timestamp 1
transform 1 0 89240 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_119_966
timestamp 1
transform 1 0 89976 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_119_972
timestamp 1
transform 1 0 90528 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_982
timestamp 1636968456
transform 1 0 91448 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_994
timestamp 1
transform 1 0 92552 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1009
timestamp 1636968456
transform 1 0 93932 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_1021
timestamp 1
transform 1 0 95036 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1032
timestamp 1
transform 1 0 96048 0 -1 67456
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1047
timestamp 1636968456
transform 1 0 97428 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_1059
timestamp 1
transform 1 0 98532 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1063
timestamp 1
transform 1 0 98900 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_1065
timestamp 1
transform 1 0 99084 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_1086
timestamp 1
transform 1 0 101016 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1090
timestamp 1
transform 1 0 101384 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_119_1099
timestamp 1
transform 1 0 102212 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_119_1118
timestamp 1
transform 1 0 103960 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1121
timestamp 1636968456
transform 1 0 104236 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1133
timestamp 1636968456
transform 1 0 105340 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1145
timestamp 1636968456
transform 1 0 106444 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_1157
timestamp 1
transform 1 0 107548 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_1165
timestamp 1
transform 1 0 108284 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1636968456
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1636968456
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636968456
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1636968456
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1636968456
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_65
timestamp 1636968456
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1636968456
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1636968456
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_109
timestamp 1636968456
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_121
timestamp 1636968456
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1636968456
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_153
timestamp 1636968456
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_165
timestamp 1636968456
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_177
timestamp 1636968456
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_197
timestamp 1636968456
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_209
timestamp 1636968456
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_221
timestamp 1636968456
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_233
timestamp 1636968456
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_253
timestamp 1636968456
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_265
timestamp 1636968456
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_277
timestamp 1636968456
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_289
timestamp 1636968456
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_309
timestamp 1636968456
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_321
timestamp 1636968456
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_333
timestamp 1636968456
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_345
timestamp 1636968456
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_365
timestamp 1636968456
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_377
timestamp 1636968456
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_389
timestamp 1636968456
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_401
timestamp 1636968456
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_421
timestamp 1636968456
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_433
timestamp 1636968456
transform 1 0 40940 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_445
timestamp 1636968456
transform 1 0 42044 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_457
timestamp 1636968456
transform 1 0 43148 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1
transform 1 0 44252 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1
transform 1 0 44804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_477
timestamp 1636968456
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_489
timestamp 1636968456
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_501
timestamp 1636968456
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_513
timestamp 1636968456
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_533
timestamp 1636968456
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_545
timestamp 1636968456
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_557
timestamp 1636968456
transform 1 0 52348 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_569
timestamp 1636968456
transform 1 0 53452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1
transform 1 0 54556 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1
transform 1 0 55108 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_589
timestamp 1636968456
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_601
timestamp 1636968456
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_613
timestamp 1636968456
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_625
timestamp 1636968456
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_645
timestamp 1636968456
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_657
timestamp 1636968456
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_669
timestamp 1636968456
transform 1 0 62652 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_681
timestamp 1636968456
transform 1 0 63756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1
transform 1 0 64860 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_701
timestamp 1636968456
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_713
timestamp 1636968456
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_725
timestamp 1636968456
transform 1 0 67804 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_737
timestamp 1636968456
transform 1 0 68908 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_749
timestamp 1
transform 1 0 70012 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_755
timestamp 1
transform 1 0 70564 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_757
timestamp 1636968456
transform 1 0 70748 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_769
timestamp 1636968456
transform 1 0 71852 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_781
timestamp 1636968456
transform 1 0 72956 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_793
timestamp 1636968456
transform 1 0 74060 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_805
timestamp 1
transform 1 0 75164 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_811
timestamp 1
transform 1 0 75716 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_813
timestamp 1636968456
transform 1 0 75900 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_825
timestamp 1636968456
transform 1 0 77004 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_837
timestamp 1636968456
transform 1 0 78108 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_849
timestamp 1636968456
transform 1 0 79212 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_861
timestamp 1
transform 1 0 80316 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_867
timestamp 1
transform 1 0 80868 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_869
timestamp 1636968456
transform 1 0 81052 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_881
timestamp 1
transform 1 0 82156 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_887
timestamp 1
transform 1 0 82708 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_912
timestamp 1636968456
transform 1 0 85008 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_925
timestamp 1
transform 1 0 86204 0 1 67456
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_120_966
timestamp 1636968456
transform 1 0 89976 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_120_978
timestamp 1
transform 1 0 91080 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_981
timestamp 1636968456
transform 1 0 91356 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_993
timestamp 1636968456
transform 1 0 92460 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_1005
timestamp 1
transform 1 0 93564 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_120_1013
timestamp 1
transform 1 0 94300 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_1032
timestamp 1
transform 1 0 96048 0 1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1037
timestamp 1636968456
transform 1 0 96508 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_1049
timestamp 1
transform 1 0 97612 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_1065
timestamp 1
transform 1 0 99084 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1069
timestamp 1
transform 1 0 99452 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1079
timestamp 1
transform 1 0 100372 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_120_1090
timestamp 1
transform 1 0 101384 0 1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1111
timestamp 1636968456
transform 1 0 103316 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1123
timestamp 1636968456
transform 1 0 104420 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1135
timestamp 1636968456
transform 1 0 105524 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1147
timestamp 1
transform 1 0 106628 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1149
timestamp 1636968456
transform 1 0 106812 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636968456
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636968456
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1636968456
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_39
timestamp 1636968456
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1636968456
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_69
timestamp 1636968456
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_81
timestamp 1636968456
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_93
timestamp 1636968456
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_113
timestamp 1636968456
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_125
timestamp 1636968456
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_137
timestamp 1636968456
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_149
timestamp 1636968456
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_169
timestamp 1636968456
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_181
timestamp 1636968456
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_193
timestamp 1636968456
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_205
timestamp 1636968456
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_225
timestamp 1636968456
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_237
timestamp 1636968456
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_249
timestamp 1636968456
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_261
timestamp 1636968456
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_281
timestamp 1636968456
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_293
timestamp 1636968456
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_305
timestamp 1636968456
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_317
timestamp 1636968456
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_337
timestamp 1636968456
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_349
timestamp 1636968456
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_361
timestamp 1636968456
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_373
timestamp 1636968456
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_393
timestamp 1636968456
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_405
timestamp 1
transform 1 0 38364 0 -1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_121_426
timestamp 1636968456
transform 1 0 40296 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_438
timestamp 1
transform 1 0 41400 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_121_446
timestamp 1
transform 1 0 42136 0 -1 68544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_121_449
timestamp 1636968456
transform 1 0 42412 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_461
timestamp 1636968456
transform 1 0 43516 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_473
timestamp 1636968456
transform 1 0 44620 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_485
timestamp 1636968456
transform 1 0 45724 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1
transform 1 0 46828 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1
transform 1 0 47380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_505
timestamp 1636968456
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_517
timestamp 1636968456
transform 1 0 48668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_529
timestamp 1636968456
transform 1 0 49772 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_541
timestamp 1636968456
transform 1 0 50876 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_553
timestamp 1
transform 1 0 51980 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_559
timestamp 1
transform 1 0 52532 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_561
timestamp 1636968456
transform 1 0 52716 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_573
timestamp 1636968456
transform 1 0 53820 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_585
timestamp 1636968456
transform 1 0 54924 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_597
timestamp 1636968456
transform 1 0 56028 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_609
timestamp 1
transform 1 0 57132 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1
transform 1 0 57684 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_617
timestamp 1636968456
transform 1 0 57868 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_629
timestamp 1636968456
transform 1 0 58972 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_641
timestamp 1636968456
transform 1 0 60076 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_653
timestamp 1636968456
transform 1 0 61180 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_665
timestamp 1
transform 1 0 62284 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_671
timestamp 1
transform 1 0 62836 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_673
timestamp 1636968456
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_685
timestamp 1636968456
transform 1 0 64124 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_697
timestamp 1636968456
transform 1 0 65228 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_709
timestamp 1636968456
transform 1 0 66332 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_729
timestamp 1636968456
transform 1 0 68172 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_741
timestamp 1636968456
transform 1 0 69276 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_753
timestamp 1636968456
transform 1 0 70380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_765
timestamp 1636968456
transform 1 0 71484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_777
timestamp 1
transform 1 0 72588 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_783
timestamp 1
transform 1 0 73140 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_785
timestamp 1636968456
transform 1 0 73324 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_797
timestamp 1636968456
transform 1 0 74428 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_809
timestamp 1636968456
transform 1 0 75532 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_821
timestamp 1636968456
transform 1 0 76636 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_833
timestamp 1
transform 1 0 77740 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_839
timestamp 1
transform 1 0 78292 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_841
timestamp 1636968456
transform 1 0 78476 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_853
timestamp 1636968456
transform 1 0 79580 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_865
timestamp 1636968456
transform 1 0 80684 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_877
timestamp 1636968456
transform 1 0 81788 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_889
timestamp 1
transform 1 0 82892 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_895
timestamp 1
transform 1 0 83444 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_897
timestamp 1636968456
transform 1 0 83628 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_909
timestamp 1636968456
transform 1 0 84732 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_921
timestamp 1636968456
transform 1 0 85836 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_933
timestamp 1636968456
transform 1 0 86940 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_945
timestamp 1
transform 1 0 88044 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_951
timestamp 1
transform 1 0 88596 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_953
timestamp 1636968456
transform 1 0 88780 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_965
timestamp 1636968456
transform 1 0 89884 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_977
timestamp 1
transform 1 0 90988 0 -1 68544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_121_988
timestamp 1636968456
transform 1 0 92000 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_1000
timestamp 1
transform 1 0 93104 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_121_1009
timestamp 1
transform 1 0 93932 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_121_1017
timestamp 1
transform 1 0 94668 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_121_1026
timestamp 1
transform 1 0 95496 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1032
timestamp 1
transform 1 0 96048 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_121_1045
timestamp 1
transform 1 0 97244 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_121_1056
timestamp 1
transform 1 0 98256 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_121_1099
timestamp 1
transform 1 0 102212 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_121_1113
timestamp 1
transform 1 0 103500 0 -1 68544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1132
timestamp 1636968456
transform 1 0 105248 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1144
timestamp 1636968456
transform 1 0 106352 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1156
timestamp 1636968456
transform 1 0 107456 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1636968456
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1636968456
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636968456
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1636968456
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1636968456
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_65
timestamp 1636968456
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_85
timestamp 1636968456
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_97
timestamp 1636968456
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_109
timestamp 1636968456
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_121
timestamp 1636968456
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_141
timestamp 1636968456
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_153
timestamp 1636968456
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_165
timestamp 1636968456
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_177
timestamp 1636968456
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_197
timestamp 1636968456
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_209
timestamp 1636968456
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_221
timestamp 1636968456
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_233
timestamp 1636968456
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_253
timestamp 1636968456
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_265
timestamp 1636968456
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_277
timestamp 1636968456
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_289
timestamp 1636968456
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_309
timestamp 1636968456
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_321
timestamp 1636968456
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_333
timestamp 1636968456
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_345
timestamp 1636968456
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_365
timestamp 1636968456
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_377
timestamp 1636968456
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_389
timestamp 1636968456
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_401
timestamp 1636968456
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_421
timestamp 1636968456
transform 1 0 39836 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_433
timestamp 1636968456
transform 1 0 40940 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_445
timestamp 1
transform 1 0 42044 0 1 68544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_122_451
timestamp 1636968456
transform 1 0 42596 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_463
timestamp 1
transform 1 0 43700 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_471
timestamp 1
transform 1 0 44436 0 1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_122_495
timestamp 1636968456
transform 1 0 46644 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_507
timestamp 1636968456
transform 1 0 47748 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_519
timestamp 1636968456
transform 1 0 48852 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_531
timestamp 1
transform 1 0 49956 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_533
timestamp 1636968456
transform 1 0 50140 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_545
timestamp 1636968456
transform 1 0 51244 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_557
timestamp 1636968456
transform 1 0 52348 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_569
timestamp 1636968456
transform 1 0 53452 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_581
timestamp 1
transform 1 0 54556 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1
transform 1 0 55108 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_589
timestamp 1636968456
transform 1 0 55292 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_601
timestamp 1636968456
transform 1 0 56396 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_613
timestamp 1
transform 1 0 57500 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_621
timestamp 1
transform 1 0 58236 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_645
timestamp 1
transform 1 0 60444 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_653
timestamp 1
transform 1 0 61180 0 1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_122_658
timestamp 1636968456
transform 1 0 61640 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_670
timestamp 1636968456
transform 1 0 62744 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_682
timestamp 1636968456
transform 1 0 63848 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_694
timestamp 1
transform 1 0 64952 0 1 68544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_122_721
timestamp 1636968456
transform 1 0 67436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_733
timestamp 1636968456
transform 1 0 68540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_745
timestamp 1
transform 1 0 69644 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_753
timestamp 1
transform 1 0 70380 0 1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_122_757
timestamp 1636968456
transform 1 0 70748 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_769
timestamp 1636968456
transform 1 0 71852 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_781
timestamp 1636968456
transform 1 0 72956 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_793
timestamp 1636968456
transform 1 0 74060 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_805
timestamp 1
transform 1 0 75164 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_811
timestamp 1
transform 1 0 75716 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_813
timestamp 1636968456
transform 1 0 75900 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_825
timestamp 1636968456
transform 1 0 77004 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_837
timestamp 1636968456
transform 1 0 78108 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_849
timestamp 1636968456
transform 1 0 79212 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_861
timestamp 1
transform 1 0 80316 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_867
timestamp 1
transform 1 0 80868 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_869
timestamp 1636968456
transform 1 0 81052 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_881
timestamp 1636968456
transform 1 0 82156 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_893
timestamp 1636968456
transform 1 0 83260 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_905
timestamp 1636968456
transform 1 0 84364 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_917
timestamp 1
transform 1 0 85468 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_923
timestamp 1
transform 1 0 86020 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_925
timestamp 1
transform 1 0 86204 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_929
timestamp 1
transform 1 0 86572 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_935
timestamp 1636968456
transform 1 0 87124 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_947
timestamp 1636968456
transform 1 0 88228 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_959
timestamp 1
transform 1 0 89332 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_963
timestamp 1
transform 1 0 89700 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_969
timestamp 1
transform 1 0 90252 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_977
timestamp 1
transform 1 0 90988 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_1006
timestamp 1
transform 1 0 93656 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_1023
timestamp 1
transform 1 0 95220 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_122_1033
timestamp 1
transform 1 0 96140 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_1037
timestamp 1
transform 1 0 96508 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1048
timestamp 1
transform 1 0 97520 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1054
timestamp 1
transform 1 0 98072 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_1058
timestamp 1
transform 1 0 98440 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_1066
timestamp 1
transform 1 0 99176 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_122_1076
timestamp 1
transform 1 0 100096 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_1088
timestamp 1
transform 1 0 101200 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1102
timestamp 1
transform 1 0 102488 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_122_1119
timestamp 1
transform 1 0 104052 0 1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1135
timestamp 1636968456
transform 1 0 105524 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1147
timestamp 1
transform 1 0 106628 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1149
timestamp 1636968456
transform 1 0 106812 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1161
timestamp 1
transform 1 0 107916 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1167
timestamp 1
transform 1 0 108468 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636968456
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636968456
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636968456
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_39
timestamp 1636968456
transform 1 0 4692 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1
transform 1 0 5796 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1636968456
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_69
timestamp 1636968456
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_81
timestamp 1636968456
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_93
timestamp 1636968456
transform 1 0 9660 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_105
timestamp 1
transform 1 0 10764 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_111
timestamp 1
transform 1 0 11316 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_113
timestamp 1636968456
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_125
timestamp 1636968456
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_137
timestamp 1636968456
transform 1 0 13708 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_149
timestamp 1636968456
transform 1 0 14812 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1
transform 1 0 15916 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_169
timestamp 1636968456
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_181
timestamp 1636968456
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_193
timestamp 1636968456
transform 1 0 18860 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_205
timestamp 1636968456
transform 1 0 19964 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_217
timestamp 1
transform 1 0 21068 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_223
timestamp 1
transform 1 0 21620 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_225
timestamp 1636968456
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_237
timestamp 1636968456
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_249
timestamp 1636968456
transform 1 0 24012 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_261
timestamp 1636968456
transform 1 0 25116 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_273
timestamp 1
transform 1 0 26220 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_279
timestamp 1
transform 1 0 26772 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_281
timestamp 1636968456
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_293
timestamp 1636968456
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_305
timestamp 1636968456
transform 1 0 29164 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_317
timestamp 1636968456
transform 1 0 30268 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_329
timestamp 1
transform 1 0 31372 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_335
timestamp 1
transform 1 0 31924 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_337
timestamp 1636968456
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_349
timestamp 1636968456
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_361
timestamp 1636968456
transform 1 0 34316 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_373
timestamp 1636968456
transform 1 0 35420 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_385
timestamp 1
transform 1 0 36524 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_391
timestamp 1
transform 1 0 37076 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_393
timestamp 1636968456
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_405
timestamp 1636968456
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_417
timestamp 1636968456
transform 1 0 39468 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_429
timestamp 1636968456
transform 1 0 40572 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_441
timestamp 1
transform 1 0 41676 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_445
timestamp 1
transform 1 0 42044 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_465
timestamp 1636968456
transform 1 0 43884 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_477
timestamp 1636968456
transform 1 0 44988 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_489
timestamp 1636968456
transform 1 0 46092 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_501
timestamp 1
transform 1 0 47196 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_505
timestamp 1636968456
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_517
timestamp 1636968456
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_529
timestamp 1636968456
transform 1 0 49772 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_541
timestamp 1636968456
transform 1 0 50876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_553
timestamp 1
transform 1 0 51980 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_559
timestamp 1
transform 1 0 52532 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_561
timestamp 1636968456
transform 1 0 52716 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_573
timestamp 1636968456
transform 1 0 53820 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_585
timestamp 1636968456
transform 1 0 54924 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_597
timestamp 1636968456
transform 1 0 56028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_609
timestamp 1
transform 1 0 57132 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_615
timestamp 1
transform 1 0 57684 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_617
timestamp 1636968456
transform 1 0 57868 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_629
timestamp 1636968456
transform 1 0 58972 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_641
timestamp 1636968456
transform 1 0 60076 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_653
timestamp 1
transform 1 0 61180 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_675
timestamp 1636968456
transform 1 0 63204 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_687
timestamp 1636968456
transform 1 0 64308 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_699
timestamp 1
transform 1 0 65412 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_707
timestamp 1
transform 1 0 66148 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_731
timestamp 1636968456
transform 1 0 68356 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_743
timestamp 1636968456
transform 1 0 69460 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_755
timestamp 1636968456
transform 1 0 70564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_767
timestamp 1636968456
transform 1 0 71668 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_779
timestamp 1
transform 1 0 72772 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_783
timestamp 1
transform 1 0 73140 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_785
timestamp 1636968456
transform 1 0 73324 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_797
timestamp 1636968456
transform 1 0 74428 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_809
timestamp 1636968456
transform 1 0 75532 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_821
timestamp 1636968456
transform 1 0 76636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_833
timestamp 1
transform 1 0 77740 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_839
timestamp 1
transform 1 0 78292 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_841
timestamp 1
transform 1 0 78476 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_849
timestamp 1
transform 1 0 79212 0 -1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_854
timestamp 1636968456
transform 1 0 79672 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_866
timestamp 1636968456
transform 1 0 80776 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_878
timestamp 1636968456
transform 1 0 81880 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_890
timestamp 1
transform 1 0 82984 0 -1 69632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_123_897
timestamp 1636968456
transform 1 0 83628 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_909
timestamp 1636968456
transform 1 0 84732 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_921
timestamp 1636968456
transform 1 0 85836 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_933
timestamp 1636968456
transform 1 0 86940 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_945
timestamp 1
transform 1 0 88044 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_951
timestamp 1
transform 1 0 88596 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_123_963
timestamp 1
transform 1 0 89700 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_999
timestamp 1
transform 1 0 93012 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1007
timestamp 1
transform 1 0 93748 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1009
timestamp 1636968456
transform 1 0 93932 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1021
timestamp 1636968456
transform 1 0 95036 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1033
timestamp 1636968456
transform 1 0 96140 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1045
timestamp 1
transform 1 0 97244 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1068
timestamp 1
transform 1 0 99360 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_123_1075
timestamp 1
transform 1 0 100004 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1081
timestamp 1636968456
transform 1 0 100556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_1096
timestamp 1
transform 1 0 101936 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1100
timestamp 1
transform 1 0 102304 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1108
timestamp 1
transform 1 0 103040 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1119
timestamp 1
transform 1 0 104052 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_1121
timestamp 1
transform 1 0 104236 0 -1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1130
timestamp 1636968456
transform 1 0 105064 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1142
timestamp 1636968456
transform 1 0 106168 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1154
timestamp 1636968456
transform 1 0 107272 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_1166
timestamp 1
transform 1 0 108376 0 -1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636968456
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636968456
transform 1 0 2484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 1
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1636968456
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_41
timestamp 1636968456
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_53
timestamp 1636968456
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_65
timestamp 1636968456
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_85
timestamp 1636968456
transform 1 0 8924 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_97
timestamp 1636968456
transform 1 0 10028 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_109
timestamp 1636968456
transform 1 0 11132 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_121
timestamp 1636968456
transform 1 0 12236 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_133
timestamp 1
transform 1 0 13340 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_139
timestamp 1
transform 1 0 13892 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_141
timestamp 1636968456
transform 1 0 14076 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_153
timestamp 1636968456
transform 1 0 15180 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_165
timestamp 1636968456
transform 1 0 16284 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_177
timestamp 1636968456
transform 1 0 17388 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_189
timestamp 1
transform 1 0 18492 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_195
timestamp 1
transform 1 0 19044 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_197
timestamp 1636968456
transform 1 0 19228 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_209
timestamp 1636968456
transform 1 0 20332 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_221
timestamp 1636968456
transform 1 0 21436 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_233
timestamp 1636968456
transform 1 0 22540 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_245
timestamp 1
transform 1 0 23644 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_251
timestamp 1
transform 1 0 24196 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_253
timestamp 1636968456
transform 1 0 24380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_265
timestamp 1636968456
transform 1 0 25484 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_277
timestamp 1636968456
transform 1 0 26588 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_289
timestamp 1636968456
transform 1 0 27692 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_301
timestamp 1
transform 1 0 28796 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_307
timestamp 1
transform 1 0 29348 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_309
timestamp 1
transform 1 0 29532 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_124_317
timestamp 1
transform 1 0 30268 0 1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_124_322
timestamp 1636968456
transform 1 0 30728 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_124_334
timestamp 1
transform 1 0 31832 0 1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_124_340
timestamp 1636968456
transform 1 0 32384 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_352
timestamp 1636968456
transform 1 0 33488 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_365
timestamp 1
transform 1 0 34684 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_373
timestamp 1
transform 1 0 35420 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_392
timestamp 1636968456
transform 1 0 37168 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_404
timestamp 1636968456
transform 1 0 38272 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_416
timestamp 1
transform 1 0 39376 0 1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_124_421
timestamp 1636968456
transform 1 0 39836 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_433
timestamp 1636968456
transform 1 0 40940 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_445
timestamp 1636968456
transform 1 0 42044 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_457
timestamp 1636968456
transform 1 0 43148 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_469
timestamp 1
transform 1 0 44252 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_475
timestamp 1
transform 1 0 44804 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_477
timestamp 1636968456
transform 1 0 44988 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_489
timestamp 1636968456
transform 1 0 46092 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_501
timestamp 1636968456
transform 1 0 47196 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_513
timestamp 1636968456
transform 1 0 48300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_525
timestamp 1
transform 1 0 49404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_531
timestamp 1
transform 1 0 49956 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_533
timestamp 1636968456
transform 1 0 50140 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_545
timestamp 1636968456
transform 1 0 51244 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_557
timestamp 1636968456
transform 1 0 52348 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_569
timestamp 1636968456
transform 1 0 53452 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_581
timestamp 1
transform 1 0 54556 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_587
timestamp 1
transform 1 0 55108 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_589
timestamp 1636968456
transform 1 0 55292 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_601
timestamp 1636968456
transform 1 0 56396 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_613
timestamp 1636968456
transform 1 0 57500 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_625
timestamp 1636968456
transform 1 0 58604 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_637
timestamp 1
transform 1 0 59708 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_643
timestamp 1
transform 1 0 60260 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_645
timestamp 1636968456
transform 1 0 60444 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_657
timestamp 1636968456
transform 1 0 61548 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_669
timestamp 1636968456
transform 1 0 62652 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_681
timestamp 1636968456
transform 1 0 63756 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_693
timestamp 1
transform 1 0 64860 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_699
timestamp 1
transform 1 0 65412 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_701
timestamp 1
transform 1 0 65596 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_124_709
timestamp 1
transform 1 0 66332 0 1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_124_714
timestamp 1636968456
transform 1 0 66792 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_726
timestamp 1636968456
transform 1 0 67896 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_738
timestamp 1636968456
transform 1 0 69000 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_750
timestamp 1
transform 1 0 70104 0 1 69632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_124_757
timestamp 1636968456
transform 1 0 70748 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_769
timestamp 1636968456
transform 1 0 71852 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_781
timestamp 1
transform 1 0 72956 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_124_805
timestamp 1
transform 1 0 75164 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_811
timestamp 1
transform 1 0 75716 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_813
timestamp 1636968456
transform 1 0 75900 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_825
timestamp 1
transform 1 0 77004 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_124_849
timestamp 1
transform 1 0 79212 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_871
timestamp 1636968456
transform 1 0 81236 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_883
timestamp 1636968456
transform 1 0 82340 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_895
timestamp 1636968456
transform 1 0 83444 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_907
timestamp 1636968456
transform 1 0 84548 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_919
timestamp 1
transform 1 0 85652 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_124_923
timestamp 1
transform 1 0 86020 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_925
timestamp 1636968456
transform 1 0 86204 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_937
timestamp 1636968456
transform 1 0 87308 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_949
timestamp 1636968456
transform 1 0 88412 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_979
timestamp 1
transform 1 0 91172 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_985
timestamp 1636968456
transform 1 0 91724 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_997
timestamp 1636968456
transform 1 0 92828 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1009
timestamp 1
transform 1 0 93932 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1015
timestamp 1
transform 1 0 94484 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1025
timestamp 1
transform 1 0 95404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1031
timestamp 1
transform 1 0 95956 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1044
timestamp 1
transform 1 0 97152 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_124_1053
timestamp 1
transform 1 0 97980 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1057
timestamp 1
transform 1 0 98348 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_124_1061
timestamp 1
transform 1 0 98716 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_124_1068
timestamp 1
transform 1 0 99360 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1088
timestamp 1
transform 1 0 101200 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1100
timestamp 1636968456
transform 1 0 102304 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1112
timestamp 1
transform 1 0 103408 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1118
timestamp 1
transform 1 0 103960 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1134
timestamp 1636968456
transform 1 0 105432 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_124_1146
timestamp 1
transform 1 0 106536 0 1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1149
timestamp 1636968456
transform 1 0 106812 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_124_1161
timestamp 1
transform 1 0 107916 0 1 69632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_125_3
timestamp 1636968456
transform 1 0 1380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_15
timestamp 1636968456
transform 1 0 2484 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_27
timestamp 1636968456
transform 1 0 3588 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_39
timestamp 1636968456
transform 1 0 4692 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1
transform 1 0 5796 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1636968456
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_69
timestamp 1636968456
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_81
timestamp 1636968456
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_93
timestamp 1636968456
transform 1 0 9660 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1
transform 1 0 10764 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1
transform 1 0 11316 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_113
timestamp 1636968456
transform 1 0 11500 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_125
timestamp 1636968456
transform 1 0 12604 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_137
timestamp 1636968456
transform 1 0 13708 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_149
timestamp 1636968456
transform 1 0 14812 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_161
timestamp 1
transform 1 0 15916 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_167
timestamp 1
transform 1 0 16468 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_169
timestamp 1636968456
transform 1 0 16652 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_181
timestamp 1636968456
transform 1 0 17756 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_193
timestamp 1636968456
transform 1 0 18860 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_205
timestamp 1636968456
transform 1 0 19964 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_217
timestamp 1
transform 1 0 21068 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_223
timestamp 1
transform 1 0 21620 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_225
timestamp 1636968456
transform 1 0 21804 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_237
timestamp 1636968456
transform 1 0 22908 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_249
timestamp 1636968456
transform 1 0 24012 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_261
timestamp 1636968456
transform 1 0 25116 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_273
timestamp 1
transform 1 0 26220 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_279
timestamp 1
transform 1 0 26772 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_281
timestamp 1636968456
transform 1 0 26956 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_293
timestamp 1636968456
transform 1 0 28060 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_305
timestamp 1636968456
transform 1 0 29164 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_125_317
timestamp 1
transform 1 0 30268 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_125_353
timestamp 1
transform 1 0 33580 0 -1 70720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_125_379
timestamp 1636968456
transform 1 0 35972 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_391
timestamp 1
transform 1 0 37076 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_393
timestamp 1636968456
transform 1 0 37260 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_405
timestamp 1636968456
transform 1 0 38364 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_417
timestamp 1636968456
transform 1 0 39468 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_429
timestamp 1636968456
transform 1 0 40572 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_441
timestamp 1
transform 1 0 41676 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_447
timestamp 1
transform 1 0 42228 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_449
timestamp 1636968456
transform 1 0 42412 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_461
timestamp 1636968456
transform 1 0 43516 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_473
timestamp 1636968456
transform 1 0 44620 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_485
timestamp 1636968456
transform 1 0 45724 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_497
timestamp 1
transform 1 0 46828 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_503
timestamp 1
transform 1 0 47380 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_505
timestamp 1636968456
transform 1 0 47564 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_517
timestamp 1636968456
transform 1 0 48668 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_529
timestamp 1636968456
transform 1 0 49772 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_541
timestamp 1636968456
transform 1 0 50876 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_553
timestamp 1
transform 1 0 51980 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_559
timestamp 1
transform 1 0 52532 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_561
timestamp 1636968456
transform 1 0 52716 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_573
timestamp 1636968456
transform 1 0 53820 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_585
timestamp 1636968456
transform 1 0 54924 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_597
timestamp 1636968456
transform 1 0 56028 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_609
timestamp 1
transform 1 0 57132 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_615
timestamp 1
transform 1 0 57684 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_617
timestamp 1636968456
transform 1 0 57868 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_629
timestamp 1636968456
transform 1 0 58972 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_641
timestamp 1636968456
transform 1 0 60076 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_653
timestamp 1636968456
transform 1 0 61180 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_665
timestamp 1
transform 1 0 62284 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_671
timestamp 1
transform 1 0 62836 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_673
timestamp 1636968456
transform 1 0 63020 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_685
timestamp 1636968456
transform 1 0 64124 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_697
timestamp 1636968456
transform 1 0 65228 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_709
timestamp 1636968456
transform 1 0 66332 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_721
timestamp 1
transform 1 0 67436 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_727
timestamp 1
transform 1 0 67988 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_729
timestamp 1636968456
transform 1 0 68172 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_741
timestamp 1636968456
transform 1 0 69276 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_753
timestamp 1636968456
transform 1 0 70380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_765
timestamp 1636968456
transform 1 0 71484 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_777
timestamp 1
transform 1 0 72588 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_783
timestamp 1
transform 1 0 73140 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_785
timestamp 1636968456
transform 1 0 73324 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_797
timestamp 1636968456
transform 1 0 74428 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_809
timestamp 1636968456
transform 1 0 75532 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_821
timestamp 1636968456
transform 1 0 76636 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_833
timestamp 1
transform 1 0 77740 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_839
timestamp 1
transform 1 0 78292 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_841
timestamp 1636968456
transform 1 0 78476 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_853
timestamp 1636968456
transform 1 0 79580 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_865
timestamp 1636968456
transform 1 0 80684 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_877
timestamp 1636968456
transform 1 0 81788 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_889
timestamp 1
transform 1 0 82892 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_895
timestamp 1
transform 1 0 83444 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_897
timestamp 1636968456
transform 1 0 83628 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_909
timestamp 1636968456
transform 1 0 84732 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_921
timestamp 1636968456
transform 1 0 85836 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_933
timestamp 1
transform 1 0 86940 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_941
timestamp 1
transform 1 0 87676 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_125_949
timestamp 1
transform 1 0 88412 0 -1 70720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_125_953
timestamp 1636968456
transform 1 0 88780 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_965
timestamp 1
transform 1 0 89884 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_981
timestamp 1636968456
transform 1 0 91356 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_993
timestamp 1
transform 1 0 92460 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_125_1003
timestamp 1
transform 1 0 93380 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1007
timestamp 1
transform 1 0 93748 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1009
timestamp 1636968456
transform 1 0 93932 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_1021
timestamp 1
transform 1 0 95036 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1029
timestamp 1
transform 1 0 95772 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1037
timestamp 1
transform 1 0 96508 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_125_1062
timestamp 1
transform 1 0 98808 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_125_1071
timestamp 1
transform 1 0 99636 0 -1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1078
timestamp 1636968456
transform 1 0 100280 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_1090
timestamp 1
transform 1 0 101384 0 -1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1101
timestamp 1636968456
transform 1 0 102396 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1113
timestamp 1
transform 1 0 103500 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1119
timestamp 1
transform 1 0 104052 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_1121
timestamp 1
transform 1 0 104236 0 -1 70720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1144
timestamp 1636968456
transform 1 0 106352 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1156
timestamp 1
transform 1 0 107456 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1162
timestamp 1
transform 1 0 108008 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636968456
transform 1 0 1380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636968456
transform 1 0 2484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 1
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636968456
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1636968456
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_53
timestamp 1636968456
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_65
timestamp 1636968456
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_85
timestamp 1636968456
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_97
timestamp 1636968456
transform 1 0 10028 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_109
timestamp 1636968456
transform 1 0 11132 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_121
timestamp 1636968456
transform 1 0 12236 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_133
timestamp 1
transform 1 0 13340 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_139
timestamp 1
transform 1 0 13892 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_141
timestamp 1636968456
transform 1 0 14076 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_153
timestamp 1636968456
transform 1 0 15180 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_165
timestamp 1636968456
transform 1 0 16284 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_177
timestamp 1636968456
transform 1 0 17388 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_189
timestamp 1
transform 1 0 18492 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_195
timestamp 1
transform 1 0 19044 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_197
timestamp 1636968456
transform 1 0 19228 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_209
timestamp 1636968456
transform 1 0 20332 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_221
timestamp 1636968456
transform 1 0 21436 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_233
timestamp 1636968456
transform 1 0 22540 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_245
timestamp 1
transform 1 0 23644 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_251
timestamp 1
transform 1 0 24196 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_253
timestamp 1636968456
transform 1 0 24380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_265
timestamp 1636968456
transform 1 0 25484 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_277
timestamp 1636968456
transform 1 0 26588 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_289
timestamp 1636968456
transform 1 0 27692 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_301
timestamp 1
transform 1 0 28796 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_307
timestamp 1
transform 1 0 29348 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_309
timestamp 1636968456
transform 1 0 29532 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_321
timestamp 1
transform 1 0 30636 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_126_325
timestamp 1
transform 1 0 31004 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_350
timestamp 1636968456
transform 1 0 33304 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_126_362
timestamp 1
transform 1 0 34408 0 1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_126_365
timestamp 1636968456
transform 1 0 34684 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_377
timestamp 1636968456
transform 1 0 35788 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_389
timestamp 1636968456
transform 1 0 36892 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_401
timestamp 1636968456
transform 1 0 37996 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_413
timestamp 1
transform 1 0 39100 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_419
timestamp 1
transform 1 0 39652 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_421
timestamp 1636968456
transform 1 0 39836 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_433
timestamp 1636968456
transform 1 0 40940 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_445
timestamp 1636968456
transform 1 0 42044 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_457
timestamp 1636968456
transform 1 0 43148 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_469
timestamp 1
transform 1 0 44252 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_475
timestamp 1
transform 1 0 44804 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_477
timestamp 1636968456
transform 1 0 44988 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_489
timestamp 1636968456
transform 1 0 46092 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_501
timestamp 1
transform 1 0 47196 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_517
timestamp 1636968456
transform 1 0 48668 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_126_529
timestamp 1
transform 1 0 49772 0 1 70720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_126_533
timestamp 1636968456
transform 1 0 50140 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_545
timestamp 1636968456
transform 1 0 51244 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_557
timestamp 1636968456
transform 1 0 52348 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_569
timestamp 1636968456
transform 1 0 53452 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_581
timestamp 1
transform 1 0 54556 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_587
timestamp 1
transform 1 0 55108 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_589
timestamp 1636968456
transform 1 0 55292 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_601
timestamp 1636968456
transform 1 0 56396 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_613
timestamp 1636968456
transform 1 0 57500 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_625
timestamp 1636968456
transform 1 0 58604 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_637
timestamp 1
transform 1 0 59708 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_643
timestamp 1
transform 1 0 60260 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_645
timestamp 1636968456
transform 1 0 60444 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_657
timestamp 1636968456
transform 1 0 61548 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_669
timestamp 1636968456
transform 1 0 62652 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_681
timestamp 1636968456
transform 1 0 63756 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_693
timestamp 1
transform 1 0 64860 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_699
timestamp 1
transform 1 0 65412 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_701
timestamp 1636968456
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_713
timestamp 1636968456
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_725
timestamp 1636968456
transform 1 0 67804 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_737
timestamp 1636968456
transform 1 0 68908 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_749
timestamp 1
transform 1 0 70012 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_755
timestamp 1
transform 1 0 70564 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_757
timestamp 1636968456
transform 1 0 70748 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_769
timestamp 1
transform 1 0 71852 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_775
timestamp 1
transform 1 0 72404 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_796
timestamp 1636968456
transform 1 0 74336 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_808
timestamp 1
transform 1 0 75440 0 1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_126_813
timestamp 1636968456
transform 1 0 75900 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_825
timestamp 1636968456
transform 1 0 77004 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_837
timestamp 1636968456
transform 1 0 78108 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_867
timestamp 1
transform 1 0 80868 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_871
timestamp 1636968456
transform 1 0 81236 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_883
timestamp 1636968456
transform 1 0 82340 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_895
timestamp 1636968456
transform 1 0 83444 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_907
timestamp 1
transform 1 0 84548 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_126_915
timestamp 1
transform 1 0 85284 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_126_921
timestamp 1
transform 1 0 85836 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_946
timestamp 1636968456
transform 1 0 88136 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_958
timestamp 1636968456
transform 1 0 89240 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_970
timestamp 1
transform 1 0 90344 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_126_978
timestamp 1
transform 1 0 91080 0 1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_126_981
timestamp 1636968456
transform 1 0 91356 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_993
timestamp 1
transform 1 0 92460 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1016
timestamp 1636968456
transform 1 0 94576 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_1028
timestamp 1
transform 1 0 95680 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1043
timestamp 1
transform 1 0 97060 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_126_1055
timestamp 1
transform 1 0 98164 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_126_1061
timestamp 1
transform 1 0 98716 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_126_1071
timestamp 1
transform 1 0 99636 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_126_1080
timestamp 1
transform 1 0 100464 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1084
timestamp 1
transform 1 0 100832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_126_1093
timestamp 1
transform 1 0 101660 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_126_1104
timestamp 1
transform 1 0 102672 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1108
timestamp 1
transform 1 0 103040 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_126_1125
timestamp 1
transform 1 0 104604 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_126_1145
timestamp 1
transform 1 0 106444 0 1 70720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1149
timestamp 1636968456
transform 1 0 106812 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_126_1161
timestamp 1
transform 1 0 107916 0 1 70720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_127_11
timestamp 1636968456
transform 1 0 2116 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_23
timestamp 1636968456
transform 1 0 3220 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_35
timestamp 1636968456
transform 1 0 4324 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_47
timestamp 1
transform 1 0 5428 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1636968456
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_69
timestamp 1636968456
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_81
timestamp 1636968456
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_93
timestamp 1636968456
transform 1 0 9660 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_105
timestamp 1
transform 1 0 10764 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_111
timestamp 1
transform 1 0 11316 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_113
timestamp 1636968456
transform 1 0 11500 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_125
timestamp 1636968456
transform 1 0 12604 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_137
timestamp 1636968456
transform 1 0 13708 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_149
timestamp 1636968456
transform 1 0 14812 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_161
timestamp 1
transform 1 0 15916 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_167
timestamp 1
transform 1 0 16468 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_169
timestamp 1636968456
transform 1 0 16652 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_181
timestamp 1636968456
transform 1 0 17756 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_193
timestamp 1636968456
transform 1 0 18860 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_205
timestamp 1636968456
transform 1 0 19964 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_217
timestamp 1
transform 1 0 21068 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_223
timestamp 1
transform 1 0 21620 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_225
timestamp 1636968456
transform 1 0 21804 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_237
timestamp 1636968456
transform 1 0 22908 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_249
timestamp 1636968456
transform 1 0 24012 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_261
timestamp 1636968456
transform 1 0 25116 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_273
timestamp 1
transform 1 0 26220 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_279
timestamp 1
transform 1 0 26772 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_281
timestamp 1636968456
transform 1 0 26956 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_293
timestamp 1636968456
transform 1 0 28060 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_305
timestamp 1636968456
transform 1 0 29164 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_317
timestamp 1636968456
transform 1 0 30268 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_329
timestamp 1
transform 1 0 31372 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_335
timestamp 1
transform 1 0 31924 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_337
timestamp 1636968456
transform 1 0 32108 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_349
timestamp 1636968456
transform 1 0 33212 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_361
timestamp 1636968456
transform 1 0 34316 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_373
timestamp 1636968456
transform 1 0 35420 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_385
timestamp 1
transform 1 0 36524 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_391
timestamp 1
transform 1 0 37076 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_393
timestamp 1636968456
transform 1 0 37260 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_405
timestamp 1636968456
transform 1 0 38364 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_417
timestamp 1636968456
transform 1 0 39468 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_429
timestamp 1636968456
transform 1 0 40572 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_441
timestamp 1
transform 1 0 41676 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_447
timestamp 1
transform 1 0 42228 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_449
timestamp 1636968456
transform 1 0 42412 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_461
timestamp 1636968456
transform 1 0 43516 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_473
timestamp 1636968456
transform 1 0 44620 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_485
timestamp 1636968456
transform 1 0 45724 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_497
timestamp 1
transform 1 0 46828 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_503
timestamp 1
transform 1 0 47380 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_505
timestamp 1636968456
transform 1 0 47564 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_517
timestamp 1636968456
transform 1 0 48668 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_529
timestamp 1636968456
transform 1 0 49772 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_541
timestamp 1636968456
transform 1 0 50876 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_553
timestamp 1
transform 1 0 51980 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_559
timestamp 1
transform 1 0 52532 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_561
timestamp 1636968456
transform 1 0 52716 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_573
timestamp 1636968456
transform 1 0 53820 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_585
timestamp 1636968456
transform 1 0 54924 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_597
timestamp 1636968456
transform 1 0 56028 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_609
timestamp 1
transform 1 0 57132 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_615
timestamp 1
transform 1 0 57684 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_617
timestamp 1636968456
transform 1 0 57868 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_629
timestamp 1636968456
transform 1 0 58972 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_641
timestamp 1636968456
transform 1 0 60076 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_653
timestamp 1636968456
transform 1 0 61180 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_665
timestamp 1
transform 1 0 62284 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_671
timestamp 1
transform 1 0 62836 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_673
timestamp 1636968456
transform 1 0 63020 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_685
timestamp 1636968456
transform 1 0 64124 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_697
timestamp 1636968456
transform 1 0 65228 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_709
timestamp 1636968456
transform 1 0 66332 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_721
timestamp 1
transform 1 0 67436 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_727
timestamp 1
transform 1 0 67988 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_729
timestamp 1636968456
transform 1 0 68172 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_741
timestamp 1636968456
transform 1 0 69276 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_753
timestamp 1636968456
transform 1 0 70380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_765
timestamp 1636968456
transform 1 0 71484 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_777
timestamp 1
transform 1 0 72588 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_783
timestamp 1
transform 1 0 73140 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_785
timestamp 1636968456
transform 1 0 73324 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_797
timestamp 1636968456
transform 1 0 74428 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_809
timestamp 1636968456
transform 1 0 75532 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_821
timestamp 1636968456
transform 1 0 76636 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_833
timestamp 1
transform 1 0 77740 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_839
timestamp 1
transform 1 0 78292 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_841
timestamp 1636968456
transform 1 0 78476 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_853
timestamp 1636968456
transform 1 0 79580 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_865
timestamp 1636968456
transform 1 0 80684 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_877
timestamp 1636968456
transform 1 0 81788 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_889
timestamp 1
transform 1 0 82892 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_895
timestamp 1
transform 1 0 83444 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_897
timestamp 1636968456
transform 1 0 83628 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_909
timestamp 1636968456
transform 1 0 84732 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_921
timestamp 1636968456
transform 1 0 85836 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_933
timestamp 1636968456
transform 1 0 86940 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_945
timestamp 1
transform 1 0 88044 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_951
timestamp 1
transform 1 0 88596 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_953
timestamp 1
transform 1 0 88780 0 -1 71808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_127_984
timestamp 1636968456
transform 1 0 91632 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_996
timestamp 1636968456
transform 1 0 92736 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1009
timestamp 1636968456
transform 1 0 93932 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_1021
timestamp 1
transform 1 0 95036 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1027
timestamp 1
transform 1 0 95588 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_127_1034
timestamp 1
transform 1 0 96232 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1040
timestamp 1
transform 1 0 96784 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_1046
timestamp 1
transform 1 0 97336 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1050
timestamp 1
transform 1 0 97704 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_127_1056
timestamp 1
transform 1 0 98256 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_127_1065
timestamp 1
transform 1 0 99084 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_127_1074
timestamp 1
transform 1 0 99912 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_127_1087
timestamp 1
transform 1 0 101108 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_127_1108
timestamp 1
transform 1 0 103040 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1119
timestamp 1
transform 1 0 104052 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_1127
timestamp 1
transform 1 0 104788 0 -1 71808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1140
timestamp 1636968456
transform 1 0 105984 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_1152
timestamp 1
transform 1 0 107088 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1156
timestamp 1
transform 1 0 107456 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1160
timestamp 1
transform 1 0 107824 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636968456
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636968456
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1636968456
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_41
timestamp 1636968456
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_53
timestamp 1636968456
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_65
timestamp 1636968456
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_85
timestamp 1636968456
transform 1 0 8924 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_97
timestamp 1636968456
transform 1 0 10028 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_109
timestamp 1636968456
transform 1 0 11132 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_121
timestamp 1636968456
transform 1 0 12236 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_133
timestamp 1
transform 1 0 13340 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_139
timestamp 1
transform 1 0 13892 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_141
timestamp 1636968456
transform 1 0 14076 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_153
timestamp 1636968456
transform 1 0 15180 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_165
timestamp 1636968456
transform 1 0 16284 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_177
timestamp 1636968456
transform 1 0 17388 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_189
timestamp 1
transform 1 0 18492 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_195
timestamp 1
transform 1 0 19044 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_197
timestamp 1636968456
transform 1 0 19228 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_209
timestamp 1636968456
transform 1 0 20332 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_221
timestamp 1636968456
transform 1 0 21436 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_233
timestamp 1636968456
transform 1 0 22540 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_245
timestamp 1
transform 1 0 23644 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_251
timestamp 1
transform 1 0 24196 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_253
timestamp 1636968456
transform 1 0 24380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_265
timestamp 1636968456
transform 1 0 25484 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_277
timestamp 1636968456
transform 1 0 26588 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_289
timestamp 1636968456
transform 1 0 27692 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_301
timestamp 1
transform 1 0 28796 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_307
timestamp 1
transform 1 0 29348 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_309
timestamp 1636968456
transform 1 0 29532 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_321
timestamp 1636968456
transform 1 0 30636 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_333
timestamp 1636968456
transform 1 0 31740 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_345
timestamp 1636968456
transform 1 0 32844 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_357
timestamp 1
transform 1 0 33948 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_363
timestamp 1
transform 1 0 34500 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_365
timestamp 1636968456
transform 1 0 34684 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_377
timestamp 1636968456
transform 1 0 35788 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_389
timestamp 1636968456
transform 1 0 36892 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_401
timestamp 1636968456
transform 1 0 37996 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_413
timestamp 1
transform 1 0 39100 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_419
timestamp 1
transform 1 0 39652 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_421
timestamp 1636968456
transform 1 0 39836 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_433
timestamp 1636968456
transform 1 0 40940 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_445
timestamp 1636968456
transform 1 0 42044 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_457
timestamp 1636968456
transform 1 0 43148 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_469
timestamp 1
transform 1 0 44252 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_475
timestamp 1
transform 1 0 44804 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_477
timestamp 1636968456
transform 1 0 44988 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_489
timestamp 1636968456
transform 1 0 46092 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_501
timestamp 1636968456
transform 1 0 47196 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_513
timestamp 1636968456
transform 1 0 48300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_525
timestamp 1
transform 1 0 49404 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_531
timestamp 1
transform 1 0 49956 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_533
timestamp 1636968456
transform 1 0 50140 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_545
timestamp 1636968456
transform 1 0 51244 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_557
timestamp 1636968456
transform 1 0 52348 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_569
timestamp 1636968456
transform 1 0 53452 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_581
timestamp 1
transform 1 0 54556 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_587
timestamp 1
transform 1 0 55108 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_589
timestamp 1636968456
transform 1 0 55292 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_601
timestamp 1636968456
transform 1 0 56396 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_613
timestamp 1636968456
transform 1 0 57500 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_625
timestamp 1636968456
transform 1 0 58604 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_637
timestamp 1
transform 1 0 59708 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_643
timestamp 1
transform 1 0 60260 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_645
timestamp 1636968456
transform 1 0 60444 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_657
timestamp 1636968456
transform 1 0 61548 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_669
timestamp 1636968456
transform 1 0 62652 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_681
timestamp 1636968456
transform 1 0 63756 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_693
timestamp 1
transform 1 0 64860 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_699
timestamp 1
transform 1 0 65412 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_701
timestamp 1636968456
transform 1 0 65596 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_713
timestamp 1636968456
transform 1 0 66700 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_725
timestamp 1636968456
transform 1 0 67804 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_737
timestamp 1636968456
transform 1 0 68908 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_749
timestamp 1
transform 1 0 70012 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_755
timestamp 1
transform 1 0 70564 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_757
timestamp 1636968456
transform 1 0 70748 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_769
timestamp 1636968456
transform 1 0 71852 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_781
timestamp 1636968456
transform 1 0 72956 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_793
timestamp 1636968456
transform 1 0 74060 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_805
timestamp 1
transform 1 0 75164 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_811
timestamp 1
transform 1 0 75716 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_813
timestamp 1636968456
transform 1 0 75900 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_825
timestamp 1636968456
transform 1 0 77004 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_837
timestamp 1636968456
transform 1 0 78108 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_849
timestamp 1636968456
transform 1 0 79212 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_861
timestamp 1
transform 1 0 80316 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_867
timestamp 1
transform 1 0 80868 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_869
timestamp 1
transform 1 0 81052 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_128_877
timestamp 1
transform 1 0 81788 0 1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_897
timestamp 1636968456
transform 1 0 83628 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_909
timestamp 1
transform 1 0 84732 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_915
timestamp 1
transform 1 0 85284 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_128_921
timestamp 1
transform 1 0 85836 0 1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_128_925
timestamp 1636968456
transform 1 0 86204 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_937
timestamp 1636968456
transform 1 0 87308 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_954
timestamp 1636968456
transform 1 0 88872 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_966
timestamp 1636968456
transform 1 0 89976 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_128_978
timestamp 1
transform 1 0 91080 0 1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_981
timestamp 1636968456
transform 1 0 91356 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_993
timestamp 1
transform 1 0 92460 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_128_1001
timestamp 1
transform 1 0 93196 0 1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1011
timestamp 1636968456
transform 1 0 94116 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1023
timestamp 1636968456
transform 1 0 95220 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1035
timestamp 1
transform 1 0 96324 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1044
timestamp 1
transform 1 0 97152 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_128_1067
timestamp 1
transform 1 0 99268 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_128_1078
timestamp 1
transform 1 0 100280 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1086
timestamp 1
transform 1 0 101016 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_128_1090
timestamp 1
transform 1 0 101384 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_128_1093
timestamp 1
transform 1 0 101660 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_128_1102
timestamp 1
transform 1 0 102488 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_128_1114
timestamp 1
transform 1 0 103592 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_128_1125
timestamp 1
transform 1 0 104604 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_128_1143
timestamp 1
transform 1 0 106260 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1147
timestamp 1
transform 1 0 106628 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1149
timestamp 1636968456
transform 1 0 106812 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_1161
timestamp 1
transform 1 0 107916 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1167
timestamp 1
transform 1 0 108468 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_9
timestamp 1636968456
transform 1 0 1932 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_21
timestamp 1636968456
transform 1 0 3036 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_33
timestamp 1636968456
transform 1 0 4140 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_45
timestamp 1
transform 1 0 5244 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_129_53
timestamp 1
transform 1 0 5980 0 -1 72896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_129_57
timestamp 1636968456
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_69
timestamp 1636968456
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_81
timestamp 1636968456
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_93
timestamp 1636968456
transform 1 0 9660 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_105
timestamp 1
transform 1 0 10764 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_111
timestamp 1
transform 1 0 11316 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_113
timestamp 1636968456
transform 1 0 11500 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_125
timestamp 1636968456
transform 1 0 12604 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_137
timestamp 1636968456
transform 1 0 13708 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_149
timestamp 1636968456
transform 1 0 14812 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_161
timestamp 1
transform 1 0 15916 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_167
timestamp 1
transform 1 0 16468 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_169
timestamp 1636968456
transform 1 0 16652 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_181
timestamp 1636968456
transform 1 0 17756 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_193
timestamp 1636968456
transform 1 0 18860 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_205
timestamp 1636968456
transform 1 0 19964 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_217
timestamp 1
transform 1 0 21068 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_223
timestamp 1
transform 1 0 21620 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_225
timestamp 1636968456
transform 1 0 21804 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_237
timestamp 1636968456
transform 1 0 22908 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_249
timestamp 1636968456
transform 1 0 24012 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_261
timestamp 1636968456
transform 1 0 25116 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_273
timestamp 1
transform 1 0 26220 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_279
timestamp 1
transform 1 0 26772 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_281
timestamp 1636968456
transform 1 0 26956 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_293
timestamp 1636968456
transform 1 0 28060 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_305
timestamp 1636968456
transform 1 0 29164 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_317
timestamp 1636968456
transform 1 0 30268 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_329
timestamp 1
transform 1 0 31372 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_335
timestamp 1
transform 1 0 31924 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_337
timestamp 1636968456
transform 1 0 32108 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_349
timestamp 1636968456
transform 1 0 33212 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_361
timestamp 1636968456
transform 1 0 34316 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_373
timestamp 1636968456
transform 1 0 35420 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_385
timestamp 1
transform 1 0 36524 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_391
timestamp 1
transform 1 0 37076 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_393
timestamp 1636968456
transform 1 0 37260 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_405
timestamp 1636968456
transform 1 0 38364 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_417
timestamp 1636968456
transform 1 0 39468 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_429
timestamp 1636968456
transform 1 0 40572 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_441
timestamp 1
transform 1 0 41676 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_447
timestamp 1
transform 1 0 42228 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_449
timestamp 1636968456
transform 1 0 42412 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_461
timestamp 1636968456
transform 1 0 43516 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_473
timestamp 1636968456
transform 1 0 44620 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_485
timestamp 1636968456
transform 1 0 45724 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_497
timestamp 1
transform 1 0 46828 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_503
timestamp 1
transform 1 0 47380 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_505
timestamp 1636968456
transform 1 0 47564 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_517
timestamp 1636968456
transform 1 0 48668 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_529
timestamp 1636968456
transform 1 0 49772 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_541
timestamp 1636968456
transform 1 0 50876 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_553
timestamp 1
transform 1 0 51980 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_559
timestamp 1
transform 1 0 52532 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_561
timestamp 1636968456
transform 1 0 52716 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_573
timestamp 1636968456
transform 1 0 53820 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_585
timestamp 1636968456
transform 1 0 54924 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_597
timestamp 1636968456
transform 1 0 56028 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_609
timestamp 1
transform 1 0 57132 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_615
timestamp 1
transform 1 0 57684 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_617
timestamp 1636968456
transform 1 0 57868 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_629
timestamp 1636968456
transform 1 0 58972 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_641
timestamp 1636968456
transform 1 0 60076 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_653
timestamp 1636968456
transform 1 0 61180 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_665
timestamp 1
transform 1 0 62284 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_671
timestamp 1
transform 1 0 62836 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_673
timestamp 1636968456
transform 1 0 63020 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_685
timestamp 1636968456
transform 1 0 64124 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_697
timestamp 1636968456
transform 1 0 65228 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_709
timestamp 1636968456
transform 1 0 66332 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_721
timestamp 1
transform 1 0 67436 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_727
timestamp 1
transform 1 0 67988 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_129_729
timestamp 1
transform 1 0 68172 0 -1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_129_740
timestamp 1636968456
transform 1 0 69184 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_752
timestamp 1636968456
transform 1 0 70288 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_764
timestamp 1636968456
transform 1 0 71392 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_776
timestamp 1
transform 1 0 72496 0 -1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_129_785
timestamp 1636968456
transform 1 0 73324 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_797
timestamp 1636968456
transform 1 0 74428 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_809
timestamp 1636968456
transform 1 0 75532 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_821
timestamp 1636968456
transform 1 0 76636 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_833
timestamp 1
transform 1 0 77740 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_839
timestamp 1
transform 1 0 78292 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_841
timestamp 1636968456
transform 1 0 78476 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_853
timestamp 1636968456
transform 1 0 79580 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_865
timestamp 1636968456
transform 1 0 80684 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_877
timestamp 1636968456
transform 1 0 81788 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_889
timestamp 1
transform 1 0 82892 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_895
timestamp 1
transform 1 0 83444 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_897
timestamp 1636968456
transform 1 0 83628 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_909
timestamp 1636968456
transform 1 0 84732 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_921
timestamp 1
transform 1 0 85836 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_129_949
timestamp 1
transform 1 0 88412 0 -1 72896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_129_953
timestamp 1636968456
transform 1 0 88780 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_965
timestamp 1636968456
transform 1 0 89884 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_977
timestamp 1636968456
transform 1 0 90988 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_989
timestamp 1636968456
transform 1 0 92092 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_1001
timestamp 1
transform 1 0 93196 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1007
timestamp 1
transform 1 0 93748 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1009
timestamp 1636968456
transform 1 0 93932 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1021
timestamp 1636968456
transform 1 0 95036 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1033
timestamp 1
transform 1 0 96140 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_129_1041
timestamp 1
transform 1 0 96876 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_129_1062
timestamp 1
transform 1 0 98808 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_129_1070
timestamp 1
transform 1 0 99544 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1074
timestamp 1
transform 1 0 99912 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_129_1089
timestamp 1
transform 1 0 101292 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_129_1096
timestamp 1
transform 1 0 101936 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1102
timestamp 1
transform 1 0 102488 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_129_1108
timestamp 1
transform 1 0 103040 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1112
timestamp 1
transform 1 0 103408 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1146
timestamp 1636968456
transform 1 0 106536 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_1158
timestamp 1
transform 1 0 107640 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1162
timestamp 1
transform 1 0 108008 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_9
timestamp 1636968456
transform 1 0 1932 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_21
timestamp 1
transform 1 0 3036 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1636968456
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_41
timestamp 1636968456
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_53
timestamp 1636968456
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_65
timestamp 1636968456
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_85
timestamp 1636968456
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_97
timestamp 1636968456
transform 1 0 10028 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_109
timestamp 1636968456
transform 1 0 11132 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_121
timestamp 1636968456
transform 1 0 12236 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_133
timestamp 1
transform 1 0 13340 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_139
timestamp 1
transform 1 0 13892 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_141
timestamp 1636968456
transform 1 0 14076 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_153
timestamp 1636968456
transform 1 0 15180 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_165
timestamp 1636968456
transform 1 0 16284 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_177
timestamp 1636968456
transform 1 0 17388 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_189
timestamp 1
transform 1 0 18492 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_195
timestamp 1
transform 1 0 19044 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_197
timestamp 1636968456
transform 1 0 19228 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_209
timestamp 1636968456
transform 1 0 20332 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_245
timestamp 1
transform 1 0 23644 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_251
timestamp 1
transform 1 0 24196 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_253
timestamp 1636968456
transform 1 0 24380 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_265
timestamp 1636968456
transform 1 0 25484 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_277
timestamp 1636968456
transform 1 0 26588 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_289
timestamp 1636968456
transform 1 0 27692 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_301
timestamp 1
transform 1 0 28796 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_307
timestamp 1
transform 1 0 29348 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_309
timestamp 1636968456
transform 1 0 29532 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_321
timestamp 1636968456
transform 1 0 30636 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_333
timestamp 1636968456
transform 1 0 31740 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_345
timestamp 1636968456
transform 1 0 32844 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_357
timestamp 1
transform 1 0 33948 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_363
timestamp 1
transform 1 0 34500 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_365
timestamp 1636968456
transform 1 0 34684 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_377
timestamp 1636968456
transform 1 0 35788 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_389
timestamp 1
transform 1 0 36892 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_393
timestamp 1
transform 1 0 37260 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_405
timestamp 1636968456
transform 1 0 38364 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_130_417
timestamp 1
transform 1 0 39468 0 1 72896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_130_432
timestamp 1636968456
transform 1 0 40848 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_444
timestamp 1636968456
transform 1 0 41952 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_456
timestamp 1636968456
transform 1 0 43056 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_468
timestamp 1
transform 1 0 44160 0 1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_130_477
timestamp 1636968456
transform 1 0 44988 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_489
timestamp 1636968456
transform 1 0 46092 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_501
timestamp 1636968456
transform 1 0 47196 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_513
timestamp 1636968456
transform 1 0 48300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_525
timestamp 1
transform 1 0 49404 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_531
timestamp 1
transform 1 0 49956 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_533
timestamp 1636968456
transform 1 0 50140 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_545
timestamp 1636968456
transform 1 0 51244 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_557
timestamp 1636968456
transform 1 0 52348 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_569
timestamp 1636968456
transform 1 0 53452 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_581
timestamp 1
transform 1 0 54556 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_587
timestamp 1
transform 1 0 55108 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_589
timestamp 1636968456
transform 1 0 55292 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_601
timestamp 1636968456
transform 1 0 56396 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_613
timestamp 1636968456
transform 1 0 57500 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_625
timestamp 1636968456
transform 1 0 58604 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_637
timestamp 1
transform 1 0 59708 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_643
timestamp 1
transform 1 0 60260 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_645
timestamp 1636968456
transform 1 0 60444 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_657
timestamp 1636968456
transform 1 0 61548 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_669
timestamp 1636968456
transform 1 0 62652 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_681
timestamp 1636968456
transform 1 0 63756 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_693
timestamp 1
transform 1 0 64860 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_699
timestamp 1
transform 1 0 65412 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_701
timestamp 1636968456
transform 1 0 65596 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_713
timestamp 1636968456
transform 1 0 66700 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_725
timestamp 1
transform 1 0 67804 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_755
timestamp 1
transform 1 0 70564 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_757
timestamp 1636968456
transform 1 0 70748 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_769
timestamp 1
transform 1 0 71852 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_773
timestamp 1
transform 1 0 72220 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_785
timestamp 1636968456
transform 1 0 73324 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_797
timestamp 1636968456
transform 1 0 74428 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_130_809
timestamp 1
transform 1 0 75532 0 1 72896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_130_813
timestamp 1636968456
transform 1 0 75900 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_825
timestamp 1636968456
transform 1 0 77004 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_837
timestamp 1
transform 1 0 78108 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_841
timestamp 1
transform 1 0 78476 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_860
timestamp 1
transform 1 0 80224 0 1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_130_869
timestamp 1636968456
transform 1 0 81052 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_881
timestamp 1636968456
transform 1 0 82156 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_893
timestamp 1636968456
transform 1 0 83260 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_905
timestamp 1636968456
transform 1 0 84364 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_917
timestamp 1
transform 1 0 85468 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_923
timestamp 1
transform 1 0 86020 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_925
timestamp 1636968456
transform 1 0 86204 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_937
timestamp 1
transform 1 0 87308 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_941
timestamp 1
transform 1 0 87676 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_947
timestamp 1636968456
transform 1 0 88228 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_959
timestamp 1636968456
transform 1 0 89332 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_971
timestamp 1
transform 1 0 90436 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_979
timestamp 1
transform 1 0 91172 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_981
timestamp 1636968456
transform 1 0 91356 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_993
timestamp 1636968456
transform 1 0 92460 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_130_1005
timestamp 1
transform 1 0 93564 0 1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1009
timestamp 1636968456
transform 1 0 93932 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_1021
timestamp 1
transform 1 0 95036 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1025
timestamp 1
transform 1 0 95404 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_130_1031
timestamp 1
transform 1 0 95956 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1035
timestamp 1
transform 1 0 96324 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_130_1037
timestamp 1
transform 1 0 96508 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_130_1063
timestamp 1
transform 1 0 98900 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_130_1073
timestamp 1
transform 1 0 99820 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1077
timestamp 1
transform 1 0 100188 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1091
timestamp 1
transform 1 0 101476 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1110
timestamp 1
transform 1 0 103224 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1118
timestamp 1
transform 1 0 103960 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_1125
timestamp 1
transform 1 0 104604 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_130_1144
timestamp 1
transform 1 0 106352 0 1 72896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1149
timestamp 1636968456
transform 1 0 106812 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_130_1161
timestamp 1
transform 1 0 107916 0 1 72896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_131_9
timestamp 1636968456
transform 1 0 1932 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_21
timestamp 1636968456
transform 1 0 3036 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_33
timestamp 1636968456
transform 1 0 4140 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_45
timestamp 1
transform 1 0 5244 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_131_53
timestamp 1
transform 1 0 5980 0 -1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_131_57
timestamp 1636968456
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_69
timestamp 1636968456
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_81
timestamp 1636968456
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_93
timestamp 1636968456
transform 1 0 9660 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_105
timestamp 1
transform 1 0 10764 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_109
timestamp 1
transform 1 0 11132 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_131_113
timestamp 1
transform 1 0 11500 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_136
timestamp 1636968456
transform 1 0 13616 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_148
timestamp 1636968456
transform 1 0 14720 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_160
timestamp 1
transform 1 0 15824 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_131_169
timestamp 1
transform 1 0 16652 0 -1 73984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_131_195
timestamp 1636968456
transform 1 0 19044 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_207
timestamp 1636968456
transform 1 0 20148 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_219
timestamp 1
transform 1 0 21252 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_223
timestamp 1
transform 1 0 21620 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_225
timestamp 1636968456
transform 1 0 21804 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_237
timestamp 1
transform 1 0 22908 0 -1 73984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_131_265
timestamp 1636968456
transform 1 0 25484 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_277
timestamp 1
transform 1 0 26588 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_131_281
timestamp 1
transform 1 0 26956 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_131_289
timestamp 1
transform 1 0 27692 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_295
timestamp 1636968456
transform 1 0 28244 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_307
timestamp 1636968456
transform 1 0 29348 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_319
timestamp 1636968456
transform 1 0 30452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_331
timestamp 1
transform 1 0 31556 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_335
timestamp 1
transform 1 0 31924 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_337
timestamp 1636968456
transform 1 0 32108 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_349
timestamp 1636968456
transform 1 0 33212 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_361
timestamp 1
transform 1 0 34316 0 -1 73984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_131_380
timestamp 1636968456
transform 1 0 36064 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_393
timestamp 1636968456
transform 1 0 37260 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_405
timestamp 1636968456
transform 1 0 38364 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_417
timestamp 1636968456
transform 1 0 39468 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_429
timestamp 1636968456
transform 1 0 40572 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_441
timestamp 1
transform 1 0 41676 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_447
timestamp 1
transform 1 0 42228 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_449
timestamp 1636968456
transform 1 0 42412 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_461
timestamp 1636968456
transform 1 0 43516 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_473
timestamp 1636968456
transform 1 0 44620 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_485
timestamp 1636968456
transform 1 0 45724 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_497
timestamp 1
transform 1 0 46828 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_503
timestamp 1
transform 1 0 47380 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_505
timestamp 1636968456
transform 1 0 47564 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_517
timestamp 1636968456
transform 1 0 48668 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_529
timestamp 1636968456
transform 1 0 49772 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_541
timestamp 1636968456
transform 1 0 50876 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_553
timestamp 1
transform 1 0 51980 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_559
timestamp 1
transform 1 0 52532 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_561
timestamp 1636968456
transform 1 0 52716 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_573
timestamp 1636968456
transform 1 0 53820 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_585
timestamp 1
transform 1 0 54924 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_131_611
timestamp 1
transform 1 0 57316 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_615
timestamp 1
transform 1 0 57684 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_617
timestamp 1636968456
transform 1 0 57868 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_629
timestamp 1636968456
transform 1 0 58972 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_641
timestamp 1636968456
transform 1 0 60076 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_653
timestamp 1636968456
transform 1 0 61180 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_665
timestamp 1
transform 1 0 62284 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_671
timestamp 1
transform 1 0 62836 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_673
timestamp 1636968456
transform 1 0 63020 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_685
timestamp 1636968456
transform 1 0 64124 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_697
timestamp 1636968456
transform 1 0 65228 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_709
timestamp 1636968456
transform 1 0 66332 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_721
timestamp 1
transform 1 0 67436 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_727
timestamp 1
transform 1 0 67988 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_131_740
timestamp 1
transform 1 0 69184 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_746
timestamp 1
transform 1 0 69736 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_758
timestamp 1636968456
transform 1 0 70840 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_770
timestamp 1636968456
transform 1 0 71944 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_782
timestamp 1
transform 1 0 73048 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_131_793
timestamp 1
transform 1 0 74060 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_805
timestamp 1636968456
transform 1 0 75164 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_817
timestamp 1636968456
transform 1 0 76268 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_829
timestamp 1
transform 1 0 77372 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_131_837
timestamp 1
transform 1 0 78108 0 -1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_131_841
timestamp 1636968456
transform 1 0 78476 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_853
timestamp 1636968456
transform 1 0 79580 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_865
timestamp 1636968456
transform 1 0 80684 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_877
timestamp 1636968456
transform 1 0 81788 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_889
timestamp 1
transform 1 0 82892 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_895
timestamp 1
transform 1 0 83444 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_897
timestamp 1636968456
transform 1 0 83628 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_914
timestamp 1
transform 1 0 85192 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_131_941
timestamp 1
transform 1 0 87676 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_131_949
timestamp 1
transform 1 0 88412 0 -1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_131_982
timestamp 1636968456
transform 1 0 91448 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_994
timestamp 1
transform 1 0 92552 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1007
timestamp 1
transform 1 0 93748 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1017
timestamp 1636968456
transform 1 0 94668 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1029
timestamp 1636968456
transform 1 0 95772 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1041
timestamp 1636968456
transform 1 0 96876 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1053
timestamp 1
transform 1 0 97980 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1059
timestamp 1
transform 1 0 98532 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1083
timestamp 1636968456
transform 1 0 100740 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_1098
timestamp 1
transform 1 0 102120 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_131_1105
timestamp 1
transform 1 0 102764 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_131_1115
timestamp 1
transform 1 0 103684 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1119
timestamp 1
transform 1 0 104052 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_131_1129
timestamp 1
transform 1 0 104972 0 -1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1139
timestamp 1636968456
transform 1 0 105892 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1151
timestamp 1636968456
transform 1 0 106996 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_9
timestamp 1636968456
transform 1 0 1932 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_21
timestamp 1
transform 1 0 3036 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1636968456
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_41
timestamp 1636968456
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_53
timestamp 1636968456
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_65
timestamp 1636968456
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_85
timestamp 1636968456
transform 1 0 8924 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_97
timestamp 1636968456
transform 1 0 10028 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_109
timestamp 1636968456
transform 1 0 11132 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_121
timestamp 1636968456
transform 1 0 12236 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_133
timestamp 1
transform 1 0 13340 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_139
timestamp 1
transform 1 0 13892 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_141
timestamp 1636968456
transform 1 0 14076 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_153
timestamp 1636968456
transform 1 0 15180 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_165
timestamp 1636968456
transform 1 0 16284 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_177
timestamp 1636968456
transform 1 0 17388 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_189
timestamp 1
transform 1 0 18492 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_195
timestamp 1
transform 1 0 19044 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_197
timestamp 1636968456
transform 1 0 19228 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_209
timestamp 1636968456
transform 1 0 20332 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_132_221
timestamp 1
transform 1 0 21436 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_132_249
timestamp 1
transform 1 0 24012 0 1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_132_258
timestamp 1636968456
transform 1 0 24840 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_270
timestamp 1636968456
transform 1 0 25944 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_282
timestamp 1
transform 1 0 27048 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_132_290
timestamp 1
transform 1 0 27784 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_132_298
timestamp 1
transform 1 0 28520 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_132_306
timestamp 1
transform 1 0 29256 0 1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_132_314
timestamp 1636968456
transform 1 0 29992 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_326
timestamp 1636968456
transform 1 0 31096 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_338
timestamp 1636968456
transform 1 0 32200 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_350
timestamp 1636968456
transform 1 0 33304 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_132_362
timestamp 1
transform 1 0 34408 0 1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_132_365
timestamp 1636968456
transform 1 0 34684 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_377
timestamp 1636968456
transform 1 0 35788 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_389
timestamp 1636968456
transform 1 0 36892 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_401
timestamp 1636968456
transform 1 0 37996 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_413
timestamp 1
transform 1 0 39100 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_419
timestamp 1
transform 1 0 39652 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_421
timestamp 1636968456
transform 1 0 39836 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_433
timestamp 1636968456
transform 1 0 40940 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_445
timestamp 1636968456
transform 1 0 42044 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_457
timestamp 1636968456
transform 1 0 43148 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_469
timestamp 1
transform 1 0 44252 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_475
timestamp 1
transform 1 0 44804 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_477
timestamp 1636968456
transform 1 0 44988 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_489
timestamp 1636968456
transform 1 0 46092 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_501
timestamp 1636968456
transform 1 0 47196 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_513
timestamp 1636968456
transform 1 0 48300 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_525
timestamp 1
transform 1 0 49404 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_531
timestamp 1
transform 1 0 49956 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_533
timestamp 1636968456
transform 1 0 50140 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_545
timestamp 1636968456
transform 1 0 51244 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_557
timestamp 1636968456
transform 1 0 52348 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_569
timestamp 1636968456
transform 1 0 53452 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_581
timestamp 1
transform 1 0 54556 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_587
timestamp 1
transform 1 0 55108 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_589
timestamp 1636968456
transform 1 0 55292 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_601
timestamp 1636968456
transform 1 0 56396 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_613
timestamp 1636968456
transform 1 0 57500 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_625
timestamp 1636968456
transform 1 0 58604 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_637
timestamp 1
transform 1 0 59708 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_643
timestamp 1
transform 1 0 60260 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_645
timestamp 1636968456
transform 1 0 60444 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_657
timestamp 1636968456
transform 1 0 61548 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_669
timestamp 1636968456
transform 1 0 62652 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_681
timestamp 1636968456
transform 1 0 63756 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_693
timestamp 1
transform 1 0 64860 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_699
timestamp 1
transform 1 0 65412 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_701
timestamp 1636968456
transform 1 0 65596 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_713
timestamp 1636968456
transform 1 0 66700 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_725
timestamp 1636968456
transform 1 0 67804 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_737
timestamp 1636968456
transform 1 0 68908 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_749
timestamp 1
transform 1 0 70012 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_755
timestamp 1
transform 1 0 70564 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_757
timestamp 1636968456
transform 1 0 70748 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_769
timestamp 1636968456
transform 1 0 71852 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_781
timestamp 1636968456
transform 1 0 72956 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_793
timestamp 1
transform 1 0 74060 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_132_805
timestamp 1
transform 1 0 75164 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_811
timestamp 1
transform 1 0 75716 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_813
timestamp 1636968456
transform 1 0 75900 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_825
timestamp 1636968456
transform 1 0 77004 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_837
timestamp 1636968456
transform 1 0 78108 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_849
timestamp 1636968456
transform 1 0 79212 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_861
timestamp 1
transform 1 0 80316 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_867
timestamp 1
transform 1 0 80868 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_869
timestamp 1636968456
transform 1 0 81052 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_881
timestamp 1636968456
transform 1 0 82156 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_893
timestamp 1636968456
transform 1 0 83260 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_905
timestamp 1636968456
transform 1 0 84364 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_917
timestamp 1
transform 1 0 85468 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_132_923
timestamp 1
transform 1 0 86020 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_925
timestamp 1
transform 1 0 86204 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_132_933
timestamp 1
transform 1 0 86940 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_132_940
timestamp 1
transform 1 0 87584 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_132_972
timestamp 1
transform 1 0 90528 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_981
timestamp 1
transform 1 0 91356 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_987
timestamp 1636968456
transform 1 0 91908 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_999
timestamp 1636968456
transform 1 0 93012 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1011
timestamp 1636968456
transform 1 0 94116 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1023
timestamp 1636968456
transform 1 0 95220 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1035
timestamp 1
transform 1 0 96324 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1037
timestamp 1
transform 1 0 96508 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_132_1045
timestamp 1
transform 1 0 97244 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1049
timestamp 1
transform 1 0 97612 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1058
timestamp 1636968456
transform 1 0 98440 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_132_1070
timestamp 1
transform 1 0 99544 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_132_1082
timestamp 1
transform 1 0 100648 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1088
timestamp 1
transform 1 0 101200 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_132_1100
timestamp 1
transform 1 0 102304 0 1 73984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1111
timestamp 1636968456
transform 1 0 103316 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1127
timestamp 1
transform 1 0 104788 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_1137
timestamp 1
transform 1 0 105708 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_132_1145
timestamp 1
transform 1 0 106444 0 1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1149
timestamp 1636968456
transform 1 0 106812 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1161
timestamp 1
transform 1 0 107916 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636968456
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636968456
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1636968456
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_39
timestamp 1636968456
transform 1 0 4692 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_51
timestamp 1
transform 1 0 5796 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_55
timestamp 1
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_57
timestamp 1636968456
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_69
timestamp 1636968456
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_81
timestamp 1636968456
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_93
timestamp 1636968456
transform 1 0 9660 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_105
timestamp 1
transform 1 0 10764 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_111
timestamp 1
transform 1 0 11316 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_113
timestamp 1636968456
transform 1 0 11500 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_125
timestamp 1636968456
transform 1 0 12604 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_137
timestamp 1636968456
transform 1 0 13708 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_149
timestamp 1636968456
transform 1 0 14812 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_161
timestamp 1
transform 1 0 15916 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_167
timestamp 1
transform 1 0 16468 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_169
timestamp 1636968456
transform 1 0 16652 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_181
timestamp 1
transform 1 0 17756 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_205
timestamp 1636968456
transform 1 0 19964 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_217
timestamp 1
transform 1 0 21068 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_223
timestamp 1
transform 1 0 21620 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_225
timestamp 1636968456
transform 1 0 21804 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_237
timestamp 1636968456
transform 1 0 22908 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_249
timestamp 1636968456
transform 1 0 24012 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_261
timestamp 1636968456
transform 1 0 25116 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_273
timestamp 1
transform 1 0 26220 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_279
timestamp 1
transform 1 0 26772 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_281
timestamp 1636968456
transform 1 0 26956 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_293
timestamp 1636968456
transform 1 0 28060 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_305
timestamp 1636968456
transform 1 0 29164 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_317
timestamp 1636968456
transform 1 0 30268 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_329
timestamp 1
transform 1 0 31372 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_335
timestamp 1
transform 1 0 31924 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_337
timestamp 1636968456
transform 1 0 32108 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_349
timestamp 1636968456
transform 1 0 33212 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_361
timestamp 1636968456
transform 1 0 34316 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_373
timestamp 1636968456
transform 1 0 35420 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_385
timestamp 1
transform 1 0 36524 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_391
timestamp 1
transform 1 0 37076 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_393
timestamp 1636968456
transform 1 0 37260 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_405
timestamp 1636968456
transform 1 0 38364 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_417
timestamp 1636968456
transform 1 0 39468 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_429
timestamp 1636968456
transform 1 0 40572 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_441
timestamp 1
transform 1 0 41676 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_447
timestamp 1
transform 1 0 42228 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_449
timestamp 1636968456
transform 1 0 42412 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_461
timestamp 1636968456
transform 1 0 43516 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_473
timestamp 1636968456
transform 1 0 44620 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_485
timestamp 1636968456
transform 1 0 45724 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_497
timestamp 1
transform 1 0 46828 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_503
timestamp 1
transform 1 0 47380 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_505
timestamp 1636968456
transform 1 0 47564 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_517
timestamp 1636968456
transform 1 0 48668 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_529
timestamp 1636968456
transform 1 0 49772 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_541
timestamp 1636968456
transform 1 0 50876 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_553
timestamp 1
transform 1 0 51980 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_559
timestamp 1
transform 1 0 52532 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_561
timestamp 1636968456
transform 1 0 52716 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_573
timestamp 1636968456
transform 1 0 53820 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_585
timestamp 1636968456
transform 1 0 54924 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_597
timestamp 1636968456
transform 1 0 56028 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_609
timestamp 1
transform 1 0 57132 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_615
timestamp 1
transform 1 0 57684 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_617
timestamp 1636968456
transform 1 0 57868 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_629
timestamp 1636968456
transform 1 0 58972 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_641
timestamp 1636968456
transform 1 0 60076 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_653
timestamp 1636968456
transform 1 0 61180 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_665
timestamp 1
transform 1 0 62284 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_671
timestamp 1
transform 1 0 62836 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_673
timestamp 1636968456
transform 1 0 63020 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_685
timestamp 1636968456
transform 1 0 64124 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_697
timestamp 1636968456
transform 1 0 65228 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_709
timestamp 1636968456
transform 1 0 66332 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_721
timestamp 1
transform 1 0 67436 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_727
timestamp 1
transform 1 0 67988 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_729
timestamp 1636968456
transform 1 0 68172 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_741
timestamp 1636968456
transform 1 0 69276 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_753
timestamp 1636968456
transform 1 0 70380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_765
timestamp 1636968456
transform 1 0 71484 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_777
timestamp 1
transform 1 0 72588 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_783
timestamp 1
transform 1 0 73140 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_785
timestamp 1636968456
transform 1 0 73324 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_797
timestamp 1636968456
transform 1 0 74428 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_809
timestamp 1636968456
transform 1 0 75532 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_821
timestamp 1636968456
transform 1 0 76636 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_833
timestamp 1
transform 1 0 77740 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_839
timestamp 1
transform 1 0 78292 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_841
timestamp 1636968456
transform 1 0 78476 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_853
timestamp 1636968456
transform 1 0 79580 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_865
timestamp 1636968456
transform 1 0 80684 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_877
timestamp 1636968456
transform 1 0 81788 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_889
timestamp 1
transform 1 0 82892 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_895
timestamp 1
transform 1 0 83444 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_897
timestamp 1636968456
transform 1 0 83628 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_909
timestamp 1636968456
transform 1 0 84732 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_921
timestamp 1
transform 1 0 85836 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_133_950
timestamp 1
transform 1 0 88504 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_133_953
timestamp 1
transform 1 0 88780 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_133_966
timestamp 1
transform 1 0 89976 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_974
timestamp 1
transform 1 0 90712 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_994
timestamp 1636968456
transform 1 0 92552 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_133_1006
timestamp 1
transform 1 0 93656 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1009
timestamp 1
transform 1 0 93932 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1017
timestamp 1636968456
transform 1 0 94668 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_1029
timestamp 1
transform 1 0 95772 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1035
timestamp 1
transform 1 0 96324 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_133_1051
timestamp 1
transform 1 0 97796 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_133_1062
timestamp 1
transform 1 0 98808 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1073
timestamp 1
transform 1 0 99820 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_133_1101
timestamp 1
transform 1 0 102396 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1107
timestamp 1
transform 1 0 102948 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_133_1121
timestamp 1
transform 1 0 104236 0 -1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1136
timestamp 1636968456
transform 1 0 105616 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1148
timestamp 1636968456
transform 1 0 106720 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_1160
timestamp 1
transform 1 0 107824 0 -1 75072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_134_7
timestamp 1636968456
transform 1 0 1748 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_19
timestamp 1
transform 1 0 2852 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1636968456
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_41
timestamp 1636968456
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_53
timestamp 1636968456
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_65
timestamp 1636968456
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_85
timestamp 1636968456
transform 1 0 8924 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_97
timestamp 1636968456
transform 1 0 10028 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_109
timestamp 1636968456
transform 1 0 11132 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_121
timestamp 1636968456
transform 1 0 12236 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_133
timestamp 1
transform 1 0 13340 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_139
timestamp 1
transform 1 0 13892 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_141
timestamp 1636968456
transform 1 0 14076 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_153
timestamp 1636968456
transform 1 0 15180 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_165
timestamp 1636968456
transform 1 0 16284 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_177
timestamp 1636968456
transform 1 0 17388 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_189
timestamp 1
transform 1 0 18492 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_195
timestamp 1
transform 1 0 19044 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_197
timestamp 1636968456
transform 1 0 19228 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_209
timestamp 1636968456
transform 1 0 20332 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_221
timestamp 1
transform 1 0 21436 0 1 75072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_134_234
timestamp 1636968456
transform 1 0 22632 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_246
timestamp 1
transform 1 0 23736 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_134_253
timestamp 1
transform 1 0 24380 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_134_261
timestamp 1
transform 1 0 25116 0 1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_134_269
timestamp 1636968456
transform 1 0 25852 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_281
timestamp 1636968456
transform 1 0 26956 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_293
timestamp 1636968456
transform 1 0 28060 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_134_305
timestamp 1
transform 1 0 29164 0 1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_134_309
timestamp 1636968456
transform 1 0 29532 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_321
timestamp 1636968456
transform 1 0 30636 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_333
timestamp 1636968456
transform 1 0 31740 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_345
timestamp 1636968456
transform 1 0 32844 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_357
timestamp 1
transform 1 0 33948 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_363
timestamp 1
transform 1 0 34500 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_365
timestamp 1636968456
transform 1 0 34684 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_377
timestamp 1636968456
transform 1 0 35788 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_389
timestamp 1636968456
transform 1 0 36892 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_401
timestamp 1636968456
transform 1 0 37996 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_413
timestamp 1
transform 1 0 39100 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_419
timestamp 1
transform 1 0 39652 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_421
timestamp 1636968456
transform 1 0 39836 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_433
timestamp 1636968456
transform 1 0 40940 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_445
timestamp 1636968456
transform 1 0 42044 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_457
timestamp 1636968456
transform 1 0 43148 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_469
timestamp 1
transform 1 0 44252 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_475
timestamp 1
transform 1 0 44804 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_477
timestamp 1636968456
transform 1 0 44988 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_489
timestamp 1636968456
transform 1 0 46092 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_501
timestamp 1636968456
transform 1 0 47196 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_513
timestamp 1636968456
transform 1 0 48300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_525
timestamp 1
transform 1 0 49404 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_531
timestamp 1
transform 1 0 49956 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_533
timestamp 1636968456
transform 1 0 50140 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_545
timestamp 1636968456
transform 1 0 51244 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_557
timestamp 1636968456
transform 1 0 52348 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_569
timestamp 1636968456
transform 1 0 53452 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_581
timestamp 1
transform 1 0 54556 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_587
timestamp 1
transform 1 0 55108 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_589
timestamp 1636968456
transform 1 0 55292 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_601
timestamp 1636968456
transform 1 0 56396 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_613
timestamp 1636968456
transform 1 0 57500 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_625
timestamp 1636968456
transform 1 0 58604 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_637
timestamp 1
transform 1 0 59708 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_643
timestamp 1
transform 1 0 60260 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_645
timestamp 1636968456
transform 1 0 60444 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_657
timestamp 1636968456
transform 1 0 61548 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_669
timestamp 1636968456
transform 1 0 62652 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_681
timestamp 1636968456
transform 1 0 63756 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_693
timestamp 1
transform 1 0 64860 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_699
timestamp 1
transform 1 0 65412 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_701
timestamp 1636968456
transform 1 0 65596 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_713
timestamp 1636968456
transform 1 0 66700 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_725
timestamp 1636968456
transform 1 0 67804 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_737
timestamp 1636968456
transform 1 0 68908 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_749
timestamp 1
transform 1 0 70012 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_755
timestamp 1
transform 1 0 70564 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_757
timestamp 1636968456
transform 1 0 70748 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_769
timestamp 1636968456
transform 1 0 71852 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_781
timestamp 1636968456
transform 1 0 72956 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_793
timestamp 1636968456
transform 1 0 74060 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_805
timestamp 1
transform 1 0 75164 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_811
timestamp 1
transform 1 0 75716 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_813
timestamp 1636968456
transform 1 0 75900 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_825
timestamp 1636968456
transform 1 0 77004 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_837
timestamp 1636968456
transform 1 0 78108 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_849
timestamp 1636968456
transform 1 0 79212 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_861
timestamp 1
transform 1 0 80316 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_867
timestamp 1
transform 1 0 80868 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_869
timestamp 1636968456
transform 1 0 81052 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_881
timestamp 1636968456
transform 1 0 82156 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_893
timestamp 1636968456
transform 1 0 83260 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_905
timestamp 1636968456
transform 1 0 84364 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_917
timestamp 1
transform 1 0 85468 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_923
timestamp 1
transform 1 0 86020 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_925
timestamp 1636968456
transform 1 0 86204 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_134_937
timestamp 1
transform 1 0 87308 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_134_951
timestamp 1
transform 1 0 88596 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_134_977
timestamp 1
transform 1 0 90988 0 1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_134_981
timestamp 1636968456
transform 1 0 91356 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_134_993
timestamp 1
transform 1 0 92460 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_134_997
timestamp 1
transform 1 0 92828 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1020
timestamp 1636968456
transform 1 0 94944 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_134_1032
timestamp 1
transform 1 0 96048 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_134_1037
timestamp 1
transform 1 0 96508 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_134_1052
timestamp 1
transform 1 0 97888 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_134_1058
timestamp 1
transform 1 0 98440 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1062
timestamp 1
transform 1 0 98808 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1066
timestamp 1636968456
transform 1 0 99176 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_134_1081
timestamp 1
transform 1 0 100556 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_134_1100
timestamp 1
transform 1 0 102304 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1104
timestamp 1
transform 1 0 102672 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1134
timestamp 1636968456
transform 1 0 105432 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_134_1146
timestamp 1
transform 1 0 106536 0 1 75072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1149
timestamp 1636968456
transform 1 0 106812 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1161
timestamp 1
transform 1 0 107916 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_7
timestamp 1636968456
transform 1 0 1748 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_19
timestamp 1636968456
transform 1 0 2852 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_31
timestamp 1636968456
transform 1 0 3956 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_43
timestamp 1636968456
transform 1 0 5060 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_135_55
timestamp 1
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_57
timestamp 1636968456
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_69
timestamp 1636968456
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_81
timestamp 1636968456
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_93
timestamp 1636968456
transform 1 0 9660 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_105
timestamp 1
transform 1 0 10764 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_111
timestamp 1
transform 1 0 11316 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_113
timestamp 1636968456
transform 1 0 11500 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_125
timestamp 1636968456
transform 1 0 12604 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_137
timestamp 1
transform 1 0 13708 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_135_145
timestamp 1
transform 1 0 14444 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_169
timestamp 1636968456
transform 1 0 16652 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_181
timestamp 1636968456
transform 1 0 17756 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_193
timestamp 1636968456
transform 1 0 18860 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_205
timestamp 1636968456
transform 1 0 19964 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_217
timestamp 1
transform 1 0 21068 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_223
timestamp 1
transform 1 0 21620 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_225
timestamp 1636968456
transform 1 0 21804 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_237
timestamp 1636968456
transform 1 0 22908 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_249
timestamp 1636968456
transform 1 0 24012 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_261
timestamp 1636968456
transform 1 0 25116 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_273
timestamp 1
transform 1 0 26220 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_279
timestamp 1
transform 1 0 26772 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_281
timestamp 1636968456
transform 1 0 26956 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_293
timestamp 1636968456
transform 1 0 28060 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_305
timestamp 1636968456
transform 1 0 29164 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_317
timestamp 1636968456
transform 1 0 30268 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_329
timestamp 1
transform 1 0 31372 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_335
timestamp 1
transform 1 0 31924 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_337
timestamp 1636968456
transform 1 0 32108 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_349
timestamp 1636968456
transform 1 0 33212 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_361
timestamp 1636968456
transform 1 0 34316 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_373
timestamp 1636968456
transform 1 0 35420 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_385
timestamp 1
transform 1 0 36524 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_391
timestamp 1
transform 1 0 37076 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_393
timestamp 1636968456
transform 1 0 37260 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_405
timestamp 1636968456
transform 1 0 38364 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_417
timestamp 1636968456
transform 1 0 39468 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_429
timestamp 1636968456
transform 1 0 40572 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_441
timestamp 1
transform 1 0 41676 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_447
timestamp 1
transform 1 0 42228 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_449
timestamp 1636968456
transform 1 0 42412 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_461
timestamp 1636968456
transform 1 0 43516 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_473
timestamp 1636968456
transform 1 0 44620 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_485
timestamp 1636968456
transform 1 0 45724 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_497
timestamp 1
transform 1 0 46828 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_503
timestamp 1
transform 1 0 47380 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_505
timestamp 1636968456
transform 1 0 47564 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_517
timestamp 1636968456
transform 1 0 48668 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_529
timestamp 1636968456
transform 1 0 49772 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_541
timestamp 1636968456
transform 1 0 50876 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_553
timestamp 1
transform 1 0 51980 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_559
timestamp 1
transform 1 0 52532 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_561
timestamp 1636968456
transform 1 0 52716 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_573
timestamp 1636968456
transform 1 0 53820 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_585
timestamp 1636968456
transform 1 0 54924 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_597
timestamp 1636968456
transform 1 0 56028 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_609
timestamp 1
transform 1 0 57132 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_615
timestamp 1
transform 1 0 57684 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_617
timestamp 1636968456
transform 1 0 57868 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_629
timestamp 1636968456
transform 1 0 58972 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_641
timestamp 1636968456
transform 1 0 60076 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_653
timestamp 1636968456
transform 1 0 61180 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_665
timestamp 1
transform 1 0 62284 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_671
timestamp 1
transform 1 0 62836 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_673
timestamp 1636968456
transform 1 0 63020 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_685
timestamp 1636968456
transform 1 0 64124 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_697
timestamp 1636968456
transform 1 0 65228 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_709
timestamp 1636968456
transform 1 0 66332 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_721
timestamp 1
transform 1 0 67436 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_727
timestamp 1
transform 1 0 67988 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_729
timestamp 1636968456
transform 1 0 68172 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_741
timestamp 1636968456
transform 1 0 69276 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_753
timestamp 1636968456
transform 1 0 70380 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_765
timestamp 1636968456
transform 1 0 71484 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_777
timestamp 1
transform 1 0 72588 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_783
timestamp 1
transform 1 0 73140 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_785
timestamp 1636968456
transform 1 0 73324 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_797
timestamp 1636968456
transform 1 0 74428 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_809
timestamp 1636968456
transform 1 0 75532 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_821
timestamp 1636968456
transform 1 0 76636 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_833
timestamp 1
transform 1 0 77740 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_839
timestamp 1
transform 1 0 78292 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_841
timestamp 1636968456
transform 1 0 78476 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_853
timestamp 1636968456
transform 1 0 79580 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_865
timestamp 1636968456
transform 1 0 80684 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_877
timestamp 1636968456
transform 1 0 81788 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_889
timestamp 1
transform 1 0 82892 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_895
timestamp 1
transform 1 0 83444 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_899
timestamp 1636968456
transform 1 0 83812 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_911
timestamp 1636968456
transform 1 0 84916 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_923
timestamp 1636968456
transform 1 0 86020 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_935
timestamp 1
transform 1 0 87124 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_135_947
timestamp 1
transform 1 0 88228 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_951
timestamp 1
transform 1 0 88596 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_955
timestamp 1
transform 1 0 88964 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_963
timestamp 1
transform 1 0 89700 0 -1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_135_970
timestamp 1
transform 1 0 90344 0 -1 76160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_135_979
timestamp 1636968456
transform 1 0 91172 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_991
timestamp 1636968456
transform 1 0 92276 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_1003
timestamp 1
transform 1 0 93380 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1007
timestamp 1
transform 1 0 93748 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_1009
timestamp 1
transform 1 0 93932 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_135_1017
timestamp 1
transform 1 0 94668 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1042
timestamp 1
transform 1 0 96968 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1048
timestamp 1
transform 1 0 97520 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1073
timestamp 1
transform 1 0 99820 0 -1 76160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1084
timestamp 1636968456
transform 1 0 100832 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1096
timestamp 1636968456
transform 1 0 101936 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1108
timestamp 1636968456
transform 1 0 103040 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1121
timestamp 1636968456
transform 1 0 104236 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1133
timestamp 1636968456
transform 1 0 105340 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1145
timestamp 1636968456
transform 1 0 106444 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_1157
timestamp 1
transform 1 0 107548 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1161
timestamp 1
transform 1 0 107916 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_7
timestamp 1636968456
transform 1 0 1748 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_19
timestamp 1
transform 1 0 2852 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1636968456
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_41
timestamp 1636968456
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_53
timestamp 1636968456
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_65
timestamp 1636968456
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_85
timestamp 1636968456
transform 1 0 8924 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_97
timestamp 1636968456
transform 1 0 10028 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_109
timestamp 1636968456
transform 1 0 11132 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_121
timestamp 1636968456
transform 1 0 12236 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_133
timestamp 1
transform 1 0 13340 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_139
timestamp 1
transform 1 0 13892 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_141
timestamp 1636968456
transform 1 0 14076 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_153
timestamp 1636968456
transform 1 0 15180 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_165
timestamp 1636968456
transform 1 0 16284 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_177
timestamp 1636968456
transform 1 0 17388 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_189
timestamp 1
transform 1 0 18492 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_195
timestamp 1
transform 1 0 19044 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_197
timestamp 1636968456
transform 1 0 19228 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_209
timestamp 1636968456
transform 1 0 20332 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_221
timestamp 1636968456
transform 1 0 21436 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_233
timestamp 1
transform 1 0 22540 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_237
timestamp 1
transform 1 0 22908 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_136_251
timestamp 1
transform 1 0 24196 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_253
timestamp 1636968456
transform 1 0 24380 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_265
timestamp 1
transform 1 0 25484 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_136_273
timestamp 1
transform 1 0 26220 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_136_289
timestamp 1
transform 1 0 27692 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_297
timestamp 1
transform 1 0 28428 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_136_307
timestamp 1
transform 1 0 29348 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_311
timestamp 1636968456
transform 1 0 29716 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_323
timestamp 1636968456
transform 1 0 30820 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_335
timestamp 1636968456
transform 1 0 31924 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_347
timestamp 1636968456
transform 1 0 33028 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_359
timestamp 1
transform 1 0 34132 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_363
timestamp 1
transform 1 0 34500 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_365
timestamp 1636968456
transform 1 0 34684 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_377
timestamp 1636968456
transform 1 0 35788 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_389
timestamp 1636968456
transform 1 0 36892 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_401
timestamp 1636968456
transform 1 0 37996 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_413
timestamp 1
transform 1 0 39100 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_419
timestamp 1
transform 1 0 39652 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_441
timestamp 1636968456
transform 1 0 41676 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_453
timestamp 1
transform 1 0 42780 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_136_474
timestamp 1
transform 1 0 44712 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_136_477
timestamp 1
transform 1 0 44988 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_481
timestamp 1
transform 1 0 45356 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_502
timestamp 1636968456
transform 1 0 47288 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_514
timestamp 1636968456
transform 1 0 48392 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_526
timestamp 1
transform 1 0 49496 0 1 76160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_136_533
timestamp 1636968456
transform 1 0 50140 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_545
timestamp 1636968456
transform 1 0 51244 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_557
timestamp 1636968456
transform 1 0 52348 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_569
timestamp 1636968456
transform 1 0 53452 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_581
timestamp 1
transform 1 0 54556 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_587
timestamp 1
transform 1 0 55108 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_589
timestamp 1636968456
transform 1 0 55292 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_601
timestamp 1636968456
transform 1 0 56396 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_613
timestamp 1636968456
transform 1 0 57500 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_625
timestamp 1636968456
transform 1 0 58604 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_637
timestamp 1
transform 1 0 59708 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_641
timestamp 1
transform 1 0 60076 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_136_647
timestamp 1
transform 1 0 60628 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_136_664
timestamp 1
transform 1 0 62192 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_668
timestamp 1
transform 1 0 62560 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_689
timestamp 1
transform 1 0 64492 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_697
timestamp 1
transform 1 0 65228 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_136_719
timestamp 1
transform 1 0 67252 0 1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_136_741
timestamp 1636968456
transform 1 0 69276 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_136_753
timestamp 1
transform 1 0 70380 0 1 76160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_136_757
timestamp 1636968456
transform 1 0 70748 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_769
timestamp 1636968456
transform 1 0 71852 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_781
timestamp 1636968456
transform 1 0 72956 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_793
timestamp 1636968456
transform 1 0 74060 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_805
timestamp 1
transform 1 0 75164 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_811
timestamp 1
transform 1 0 75716 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_813
timestamp 1636968456
transform 1 0 75900 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_825
timestamp 1636968456
transform 1 0 77004 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_837
timestamp 1636968456
transform 1 0 78108 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_849
timestamp 1636968456
transform 1 0 79212 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_861
timestamp 1
transform 1 0 80316 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_867
timestamp 1
transform 1 0 80868 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_869
timestamp 1636968456
transform 1 0 81052 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_881
timestamp 1
transform 1 0 82156 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_136_916
timestamp 1
transform 1 0 85376 0 1 76160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_136_925
timestamp 1636968456
transform 1 0 86204 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_937
timestamp 1636968456
transform 1 0 87308 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_949
timestamp 1636968456
transform 1 0 88412 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_961
timestamp 1636968456
transform 1 0 89516 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_973
timestamp 1
transform 1 0 90620 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_979
timestamp 1
transform 1 0 91172 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_981
timestamp 1636968456
transform 1 0 91356 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_993
timestamp 1
transform 1 0 92460 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1016
timestamp 1636968456
transform 1 0 94576 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_1028
timestamp 1
transform 1 0 95680 0 1 76160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1037
timestamp 1636968456
transform 1 0 96508 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1049
timestamp 1
transform 1 0 97612 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_136_1090
timestamp 1
transform 1 0 101384 0 1 76160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1093
timestamp 1636968456
transform 1 0 101660 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1105
timestamp 1636968456
transform 1 0 102764 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1117
timestamp 1636968456
transform 1 0 103868 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1129
timestamp 1636968456
transform 1 0 104972 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_1141
timestamp 1
transform 1 0 106076 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1147
timestamp 1
transform 1 0 106628 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1149
timestamp 1636968456
transform 1 0 106812 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1161
timestamp 1
transform 1 0 107916 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_11
timestamp 1636968456
transform 1 0 2116 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_23
timestamp 1636968456
transform 1 0 3220 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_35
timestamp 1636968456
transform 1 0 4324 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_47
timestamp 1
transform 1 0 5428 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_57
timestamp 1636968456
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_69
timestamp 1636968456
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_81
timestamp 1636968456
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_93
timestamp 1636968456
transform 1 0 9660 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_105
timestamp 1
transform 1 0 10764 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_111
timestamp 1
transform 1 0 11316 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_113
timestamp 1636968456
transform 1 0 11500 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_125
timestamp 1636968456
transform 1 0 12604 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_137
timestamp 1636968456
transform 1 0 13708 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_149
timestamp 1636968456
transform 1 0 14812 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_161
timestamp 1
transform 1 0 15916 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_167
timestamp 1
transform 1 0 16468 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_169
timestamp 1636968456
transform 1 0 16652 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_181
timestamp 1636968456
transform 1 0 17756 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_193
timestamp 1636968456
transform 1 0 18860 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_205
timestamp 1636968456
transform 1 0 19964 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_217
timestamp 1
transform 1 0 21068 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_223
timestamp 1
transform 1 0 21620 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_137_225
timestamp 1
transform 1 0 21804 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_229
timestamp 1
transform 1 0 22172 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_235
timestamp 1636968456
transform 1 0 22724 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_247
timestamp 1
transform 1 0 23828 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_137_255
timestamp 1
transform 1 0 24564 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_137_258
timestamp 1
transform 1 0 24840 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_275
timestamp 1
transform 1 0 26404 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_279
timestamp 1
transform 1 0 26772 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_281
timestamp 1636968456
transform 1 0 26956 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_293
timestamp 1636968456
transform 1 0 28060 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_305
timestamp 1636968456
transform 1 0 29164 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_317
timestamp 1636968456
transform 1 0 30268 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_329
timestamp 1
transform 1 0 31372 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_335
timestamp 1
transform 1 0 31924 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_337
timestamp 1636968456
transform 1 0 32108 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_349
timestamp 1636968456
transform 1 0 33212 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_361
timestamp 1636968456
transform 1 0 34316 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_373
timestamp 1636968456
transform 1 0 35420 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_385
timestamp 1
transform 1 0 36524 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_391
timestamp 1
transform 1 0 37076 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_393
timestamp 1636968456
transform 1 0 37260 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_405
timestamp 1636968456
transform 1 0 38364 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_417
timestamp 1636968456
transform 1 0 39468 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_429
timestamp 1636968456
transform 1 0 40572 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_441
timestamp 1
transform 1 0 41676 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_447
timestamp 1
transform 1 0 42228 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_449
timestamp 1636968456
transform 1 0 42412 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_461
timestamp 1636968456
transform 1 0 43516 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_473
timestamp 1636968456
transform 1 0 44620 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_485
timestamp 1636968456
transform 1 0 45724 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_497
timestamp 1
transform 1 0 46828 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_503
timestamp 1
transform 1 0 47380 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_505
timestamp 1636968456
transform 1 0 47564 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_517
timestamp 1636968456
transform 1 0 48668 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_529
timestamp 1636968456
transform 1 0 49772 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_541
timestamp 1636968456
transform 1 0 50876 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_553
timestamp 1
transform 1 0 51980 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_559
timestamp 1
transform 1 0 52532 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_561
timestamp 1636968456
transform 1 0 52716 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_573
timestamp 1636968456
transform 1 0 53820 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_137_585
timestamp 1
transform 1 0 54924 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_588
timestamp 1636968456
transform 1 0 55200 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_600
timestamp 1636968456
transform 1 0 56304 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_612
timestamp 1
transform 1 0 57408 0 -1 77248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_137_617
timestamp 1636968456
transform 1 0 57868 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_629
timestamp 1636968456
transform 1 0 58972 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_641
timestamp 1636968456
transform 1 0 60076 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_653
timestamp 1636968456
transform 1 0 61180 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_665
timestamp 1
transform 1 0 62284 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_671
timestamp 1
transform 1 0 62836 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_673
timestamp 1636968456
transform 1 0 63020 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_685
timestamp 1636968456
transform 1 0 64124 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_697
timestamp 1636968456
transform 1 0 65228 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_709
timestamp 1636968456
transform 1 0 66332 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_721
timestamp 1
transform 1 0 67436 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_727
timestamp 1
transform 1 0 67988 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_729
timestamp 1636968456
transform 1 0 68172 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_741
timestamp 1636968456
transform 1 0 69276 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_753
timestamp 1636968456
transform 1 0 70380 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_765
timestamp 1636968456
transform 1 0 71484 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_777
timestamp 1
transform 1 0 72588 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_783
timestamp 1
transform 1 0 73140 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_785
timestamp 1636968456
transform 1 0 73324 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_797
timestamp 1636968456
transform 1 0 74428 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_809
timestamp 1636968456
transform 1 0 75532 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_821
timestamp 1636968456
transform 1 0 76636 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_833
timestamp 1
transform 1 0 77740 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_839
timestamp 1
transform 1 0 78292 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_841
timestamp 1636968456
transform 1 0 78476 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_853
timestamp 1636968456
transform 1 0 79580 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_865
timestamp 1636968456
transform 1 0 80684 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_877
timestamp 1636968456
transform 1 0 81788 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_889
timestamp 1
transform 1 0 82892 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_895
timestamp 1
transform 1 0 83444 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_897
timestamp 1636968456
transform 1 0 83628 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_909
timestamp 1636968456
transform 1 0 84732 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_921
timestamp 1636968456
transform 1 0 85836 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_933
timestamp 1636968456
transform 1 0 86940 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_945
timestamp 1
transform 1 0 88044 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_949
timestamp 1
transform 1 0 88412 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_137_964
timestamp 1
transform 1 0 89792 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_137_973
timestamp 1
transform 1 0 90620 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_137_990
timestamp 1
transform 1 0 92184 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_137_1002
timestamp 1
transform 1 0 93288 0 -1 77248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1014
timestamp 1636968456
transform 1 0 94392 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_1026
timestamp 1
transform 1 0 95496 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1051
timestamp 1636968456
transform 1 0 97796 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1063
timestamp 1
transform 1 0 98900 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_1071
timestamp 1
transform 1 0 99636 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1079
timestamp 1
transform 1 0 100372 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1083
timestamp 1636968456
transform 1 0 100740 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1095
timestamp 1636968456
transform 1 0 101844 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1107
timestamp 1636968456
transform 1 0 102948 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1119
timestamp 1
transform 1 0 104052 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1121
timestamp 1636968456
transform 1 0 104236 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1133
timestamp 1636968456
transform 1 0 105340 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1145
timestamp 1636968456
transform 1 0 106444 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_1157
timestamp 1
transform 1 0 107548 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1163
timestamp 1
transform 1 0 108100 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636968456
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636968456
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1636968456
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_41
timestamp 1636968456
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_53
timestamp 1
transform 1 0 5980 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_57
timestamp 1636968456
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_69
timestamp 1636968456
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_85
timestamp 1636968456
transform 1 0 8924 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_97
timestamp 1636968456
transform 1 0 10028 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_109
timestamp 1
transform 1 0 11132 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_113
timestamp 1636968456
transform 1 0 11500 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_125
timestamp 1636968456
transform 1 0 12604 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_137
timestamp 1
transform 1 0 13708 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_141
timestamp 1
transform 1 0 14076 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_145
timestamp 1
transform 1 0 14444 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_171
timestamp 1636968456
transform 1 0 16836 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_183
timestamp 1636968456
transform 1 0 17940 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_195
timestamp 1
transform 1 0 19044 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_197
timestamp 1636968456
transform 1 0 19228 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_209
timestamp 1636968456
transform 1 0 20332 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_221
timestamp 1
transform 1 0 21436 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_225
timestamp 1636968456
transform 1 0 21804 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_237
timestamp 1
transform 1 0 22908 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_138_245
timestamp 1
transform 1 0 23644 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_249
timestamp 1
transform 1 0 24012 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_273
timestamp 1
transform 1 0 26220 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_279
timestamp 1
transform 1 0 26772 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_283
timestamp 1
transform 1 0 27140 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_291
timestamp 1
transform 1 0 27876 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_296
timestamp 1636968456
transform 1 0 28336 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_311
timestamp 1
transform 1 0 29716 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_138_321
timestamp 1
transform 1 0 30636 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_329
timestamp 1
transform 1 0 31372 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_138_334
timestamp 1
transform 1 0 31832 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_138_337
timestamp 1
transform 1 0 32108 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_138_347
timestamp 1
transform 1 0 33028 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_138_355
timestamp 1
transform 1 0 33764 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_138_359
timestamp 1
transform 1 0 34132 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_363
timestamp 1
transform 1 0 34500 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_138_365
timestamp 1
transform 1 0 34684 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_369
timestamp 1
transform 1 0 35052 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_372
timestamp 1
transform 1 0 35328 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_380
timestamp 1
transform 1 0 36064 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_138_385
timestamp 1
transform 1 0 36524 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_391
timestamp 1
transform 1 0 37076 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_138_393
timestamp 1
transform 1 0 37260 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_138_397
timestamp 1
transform 1 0 37628 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_405
timestamp 1
transform 1 0 38364 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_138_410
timestamp 1
transform 1 0 38824 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_138_418
timestamp 1
transform 1 0 39560 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_138_423
timestamp 1
transform 1 0 40020 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_431
timestamp 1
transform 1 0 40756 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_138_436
timestamp 1
transform 1 0 41216 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_138_444
timestamp 1
transform 1 0 41952 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_138_449
timestamp 1
transform 1 0 42412 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_138_457
timestamp 1
transform 1 0 43148 0 1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_138_461
timestamp 1636968456
transform 1 0 43516 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_473
timestamp 1
transform 1 0 44620 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_477
timestamp 1636968456
transform 1 0 44988 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_489
timestamp 1636968456
transform 1 0 46092 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_501
timestamp 1
transform 1 0 47196 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_505
timestamp 1636968456
transform 1 0 47564 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_517
timestamp 1636968456
transform 1 0 48668 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_529
timestamp 1
transform 1 0 49772 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_533
timestamp 1636968456
transform 1 0 50140 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_545
timestamp 1636968456
transform 1 0 51244 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_557
timestamp 1
transform 1 0 52348 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_561
timestamp 1636968456
transform 1 0 52716 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_573
timestamp 1
transform 1 0 53820 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_579
timestamp 1
transform 1 0 54372 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_138_611
timestamp 1
transform 1 0 57316 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_615
timestamp 1
transform 1 0 57684 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_617
timestamp 1636968456
transform 1 0 57868 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_629
timestamp 1636968456
transform 1 0 58972 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_641
timestamp 1
transform 1 0 60076 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_645
timestamp 1636968456
transform 1 0 60444 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_657
timestamp 1636968456
transform 1 0 61548 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_669
timestamp 1
transform 1 0 62652 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_673
timestamp 1636968456
transform 1 0 63020 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_685
timestamp 1636968456
transform 1 0 64124 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_697
timestamp 1
transform 1 0 65228 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_701
timestamp 1636968456
transform 1 0 65596 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_713
timestamp 1636968456
transform 1 0 66700 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_725
timestamp 1
transform 1 0 67804 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_729
timestamp 1636968456
transform 1 0 68172 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_741
timestamp 1636968456
transform 1 0 69276 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_753
timestamp 1
transform 1 0 70380 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_757
timestamp 1636968456
transform 1 0 70748 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_769
timestamp 1636968456
transform 1 0 71852 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_781
timestamp 1
transform 1 0 72956 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_785
timestamp 1636968456
transform 1 0 73324 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_797
timestamp 1636968456
transform 1 0 74428 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_809
timestamp 1
transform 1 0 75532 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_813
timestamp 1636968456
transform 1 0 75900 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_825
timestamp 1636968456
transform 1 0 77004 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_837
timestamp 1
transform 1 0 78108 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_841
timestamp 1636968456
transform 1 0 78476 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_853
timestamp 1636968456
transform 1 0 79580 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_865
timestamp 1
transform 1 0 80684 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_869
timestamp 1636968456
transform 1 0 81052 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_881
timestamp 1636968456
transform 1 0 82156 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_893
timestamp 1
transform 1 0 83260 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_908
timestamp 1636968456
transform 1 0 84640 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_138_920
timestamp 1
transform 1 0 85744 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_138_925
timestamp 1
transform 1 0 86204 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_937
timestamp 1636968456
transform 1 0 87308 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_949
timestamp 1
transform 1 0 88412 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_138_953
timestamp 1
transform 1 0 88780 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_987
timestamp 1
transform 1 0 91908 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1009
timestamp 1
transform 1 0 93932 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1024
timestamp 1636968456
transform 1 0 95312 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_1037
timestamp 1
transform 1 0 96508 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1043
timestamp 1
transform 1 0 97060 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1067
timestamp 1636968456
transform 1 0 99268 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1079
timestamp 1636968456
transform 1 0 100372 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1091
timestamp 1
transform 1 0 101476 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1093
timestamp 1636968456
transform 1 0 101660 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1105
timestamp 1636968456
transform 1 0 102764 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_1117
timestamp 1
transform 1 0 103868 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1121
timestamp 1636968456
transform 1 0 104236 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1133
timestamp 1636968456
transform 1 0 105340 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_1145
timestamp 1
transform 1 0 106444 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1149
timestamp 1636968456
transform 1 0 106812 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_1161
timestamp 1
transform 1 0 107916 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1167
timestamp 1
transform 1 0 108468 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_11
timestamp 1636968456
transform 1 0 2116 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_23
timestamp 1636968456
transform 1 0 3220 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_35
timestamp 1636968456
transform 1 0 4324 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_47
timestamp 1
transform 1 0 5428 0 -1 78336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_139_55
timestamp 1
transform 1 0 6164 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_57
timestamp 1636968456
transform 1 0 6348 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_139_69
timestamp 1
transform 1 0 7452 0 -1 78336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1122
timestamp 1636968456
transform 1 0 104328 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1134
timestamp 1636968456
transform 1 0 105432 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1146
timestamp 1636968456
transform 1 0 106536 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_1158
timestamp 1
transform 1 0 107640 0 -1 78336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_140_11
timestamp 1636968456
transform 1 0 2116 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_140_23
timestamp 1
transform 1 0 3220 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 1
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_29
timestamp 1636968456
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_41
timestamp 1636968456
transform 1 0 4876 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_53
timestamp 1636968456
transform 1 0 5980 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_65
timestamp 1
transform 1 0 7084 0 1 78336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1122
timestamp 1636968456
transform 1 0 104328 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1134
timestamp 1636968456
transform 1 0 105432 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_1146
timestamp 1
transform 1 0 106536 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1148
timestamp 1636968456
transform 1 0 106720 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_140_1160
timestamp 1
transform 1 0 107824 0 1 78336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_141_11
timestamp 1636968456
transform 1 0 2116 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_23
timestamp 1636968456
transform 1 0 3220 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_35
timestamp 1636968456
transform 1 0 4324 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_47
timestamp 1
transform 1 0 5428 0 -1 79424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_141_55
timestamp 1
transform 1 0 6164 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_57
timestamp 1636968456
transform 1 0 6348 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_141_69
timestamp 1
transform 1 0 7452 0 -1 79424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1122
timestamp 1636968456
transform 1 0 104328 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1134
timestamp 1636968456
transform 1 0 105432 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1146
timestamp 1636968456
transform 1 0 106536 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_1158
timestamp 1
transform 1 0 107640 0 -1 79424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_142_11
timestamp 1636968456
transform 1 0 2116 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_142_23
timestamp 1
transform 1 0 3220 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 1
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_29
timestamp 1636968456
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_41
timestamp 1636968456
transform 1 0 4876 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_53
timestamp 1636968456
transform 1 0 5980 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_65
timestamp 1
transform 1 0 7084 0 1 79424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1122
timestamp 1636968456
transform 1 0 104328 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1134
timestamp 1636968456
transform 1 0 105432 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_1146
timestamp 1
transform 1 0 106536 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1148
timestamp 1636968456
transform 1 0 106720 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_142_1160
timestamp 1
transform 1 0 107824 0 1 79424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_143_5
timestamp 1636968456
transform 1 0 1564 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_17
timestamp 1636968456
transform 1 0 2668 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_29
timestamp 1636968456
transform 1 0 3772 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_41
timestamp 1636968456
transform 1 0 4876 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_143_53
timestamp 1
transform 1 0 5980 0 -1 80512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_143_57
timestamp 1636968456
transform 1 0 6348 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_143_69
timestamp 1
transform 1 0 7452 0 -1 80512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1122
timestamp 1636968456
transform 1 0 104328 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1134
timestamp 1636968456
transform 1 0 105432 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1146
timestamp 1636968456
transform 1 0 106536 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_1158
timestamp 1
transform 1 0 107640 0 -1 80512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636968456
transform 1 0 2484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 1
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_29
timestamp 1636968456
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_41
timestamp 1636968456
transform 1 0 4876 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_53
timestamp 1636968456
transform 1 0 5980 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_65
timestamp 1
transform 1 0 7084 0 1 80512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1122
timestamp 1636968456
transform 1 0 104328 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1134
timestamp 1636968456
transform 1 0 105432 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_1146
timestamp 1
transform 1 0 106536 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_144_1148
timestamp 1
transform 1 0 106720 0 1 80512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_144_1156
timestamp 1
transform 1 0 107456 0 1 80512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_145_11
timestamp 1636968456
transform 1 0 2116 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_23
timestamp 1636968456
transform 1 0 3220 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_35
timestamp 1636968456
transform 1 0 4324 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_47
timestamp 1
transform 1 0 5428 0 -1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_145_55
timestamp 1
transform 1 0 6164 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_57
timestamp 1636968456
transform 1 0 6348 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_145_69
timestamp 1
transform 1 0 7452 0 -1 81600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1122
timestamp 1636968456
transform 1 0 104328 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1134
timestamp 1636968456
transform 1 0 105432 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1146
timestamp 1636968456
transform 1 0 106536 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_1158
timestamp 1
transform 1 0 107640 0 -1 81600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_145_1166
timestamp 1
transform 1 0 108376 0 -1 81600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_11
timestamp 1636968456
transform 1 0 2116 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_146_23
timestamp 1
transform 1 0 3220 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 1
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636968456
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_41
timestamp 1636968456
transform 1 0 4876 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_53
timestamp 1636968456
transform 1 0 5980 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_65
timestamp 1
transform 1 0 7084 0 1 81600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1122
timestamp 1636968456
transform 1 0 104328 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1134
timestamp 1636968456
transform 1 0 105432 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_1146
timestamp 1
transform 1 0 106536 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1148
timestamp 1636968456
transform 1 0 106720 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_1160
timestamp 1
transform 1 0 107824 0 1 81600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_147_11
timestamp 1636968456
transform 1 0 2116 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_23
timestamp 1
transform 1 0 3220 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_147_31
timestamp 1
transform 1 0 3956 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_147_47
timestamp 1
transform 1 0 5428 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_147_55
timestamp 1
transform 1 0 6164 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_57
timestamp 1636968456
transform 1 0 6348 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_147_69
timestamp 1
transform 1 0 7452 0 -1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1122
timestamp 1636968456
transform 1 0 104328 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1134
timestamp 1636968456
transform 1 0 105432 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1146
timestamp 1636968456
transform 1 0 106536 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_1158
timestamp 1
transform 1 0 107640 0 -1 82688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_147_1166
timestamp 1
transform 1 0 108376 0 -1 82688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636968456
transform 1 0 1380 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636968456
transform 1 0 2484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 1
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636968456
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_41
timestamp 1636968456
transform 1 0 4876 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_53
timestamp 1636968456
transform 1 0 5980 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_65
timestamp 1
transform 1 0 7084 0 1 82688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1122
timestamp 1636968456
transform 1 0 104328 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1134
timestamp 1636968456
transform 1 0 105432 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_1146
timestamp 1
transform 1 0 106536 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1148
timestamp 1636968456
transform 1 0 106720 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_1160
timestamp 1
transform 1 0 107824 0 1 82688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_149_11
timestamp 1636968456
transform 1 0 2116 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_23
timestamp 1636968456
transform 1 0 3220 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_35
timestamp 1636968456
transform 1 0 4324 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_47
timestamp 1
transform 1 0 5428 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_149_55
timestamp 1
transform 1 0 6164 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_57
timestamp 1636968456
transform 1 0 6348 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_149_69
timestamp 1
transform 1 0 7452 0 -1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1122
timestamp 1636968456
transform 1 0 104328 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1134
timestamp 1636968456
transform 1 0 105432 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1146
timestamp 1636968456
transform 1 0 106536 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_1158
timestamp 1
transform 1 0 107640 0 -1 83776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_149_1166
timestamp 1
transform 1 0 108376 0 -1 83776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_150_11
timestamp 1636968456
transform 1 0 2116 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_150_23
timestamp 1
transform 1 0 3220 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 1
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636968456
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_41
timestamp 1636968456
transform 1 0 4876 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_53
timestamp 1636968456
transform 1 0 5980 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_65
timestamp 1
transform 1 0 7084 0 1 83776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1122
timestamp 1636968456
transform 1 0 104328 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1134
timestamp 1636968456
transform 1 0 105432 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_1146
timestamp 1
transform 1 0 106536 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1148
timestamp 1636968456
transform 1 0 106720 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_1160
timestamp 1
transform 1 0 107824 0 1 83776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_151_11
timestamp 1636968456
transform 1 0 2116 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_23
timestamp 1636968456
transform 1 0 3220 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_35
timestamp 1636968456
transform 1 0 4324 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_47
timestamp 1
transform 1 0 5428 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_55
timestamp 1
transform 1 0 6164 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_57
timestamp 1636968456
transform 1 0 6348 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_151_69
timestamp 1
transform 1 0 7452 0 -1 84864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1122
timestamp 1636968456
transform 1 0 104328 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1134
timestamp 1636968456
transform 1 0 105432 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1146
timestamp 1636968456
transform 1 0 106536 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_1158
timestamp 1
transform 1 0 107640 0 -1 84864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_151_1166
timestamp 1
transform 1 0 108376 0 -1 84864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_152_11
timestamp 1636968456
transform 1 0 2116 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_152_23
timestamp 1
transform 1 0 3220 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 1
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_29
timestamp 1636968456
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_41
timestamp 1636968456
transform 1 0 4876 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_53
timestamp 1636968456
transform 1 0 5980 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_65
timestamp 1
transform 1 0 7084 0 1 84864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1122
timestamp 1636968456
transform 1 0 104328 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1134
timestamp 1636968456
transform 1 0 105432 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_1146
timestamp 1
transform 1 0 106536 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1148
timestamp 1636968456
transform 1 0 106720 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_1160
timestamp 1
transform 1 0 107824 0 1 84864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_153_3
timestamp 1636968456
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_15
timestamp 1636968456
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_27
timestamp 1636968456
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_39
timestamp 1636968456
transform 1 0 4692 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_51
timestamp 1
transform 1 0 5796 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_55
timestamp 1
transform 1 0 6164 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_57
timestamp 1636968456
transform 1 0 6348 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_153_69
timestamp 1
transform 1 0 7452 0 -1 85952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1122
timestamp 1636968456
transform 1 0 104328 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1134
timestamp 1636968456
transform 1 0 105432 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1146
timestamp 1636968456
transform 1 0 106536 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_1158
timestamp 1
transform 1 0 107640 0 -1 85952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_153_1166
timestamp 1
transform 1 0 108376 0 -1 85952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_154_8
timestamp 1636968456
transform 1 0 1840 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_20
timestamp 1
transform 1 0 2944 0 1 85952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_154_29
timestamp 1636968456
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_41
timestamp 1636968456
transform 1 0 4876 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_53
timestamp 1636968456
transform 1 0 5980 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_65
timestamp 1
transform 1 0 7084 0 1 85952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1122
timestamp 1636968456
transform 1 0 104328 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1134
timestamp 1636968456
transform 1 0 105432 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_1146
timestamp 1
transform 1 0 106536 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1148
timestamp 1636968456
transform 1 0 106720 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_1160
timestamp 1
transform 1 0 107824 0 1 85952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_155_11
timestamp 1636968456
transform 1 0 2116 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_23
timestamp 1636968456
transform 1 0 3220 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_35
timestamp 1636968456
transform 1 0 4324 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_47
timestamp 1
transform 1 0 5428 0 -1 87040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_155_55
timestamp 1
transform 1 0 6164 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_57
timestamp 1636968456
transform 1 0 6348 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_155_69
timestamp 1
transform 1 0 7452 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1122
timestamp 1636968456
transform 1 0 104328 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1134
timestamp 1636968456
transform 1 0 105432 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1146
timestamp 1636968456
transform 1 0 106536 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_1158
timestamp 1
transform 1 0 107640 0 -1 87040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_155_1166
timestamp 1
transform 1 0 108376 0 -1 87040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_156_11
timestamp 1636968456
transform 1 0 2116 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_156_23
timestamp 1
transform 1 0 3220 0 1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_156_27
timestamp 1
transform 1 0 3588 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_29
timestamp 1636968456
transform 1 0 3772 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_41
timestamp 1636968456
transform 1 0 4876 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_53
timestamp 1636968456
transform 1 0 5980 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_65
timestamp 1
transform 1 0 7084 0 1 87040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1122
timestamp 1636968456
transform 1 0 104328 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1134
timestamp 1636968456
transform 1 0 105432 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_1146
timestamp 1
transform 1 0 106536 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1148
timestamp 1636968456
transform 1 0 106720 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_1160
timestamp 1
transform 1 0 107824 0 1 87040
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_157_11
timestamp 1636968456
transform 1 0 2116 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_23
timestamp 1636968456
transform 1 0 3220 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_35
timestamp 1636968456
transform 1 0 4324 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_47
timestamp 1
transform 1 0 5428 0 -1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_157_55
timestamp 1
transform 1 0 6164 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_57
timestamp 1636968456
transform 1 0 6348 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_157_69
timestamp 1
transform 1 0 7452 0 -1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1122
timestamp 1636968456
transform 1 0 104328 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1134
timestamp 1636968456
transform 1 0 105432 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1146
timestamp 1636968456
transform 1 0 106536 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_1158
timestamp 1
transform 1 0 107640 0 -1 88128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_157_1166
timestamp 1
transform 1 0 108376 0 -1 88128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_158_3
timestamp 1636968456
transform 1 0 1380 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_15
timestamp 1636968456
transform 1 0 2484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_27
timestamp 1
transform 1 0 3588 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_29
timestamp 1636968456
transform 1 0 3772 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_41
timestamp 1636968456
transform 1 0 4876 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_53
timestamp 1636968456
transform 1 0 5980 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_65
timestamp 1
transform 1 0 7084 0 1 88128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1122
timestamp 1636968456
transform 1 0 104328 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1134
timestamp 1636968456
transform 1 0 105432 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_1146
timestamp 1
transform 1 0 106536 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1148
timestamp 1636968456
transform 1 0 106720 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_1160
timestamp 1
transform 1 0 107824 0 1 88128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_159_11
timestamp 1636968456
transform 1 0 2116 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_23
timestamp 1636968456
transform 1 0 3220 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_35
timestamp 1636968456
transform 1 0 4324 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_47
timestamp 1
transform 1 0 5428 0 -1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_159_55
timestamp 1
transform 1 0 6164 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_57
timestamp 1636968456
transform 1 0 6348 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_159_69
timestamp 1
transform 1 0 7452 0 -1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1122
timestamp 1636968456
transform 1 0 104328 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1134
timestamp 1636968456
transform 1 0 105432 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1146
timestamp 1636968456
transform 1 0 106536 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_1158
timestamp 1
transform 1 0 107640 0 -1 89216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_159_1166
timestamp 1
transform 1 0 108376 0 -1 89216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_160_3
timestamp 1636968456
transform 1 0 1380 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_15
timestamp 1636968456
transform 1 0 2484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_27
timestamp 1
transform 1 0 3588 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_29
timestamp 1636968456
transform 1 0 3772 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_41
timestamp 1636968456
transform 1 0 4876 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_53
timestamp 1636968456
transform 1 0 5980 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_65
timestamp 1
transform 1 0 7084 0 1 89216
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1122
timestamp 1636968456
transform 1 0 104328 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1134
timestamp 1636968456
transform 1 0 105432 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_1146
timestamp 1
transform 1 0 106536 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1148
timestamp 1636968456
transform 1 0 106720 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_160_1160
timestamp 1
transform 1 0 107824 0 1 89216
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_161_3
timestamp 1636968456
transform 1 0 1380 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_15
timestamp 1636968456
transform 1 0 2484 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_27
timestamp 1636968456
transform 1 0 3588 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_39
timestamp 1636968456
transform 1 0 4692 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_161_51
timestamp 1
transform 1 0 5796 0 -1 90304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_161_55
timestamp 1
transform 1 0 6164 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_57
timestamp 1636968456
transform 1 0 6348 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_161_69
timestamp 1
transform 1 0 7452 0 -1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1122
timestamp 1636968456
transform 1 0 104328 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1134
timestamp 1636968456
transform 1 0 105432 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1146
timestamp 1636968456
transform 1 0 106536 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_1158
timestamp 1
transform 1 0 107640 0 -1 90304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_161_1166
timestamp 1
transform 1 0 108376 0 -1 90304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_162_3
timestamp 1636968456
transform 1 0 1380 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_15
timestamp 1636968456
transform 1 0 2484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_27
timestamp 1
transform 1 0 3588 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_29
timestamp 1636968456
transform 1 0 3772 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_41
timestamp 1636968456
transform 1 0 4876 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_53
timestamp 1636968456
transform 1 0 5980 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_65
timestamp 1
transform 1 0 7084 0 1 90304
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1122
timestamp 1636968456
transform 1 0 104328 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1134
timestamp 1636968456
transform 1 0 105432 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_1146
timestamp 1
transform 1 0 106536 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1148
timestamp 1636968456
transform 1 0 106720 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_1160
timestamp 1
transform 1 0 107824 0 1 90304
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_163_3
timestamp 1636968456
transform 1 0 1380 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_15
timestamp 1636968456
transform 1 0 2484 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_27
timestamp 1636968456
transform 1 0 3588 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_39
timestamp 1636968456
transform 1 0 4692 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_163_51
timestamp 1
transform 1 0 5796 0 -1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_163_55
timestamp 1
transform 1 0 6164 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_57
timestamp 1636968456
transform 1 0 6348 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_163_69
timestamp 1
transform 1 0 7452 0 -1 91392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1124
timestamp 1636968456
transform 1 0 104512 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1136
timestamp 1636968456
transform 1 0 105616 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1148
timestamp 1636968456
transform 1 0 106720 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_1160
timestamp 1
transform 1 0 107824 0 -1 91392
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_164_3
timestamp 1636968456
transform 1 0 1380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_15
timestamp 1636968456
transform 1 0 2484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_27
timestamp 1
transform 1 0 3588 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_29
timestamp 1636968456
transform 1 0 3772 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_41
timestamp 1636968456
transform 1 0 4876 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_53
timestamp 1636968456
transform 1 0 5980 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_65
timestamp 1
transform 1 0 7084 0 1 91392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1135
timestamp 1636968456
transform 1 0 105524 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1148
timestamp 1636968456
transform 1 0 106720 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_1160
timestamp 1
transform 1 0 107824 0 1 91392
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_165_3
timestamp 1636968456
transform 1 0 1380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_15
timestamp 1636968456
transform 1 0 2484 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_27
timestamp 1636968456
transform 1 0 3588 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_39
timestamp 1636968456
transform 1 0 4692 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_51
timestamp 1
transform 1 0 5796 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_165_55
timestamp 1
transform 1 0 6164 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_57
timestamp 1636968456
transform 1 0 6348 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_165_69
timestamp 1
transform 1 0 7452 0 -1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1122
timestamp 1636968456
transform 1 0 104328 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1134
timestamp 1636968456
transform 1 0 105432 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1146
timestamp 1636968456
transform 1 0 106536 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_1158
timestamp 1
transform 1 0 107640 0 -1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_165_1166
timestamp 1
transform 1 0 108376 0 -1 92480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_166_3
timestamp 1636968456
transform 1 0 1380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_15
timestamp 1636968456
transform 1 0 2484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_27
timestamp 1
transform 1 0 3588 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_29
timestamp 1636968456
transform 1 0 3772 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_41
timestamp 1636968456
transform 1 0 4876 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_53
timestamp 1636968456
transform 1 0 5980 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_65
timestamp 1
transform 1 0 7084 0 1 92480
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1124
timestamp 1636968456
transform 1 0 104512 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_1136
timestamp 1
transform 1 0 105616 0 1 92480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_166_1144
timestamp 1
transform 1 0 106352 0 1 92480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1148
timestamp 1636968456
transform 1 0 106720 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_1160
timestamp 1
transform 1 0 107824 0 1 92480
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_167_3
timestamp 1636968456
transform 1 0 1380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_15
timestamp 1636968456
transform 1 0 2484 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_27
timestamp 1636968456
transform 1 0 3588 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_39
timestamp 1636968456
transform 1 0 4692 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_51
timestamp 1
transform 1 0 5796 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_55
timestamp 1
transform 1 0 6164 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_57
timestamp 1
transform 1 0 6348 0 -1 93568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1122
timestamp 1636968456
transform 1 0 104328 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1134
timestamp 1636968456
transform 1 0 105432 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1146
timestamp 1636968456
transform 1 0 106536 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_1158
timestamp 1
transform 1 0 107640 0 -1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_167_1166
timestamp 1
transform 1 0 108376 0 -1 93568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_168_3
timestamp 1636968456
transform 1 0 1380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_15
timestamp 1636968456
transform 1 0 2484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_27
timestamp 1
transform 1 0 3588 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_29
timestamp 1636968456
transform 1 0 3772 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_41
timestamp 1636968456
transform 1 0 4876 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_168_53
timestamp 1
transform 1 0 5980 0 1 93568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1124
timestamp 1636968456
transform 1 0 104512 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_1136
timestamp 1
transform 1 0 105616 0 1 93568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_168_1144
timestamp 1
transform 1 0 106352 0 1 93568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1148
timestamp 1636968456
transform 1 0 106720 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_1160
timestamp 1
transform 1 0 107824 0 1 93568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_169_3
timestamp 1636968456
transform 1 0 1380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_15
timestamp 1636968456
transform 1 0 2484 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_27
timestamp 1636968456
transform 1 0 3588 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_39
timestamp 1636968456
transform 1 0 4692 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_51
timestamp 1
transform 1 0 5796 0 -1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_169_55
timestamp 1
transform 1 0 6164 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_169_57
timestamp 1
transform 1 0 6348 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1122
timestamp 1636968456
transform 1 0 104328 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1134
timestamp 1636968456
transform 1 0 105432 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1146
timestamp 1636968456
transform 1 0 106536 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_1158
timestamp 1
transform 1 0 107640 0 -1 94656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_169_1166
timestamp 1
transform 1 0 108376 0 -1 94656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_170_3
timestamp 1636968456
transform 1 0 1380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_15
timestamp 1636968456
transform 1 0 2484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_27
timestamp 1
transform 1 0 3588 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_29
timestamp 1636968456
transform 1 0 3772 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_41
timestamp 1
transform 1 0 4876 0 1 94656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1122
timestamp 1636968456
transform 1 0 104328 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1134
timestamp 1636968456
transform 1 0 105432 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1146
timestamp 1
transform 1 0 106536 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1148
timestamp 1636968456
transform 1 0 106720 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_1160
timestamp 1
transform 1 0 107824 0 1 94656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_171_3
timestamp 1636968456
transform 1 0 1380 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_15
timestamp 1636968456
transform 1 0 2484 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_27
timestamp 1636968456
transform 1 0 3588 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_39
timestamp 1636968456
transform 1 0 4692 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_171_51
timestamp 1
transform 1 0 5796 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_55
timestamp 1
transform 1 0 6164 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_57
timestamp 1636968456
transform 1 0 6348 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1124
timestamp 1636968456
transform 1 0 104512 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1136
timestamp 1636968456
transform 1 0 105616 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1148
timestamp 1636968456
transform 1 0 106720 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_1160
timestamp 1
transform 1 0 107824 0 -1 95744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_172_3
timestamp 1636968456
transform 1 0 1380 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_15
timestamp 1636968456
transform 1 0 2484 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_27
timestamp 1
transform 1 0 3588 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_29
timestamp 1636968456
transform 1 0 3772 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_41
timestamp 1636968456
transform 1 0 4876 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_53
timestamp 1636968456
transform 1 0 5980 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_65
timestamp 1
transform 1 0 7084 0 1 95744
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1124
timestamp 1636968456
transform 1 0 104512 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_1136
timestamp 1
transform 1 0 105616 0 1 95744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_172_1144
timestamp 1
transform 1 0 106352 0 1 95744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1148
timestamp 1636968456
transform 1 0 106720 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_1160
timestamp 1
transform 1 0 107824 0 1 95744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_173_3
timestamp 1636968456
transform 1 0 1380 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_15
timestamp 1636968456
transform 1 0 2484 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_27
timestamp 1636968456
transform 1 0 3588 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_39
timestamp 1636968456
transform 1 0 4692 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_173_51
timestamp 1
transform 1 0 5796 0 -1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_173_55
timestamp 1
transform 1 0 6164 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_57
timestamp 1636968456
transform 1 0 6348 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_173_69
timestamp 1
transform 1 0 7452 0 -1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1142
timestamp 1636968456
transform 1 0 106168 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1154
timestamp 1636968456
transform 1 0 107272 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_173_1166
timestamp 1
transform 1 0 108376 0 -1 96832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_174_3
timestamp 1636968456
transform 1 0 1380 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_15
timestamp 1636968456
transform 1 0 2484 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_174_27
timestamp 1
transform 1 0 3588 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_29
timestamp 1636968456
transform 1 0 3772 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_41
timestamp 1636968456
transform 1 0 4876 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_53
timestamp 1636968456
transform 1 0 5980 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_65
timestamp 1
transform 1 0 7084 0 1 96832
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1122
timestamp 1636968456
transform 1 0 104328 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1134
timestamp 1636968456
transform 1 0 105432 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_174_1146
timestamp 1
transform 1 0 106536 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1148
timestamp 1636968456
transform 1 0 106720 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_174_1160
timestamp 1
transform 1 0 107824 0 1 96832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_175_3
timestamp 1636968456
transform 1 0 1380 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_15
timestamp 1636968456
transform 1 0 2484 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_27
timestamp 1636968456
transform 1 0 3588 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_39
timestamp 1636968456
transform 1 0 4692 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_175_51
timestamp 1
transform 1 0 5796 0 -1 97920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_175_55
timestamp 1
transform 1 0 6164 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_57
timestamp 1636968456
transform 1 0 6348 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_175_69
timestamp 1
transform 1 0 7452 0 -1 97920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1122
timestamp 1636968456
transform 1 0 104328 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1134
timestamp 1636968456
transform 1 0 105432 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1146
timestamp 1636968456
transform 1 0 106536 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_1158
timestamp 1
transform 1 0 107640 0 -1 97920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_175_1166
timestamp 1
transform 1 0 108376 0 -1 97920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_176_3
timestamp 1636968456
transform 1 0 1380 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_15
timestamp 1636968456
transform 1 0 2484 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_27
timestamp 1
transform 1 0 3588 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_29
timestamp 1636968456
transform 1 0 3772 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_41
timestamp 1636968456
transform 1 0 4876 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_53
timestamp 1636968456
transform 1 0 5980 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_65
timestamp 1
transform 1 0 7084 0 1 97920
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1122
timestamp 1636968456
transform 1 0 104328 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1134
timestamp 1636968456
transform 1 0 105432 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_1146
timestamp 1
transform 1 0 106536 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1148
timestamp 1636968456
transform 1 0 106720 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_176_1160
timestamp 1
transform 1 0 107824 0 1 97920
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_177_3
timestamp 1636968456
transform 1 0 1380 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_15
timestamp 1636968456
transform 1 0 2484 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_27
timestamp 1636968456
transform 1 0 3588 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_39
timestamp 1636968456
transform 1 0 4692 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_177_51
timestamp 1
transform 1 0 5796 0 -1 99008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_177_55
timestamp 1
transform 1 0 6164 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_57
timestamp 1636968456
transform 1 0 6348 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_177_69
timestamp 1
transform 1 0 7452 0 -1 99008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1122
timestamp 1636968456
transform 1 0 104328 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1134
timestamp 1636968456
transform 1 0 105432 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1146
timestamp 1636968456
transform 1 0 106536 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_1158
timestamp 1
transform 1 0 107640 0 -1 99008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_177_1166
timestamp 1
transform 1 0 108376 0 -1 99008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_178_3
timestamp 1636968456
transform 1 0 1380 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_15
timestamp 1636968456
transform 1 0 2484 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_27
timestamp 1
transform 1 0 3588 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_29
timestamp 1636968456
transform 1 0 3772 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_41
timestamp 1636968456
transform 1 0 4876 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_53
timestamp 1636968456
transform 1 0 5980 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_65
timestamp 1
transform 1 0 7084 0 1 99008
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1122
timestamp 1636968456
transform 1 0 104328 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1134
timestamp 1636968456
transform 1 0 105432 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_1146
timestamp 1
transform 1 0 106536 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1148
timestamp 1636968456
transform 1 0 106720 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_178_1160
timestamp 1
transform 1 0 107824 0 1 99008
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_179_3
timestamp 1636968456
transform 1 0 1380 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_15
timestamp 1636968456
transform 1 0 2484 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_27
timestamp 1636968456
transform 1 0 3588 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_39
timestamp 1636968456
transform 1 0 4692 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_51
timestamp 1
transform 1 0 5796 0 -1 100096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_179_55
timestamp 1
transform 1 0 6164 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_179_57
timestamp 1
transform 1 0 6348 0 -1 100096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_179_65
timestamp 1
transform 1 0 7084 0 -1 100096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1122
timestamp 1636968456
transform 1 0 104328 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1134
timestamp 1636968456
transform 1 0 105432 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1146
timestamp 1636968456
transform 1 0 106536 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_1158
timestamp 1
transform 1 0 107640 0 -1 100096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_179_1166
timestamp 1
transform 1 0 108376 0 -1 100096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_180_3
timestamp 1636968456
transform 1 0 1380 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_15
timestamp 1636968456
transform 1 0 2484 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_180_27
timestamp 1
transform 1 0 3588 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_29
timestamp 1636968456
transform 1 0 3772 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_41
timestamp 1636968456
transform 1 0 4876 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_180_53
timestamp 1
transform 1 0 5980 0 1 100096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1124
timestamp 1636968456
transform 1 0 104512 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_180_1136
timestamp 1
transform 1 0 105616 0 1 100096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_180_1144
timestamp 1
transform 1 0 106352 0 1 100096
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1148
timestamp 1636968456
transform 1 0 106720 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_180_1160
timestamp 1
transform 1 0 107824 0 1 100096
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_181_3
timestamp 1636968456
transform 1 0 1380 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_15
timestamp 1636968456
transform 1 0 2484 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_27
timestamp 1636968456
transform 1 0 3588 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_39
timestamp 1636968456
transform 1 0 4692 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_181_51
timestamp 1
transform 1 0 5796 0 -1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_181_55
timestamp 1
transform 1 0 6164 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_57
timestamp 1636968456
transform 1 0 6348 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1142
timestamp 1636968456
transform 1 0 106168 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1154
timestamp 1636968456
transform 1 0 107272 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_181_1166
timestamp 1
transform 1 0 108376 0 -1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_182_3
timestamp 1636968456
transform 1 0 1380 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_15
timestamp 1636968456
transform 1 0 2484 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_182_27
timestamp 1
transform 1 0 3588 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_29
timestamp 1636968456
transform 1 0 3772 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_41
timestamp 1636968456
transform 1 0 4876 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_53
timestamp 1636968456
transform 1 0 5980 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_182_65
timestamp 1
transform 1 0 7084 0 1 101184
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1122
timestamp 1636968456
transform 1 0 104328 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1134
timestamp 1636968456
transform 1 0 105432 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_182_1146
timestamp 1
transform 1 0 106536 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1148
timestamp 1636968456
transform 1 0 106720 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_1160
timestamp 1
transform 1 0 107824 0 1 101184
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_183_3
timestamp 1636968456
transform 1 0 1380 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_15
timestamp 1636968456
transform 1 0 2484 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_27
timestamp 1636968456
transform 1 0 3588 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_39
timestamp 1636968456
transform 1 0 4692 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_183_51
timestamp 1
transform 1 0 5796 0 -1 102272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_183_55
timestamp 1
transform 1 0 6164 0 -1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_183_57
timestamp 1636968456
transform 1 0 6348 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_183_69
timestamp 1
transform 1 0 7452 0 -1 102272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1122
timestamp 1636968456
transform 1 0 104328 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1134
timestamp 1636968456
transform 1 0 105432 0 -1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_183_1146
timestamp 1636968456
transform 1 0 106536 0 -1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_1158
timestamp 1
transform 1 0 107640 0 -1 102272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_183_1166
timestamp 1
transform 1 0 108376 0 -1 102272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_184_3
timestamp 1636968456
transform 1 0 1380 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_15
timestamp 1636968456
transform 1 0 2484 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_184_27
timestamp 1
transform 1 0 3588 0 1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_184_29
timestamp 1636968456
transform 1 0 3772 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_41
timestamp 1636968456
transform 1 0 4876 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_53
timestamp 1636968456
transform 1 0 5980 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_184_65
timestamp 1
transform 1 0 7084 0 1 102272
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1122
timestamp 1636968456
transform 1 0 104328 0 1 102272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1134
timestamp 1636968456
transform 1 0 105432 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_184_1146
timestamp 1
transform 1 0 106536 0 1 102272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_184_1148
timestamp 1636968456
transform 1 0 106720 0 1 102272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_184_1160
timestamp 1
transform 1 0 107824 0 1 102272
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_185_3
timestamp 1636968456
transform 1 0 1380 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_15
timestamp 1636968456
transform 1 0 2484 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_27
timestamp 1636968456
transform 1 0 3588 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_39
timestamp 1636968456
transform 1 0 4692 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_185_51
timestamp 1
transform 1 0 5796 0 -1 103360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_185_55
timestamp 1
transform 1 0 6164 0 -1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_185_57
timestamp 1636968456
transform 1 0 6348 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_185_69
timestamp 1
transform 1 0 7452 0 -1 103360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1122
timestamp 1636968456
transform 1 0 104328 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1134
timestamp 1636968456
transform 1 0 105432 0 -1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_185_1146
timestamp 1636968456
transform 1 0 106536 0 -1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_1158
timestamp 1
transform 1 0 107640 0 -1 103360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_185_1166
timestamp 1
transform 1 0 108376 0 -1 103360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_186_3
timestamp 1636968456
transform 1 0 1380 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_15
timestamp 1636968456
transform 1 0 2484 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_186_27
timestamp 1
transform 1 0 3588 0 1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_186_29
timestamp 1636968456
transform 1 0 3772 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_41
timestamp 1636968456
transform 1 0 4876 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_53
timestamp 1636968456
transform 1 0 5980 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_186_65
timestamp 1
transform 1 0 7084 0 1 103360
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1122
timestamp 1636968456
transform 1 0 104328 0 1 103360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1134
timestamp 1636968456
transform 1 0 105432 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_186_1146
timestamp 1
transform 1 0 106536 0 1 103360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_186_1148
timestamp 1636968456
transform 1 0 106720 0 1 103360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_1160
timestamp 1
transform 1 0 107824 0 1 103360
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_187_8
timestamp 1636968456
transform 1 0 1840 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_20
timestamp 1636968456
transform 1 0 2944 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_32
timestamp 1636968456
transform 1 0 4048 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_44
timestamp 1636968456
transform 1 0 5152 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_57
timestamp 1636968456
transform 1 0 6348 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_187_69
timestamp 1
transform 1 0 7452 0 -1 104448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1122
timestamp 1636968456
transform 1 0 104328 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1134
timestamp 1636968456
transform 1 0 105432 0 -1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_187_1146
timestamp 1636968456
transform 1 0 106536 0 -1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_187_1158
timestamp 1
transform 1 0 107640 0 -1 104448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_187_1166
timestamp 1
transform 1 0 108376 0 -1 104448
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_188_3
timestamp 1636968456
transform 1 0 1380 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_15
timestamp 1636968456
transform 1 0 2484 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_188_27
timestamp 1
transform 1 0 3588 0 1 104448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_188_29
timestamp 1636968456
transform 1 0 3772 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_41
timestamp 1636968456
transform 1 0 4876 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_53
timestamp 1636968456
transform 1 0 5980 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_188_65
timestamp 1
transform 1 0 7084 0 1 104448
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1122
timestamp 1636968456
transform 1 0 104328 0 1 104448
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1134
timestamp 1636968456
transform 1 0 105432 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_188_1146
timestamp 1
transform 1 0 106536 0 1 104448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_188_1148
timestamp 1636968456
transform 1 0 106720 0 1 104448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_188_1160
timestamp 1
transform 1 0 107824 0 1 104448
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_189_3
timestamp 1636968456
transform 1 0 1380 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_15
timestamp 1636968456
transform 1 0 2484 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_27
timestamp 1636968456
transform 1 0 3588 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_39
timestamp 1636968456
transform 1 0 4692 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_189_51
timestamp 1
transform 1 0 5796 0 -1 105536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_189_55
timestamp 1
transform 1 0 6164 0 -1 105536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_189_57
timestamp 1636968456
transform 1 0 6348 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_189_69
timestamp 1
transform 1 0 7452 0 -1 105536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1122
timestamp 1636968456
transform 1 0 104328 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1134
timestamp 1636968456
transform 1 0 105432 0 -1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_189_1146
timestamp 1636968456
transform 1 0 106536 0 -1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_1158
timestamp 1
transform 1 0 107640 0 -1 105536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_189_1166
timestamp 1
transform 1 0 108376 0 -1 105536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_190_8
timestamp 1636968456
transform 1 0 1840 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_190_20
timestamp 1
transform 1 0 2944 0 1 105536
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_190_29
timestamp 1636968456
transform 1 0 3772 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_41
timestamp 1636968456
transform 1 0 4876 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_53
timestamp 1636968456
transform 1 0 5980 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_190_65
timestamp 1
transform 1 0 7084 0 1 105536
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1122
timestamp 1636968456
transform 1 0 104328 0 1 105536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1134
timestamp 1636968456
transform 1 0 105432 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_190_1146
timestamp 1
transform 1 0 106536 0 1 105536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_190_1148
timestamp 1636968456
transform 1 0 106720 0 1 105536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_190_1160
timestamp 1
transform 1 0 107824 0 1 105536
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_191_3
timestamp 1636968456
transform 1 0 1380 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_15
timestamp 1636968456
transform 1 0 2484 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_27
timestamp 1636968456
transform 1 0 3588 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_39
timestamp 1636968456
transform 1 0 4692 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_191_51
timestamp 1
transform 1 0 5796 0 -1 106624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_191_55
timestamp 1
transform 1 0 6164 0 -1 106624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_191_57
timestamp 1636968456
transform 1 0 6348 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_191_69
timestamp 1
transform 1 0 7452 0 -1 106624
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1122
timestamp 1636968456
transform 1 0 104328 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1134
timestamp 1636968456
transform 1 0 105432 0 -1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_191_1146
timestamp 1636968456
transform 1 0 106536 0 -1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_1158
timestamp 1
transform 1 0 107640 0 -1 106624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_191_1166
timestamp 1
transform 1 0 108376 0 -1 106624
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_192_8
timestamp 1636968456
transform 1 0 1840 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_20
timestamp 1
transform 1 0 2944 0 1 106624
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_192_29
timestamp 1636968456
transform 1 0 3772 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_41
timestamp 1636968456
transform 1 0 4876 0 1 106624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_192_53
timestamp 1636968456
transform 1 0 5980 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_192_65
timestamp 1
transform 1 0 7084 0 1 106624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_1146
timestamp 1
transform 1 0 106536 0 1 106624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_192_1148
timestamp 1636968456
transform 1 0 106720 0 1 106624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_1160
timestamp 1
transform 1 0 107824 0 1 106624
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_193_3
timestamp 1636968456
transform 1 0 1380 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_15
timestamp 1636968456
transform 1 0 2484 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_27
timestamp 1636968456
transform 1 0 3588 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_39
timestamp 1636968456
transform 1 0 4692 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_193_51
timestamp 1
transform 1 0 5796 0 -1 107712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_193_55
timestamp 1
transform 1 0 6164 0 -1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_193_57
timestamp 1636968456
transform 1 0 6348 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_193_69
timestamp 1
transform 1 0 7452 0 -1 107712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1122
timestamp 1636968456
transform 1 0 104328 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1134
timestamp 1636968456
transform 1 0 105432 0 -1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_193_1146
timestamp 1636968456
transform 1 0 106536 0 -1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_1158
timestamp 1
transform 1 0 107640 0 -1 107712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_193_1166
timestamp 1
transform 1 0 108376 0 -1 107712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_194_3
timestamp 1636968456
transform 1 0 1380 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_15
timestamp 1636968456
transform 1 0 2484 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_194_27
timestamp 1
transform 1 0 3588 0 1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_194_29
timestamp 1636968456
transform 1 0 3772 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_41
timestamp 1636968456
transform 1 0 4876 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_53
timestamp 1636968456
transform 1 0 5980 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_194_65
timestamp 1
transform 1 0 7084 0 1 107712
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1122
timestamp 1636968456
transform 1 0 104328 0 1 107712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1134
timestamp 1636968456
transform 1 0 105432 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_194_1146
timestamp 1
transform 1 0 106536 0 1 107712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_194_1148
timestamp 1636968456
transform 1 0 106720 0 1 107712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_194_1160
timestamp 1
transform 1 0 107824 0 1 107712
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_195_8
timestamp 1636968456
transform 1 0 1840 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_20
timestamp 1636968456
transform 1 0 2944 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_32
timestamp 1636968456
transform 1 0 4048 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_44
timestamp 1636968456
transform 1 0 5152 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_57
timestamp 1636968456
transform 1 0 6348 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_195_69
timestamp 1
transform 1 0 7452 0 -1 108800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1122
timestamp 1636968456
transform 1 0 104328 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1134
timestamp 1636968456
transform 1 0 105432 0 -1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_195_1146
timestamp 1636968456
transform 1 0 106536 0 -1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_195_1158
timestamp 1
transform 1 0 107640 0 -1 108800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_195_1166
timestamp 1
transform 1 0 108376 0 -1 108800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_196_3
timestamp 1636968456
transform 1 0 1380 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_15
timestamp 1636968456
transform 1 0 2484 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_196_27
timestamp 1
transform 1 0 3588 0 1 108800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_196_29
timestamp 1636968456
transform 1 0 3772 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_41
timestamp 1636968456
transform 1 0 4876 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_53
timestamp 1636968456
transform 1 0 5980 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_196_65
timestamp 1
transform 1 0 7084 0 1 108800
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1122
timestamp 1636968456
transform 1 0 104328 0 1 108800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1134
timestamp 1636968456
transform 1 0 105432 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_196_1146
timestamp 1
transform 1 0 106536 0 1 108800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_196_1148
timestamp 1636968456
transform 1 0 106720 0 1 108800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_196_1160
timestamp 1
transform 1 0 107824 0 1 108800
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_197_8
timestamp 1636968456
transform 1 0 1840 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_20
timestamp 1636968456
transform 1 0 2944 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_32
timestamp 1636968456
transform 1 0 4048 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_44
timestamp 1636968456
transform 1 0 5152 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_57
timestamp 1636968456
transform 1 0 6348 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_197_69
timestamp 1
transform 1 0 7452 0 -1 109888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1122
timestamp 1636968456
transform 1 0 104328 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1134
timestamp 1636968456
transform 1 0 105432 0 -1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_197_1146
timestamp 1636968456
transform 1 0 106536 0 -1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_1158
timestamp 1
transform 1 0 107640 0 -1 109888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_197_1166
timestamp 1
transform 1 0 108376 0 -1 109888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_198_3
timestamp 1636968456
transform 1 0 1380 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_15
timestamp 1636968456
transform 1 0 2484 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_198_27
timestamp 1
transform 1 0 3588 0 1 109888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_198_29
timestamp 1636968456
transform 1 0 3772 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_41
timestamp 1636968456
transform 1 0 4876 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_53
timestamp 1636968456
transform 1 0 5980 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_198_65
timestamp 1
transform 1 0 7084 0 1 109888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1122
timestamp 1636968456
transform 1 0 104328 0 1 109888
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1134
timestamp 1636968456
transform 1 0 105432 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_198_1146
timestamp 1
transform 1 0 106536 0 1 109888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_198_1148
timestamp 1636968456
transform 1 0 106720 0 1 109888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_198_1160
timestamp 1
transform 1 0 107824 0 1 109888
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_199_3
timestamp 1636968456
transform 1 0 1380 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_15
timestamp 1636968456
transform 1 0 2484 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_27
timestamp 1636968456
transform 1 0 3588 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_39
timestamp 1636968456
transform 1 0 4692 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_199_51
timestamp 1
transform 1 0 5796 0 -1 110976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_199_55
timestamp 1
transform 1 0 6164 0 -1 110976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_199_57
timestamp 1636968456
transform 1 0 6348 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_199_69
timestamp 1
transform 1 0 7452 0 -1 110976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1122
timestamp 1636968456
transform 1 0 104328 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1134
timestamp 1636968456
transform 1 0 105432 0 -1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_199_1146
timestamp 1636968456
transform 1 0 106536 0 -1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_1158
timestamp 1
transform 1 0 107640 0 -1 110976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_199_1166
timestamp 1
transform 1 0 108376 0 -1 110976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_200_8
timestamp 1636968456
transform 1 0 1840 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_200_20
timestamp 1
transform 1 0 2944 0 1 110976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_200_29
timestamp 1636968456
transform 1 0 3772 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_41
timestamp 1636968456
transform 1 0 4876 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_53
timestamp 1636968456
transform 1 0 5980 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_200_65
timestamp 1
transform 1 0 7084 0 1 110976
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1122
timestamp 1636968456
transform 1 0 104328 0 1 110976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1134
timestamp 1636968456
transform 1 0 105432 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_200_1146
timestamp 1
transform 1 0 106536 0 1 110976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_200_1148
timestamp 1636968456
transform 1 0 106720 0 1 110976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_200_1160
timestamp 1
transform 1 0 107824 0 1 110976
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_201_3
timestamp 1636968456
transform 1 0 1380 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_15
timestamp 1636968456
transform 1 0 2484 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_27
timestamp 1636968456
transform 1 0 3588 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_39
timestamp 1636968456
transform 1 0 4692 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_201_51
timestamp 1
transform 1 0 5796 0 -1 112064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_201_55
timestamp 1
transform 1 0 6164 0 -1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_201_57
timestamp 1636968456
transform 1 0 6348 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_201_69
timestamp 1
transform 1 0 7452 0 -1 112064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1122
timestamp 1636968456
transform 1 0 104328 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1134
timestamp 1636968456
transform 1 0 105432 0 -1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_201_1146
timestamp 1636968456
transform 1 0 106536 0 -1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_1158
timestamp 1
transform 1 0 107640 0 -1 112064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_201_1166
timestamp 1
transform 1 0 108376 0 -1 112064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_202_3
timestamp 1636968456
transform 1 0 1380 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_15
timestamp 1636968456
transform 1 0 2484 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_202_27
timestamp 1
transform 1 0 3588 0 1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_202_29
timestamp 1636968456
transform 1 0 3772 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_41
timestamp 1636968456
transform 1 0 4876 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_53
timestamp 1636968456
transform 1 0 5980 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_202_65
timestamp 1
transform 1 0 7084 0 1 112064
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1122
timestamp 1636968456
transform 1 0 104328 0 1 112064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1134
timestamp 1636968456
transform 1 0 105432 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_202_1146
timestamp 1
transform 1 0 106536 0 1 112064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_202_1148
timestamp 1636968456
transform 1 0 106720 0 1 112064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_202_1160
timestamp 1
transform 1 0 107824 0 1 112064
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_203_3
timestamp 1636968456
transform 1 0 1380 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_15
timestamp 1636968456
transform 1 0 2484 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_27
timestamp 1636968456
transform 1 0 3588 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_39
timestamp 1636968456
transform 1 0 4692 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_203_51
timestamp 1
transform 1 0 5796 0 -1 113152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_203_55
timestamp 1
transform 1 0 6164 0 -1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_203_57
timestamp 1636968456
transform 1 0 6348 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_203_69
timestamp 1
transform 1 0 7452 0 -1 113152
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1124
timestamp 1636968456
transform 1 0 104512 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1136
timestamp 1636968456
transform 1 0 105616 0 -1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_203_1148
timestamp 1636968456
transform 1 0 106720 0 -1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_203_1160
timestamp 1
transform 1 0 107824 0 -1 113152
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_204_3
timestamp 1636968456
transform 1 0 1380 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_15
timestamp 1636968456
transform 1 0 2484 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_204_27
timestamp 1
transform 1 0 3588 0 1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_204_29
timestamp 1636968456
transform 1 0 3772 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_41
timestamp 1636968456
transform 1 0 4876 0 1 113152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_204_53
timestamp 1636968456
transform 1 0 5980 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_204_65
timestamp 1
transform 1 0 7084 0 1 113152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_204_1142
timestamp 1
transform 1 0 106168 0 1 113152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_204_1146
timestamp 1
transform 1 0 106536 0 1 113152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_204_1148
timestamp 1636968456
transform 1 0 106720 0 1 113152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_204_1160
timestamp 1
transform 1 0 107824 0 1 113152
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_205_3
timestamp 1636968456
transform 1 0 1380 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_15
timestamp 1636968456
transform 1 0 2484 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_27
timestamp 1636968456
transform 1 0 3588 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_39
timestamp 1636968456
transform 1 0 4692 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_205_51
timestamp 1
transform 1 0 5796 0 -1 114240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_205_55
timestamp 1
transform 1 0 6164 0 -1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_205_57
timestamp 1636968456
transform 1 0 6348 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_205_69
timestamp 1
transform 1 0 7452 0 -1 114240
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1122
timestamp 1636968456
transform 1 0 104328 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1134
timestamp 1636968456
transform 1 0 105432 0 -1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_205_1146
timestamp 1636968456
transform 1 0 106536 0 -1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_205_1158
timestamp 1
transform 1 0 107640 0 -1 114240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_205_1166
timestamp 1
transform 1 0 108376 0 -1 114240
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_206_3
timestamp 1636968456
transform 1 0 1380 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_15
timestamp 1636968456
transform 1 0 2484 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_206_27
timestamp 1
transform 1 0 3588 0 1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_206_29
timestamp 1636968456
transform 1 0 3772 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_41
timestamp 1636968456
transform 1 0 4876 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_53
timestamp 1636968456
transform 1 0 5980 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_206_65
timestamp 1
transform 1 0 7084 0 1 114240
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1122
timestamp 1636968456
transform 1 0 104328 0 1 114240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1134
timestamp 1636968456
transform 1 0 105432 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_206_1146
timestamp 1
transform 1 0 106536 0 1 114240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_206_1148
timestamp 1636968456
transform 1 0 106720 0 1 114240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_206_1160
timestamp 1
transform 1 0 107824 0 1 114240
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_207_3
timestamp 1636968456
transform 1 0 1380 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_15
timestamp 1636968456
transform 1 0 2484 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_27
timestamp 1636968456
transform 1 0 3588 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_39
timestamp 1636968456
transform 1 0 4692 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_207_51
timestamp 1
transform 1 0 5796 0 -1 115328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_55
timestamp 1
transform 1 0 6164 0 -1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_207_57
timestamp 1636968456
transform 1 0 6348 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_207_69
timestamp 1
transform 1 0 7452 0 -1 115328
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1122
timestamp 1636968456
transform 1 0 104328 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1134
timestamp 1636968456
transform 1 0 105432 0 -1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_207_1146
timestamp 1636968456
transform 1 0 106536 0 -1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_207_1158
timestamp 1
transform 1 0 107640 0 -1 115328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_207_1166
timestamp 1
transform 1 0 108376 0 -1 115328
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_208_3
timestamp 1636968456
transform 1 0 1380 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_15
timestamp 1636968456
transform 1 0 2484 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_208_27
timestamp 1
transform 1 0 3588 0 1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_208_29
timestamp 1636968456
transform 1 0 3772 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_41
timestamp 1636968456
transform 1 0 4876 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_53
timestamp 1636968456
transform 1 0 5980 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_208_65
timestamp 1
transform 1 0 7084 0 1 115328
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1122
timestamp 1636968456
transform 1 0 104328 0 1 115328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1134
timestamp 1636968456
transform 1 0 105432 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_208_1146
timestamp 1
transform 1 0 106536 0 1 115328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_208_1148
timestamp 1636968456
transform 1 0 106720 0 1 115328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_208_1160
timestamp 1
transform 1 0 107824 0 1 115328
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_209_3
timestamp 1636968456
transform 1 0 1380 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_15
timestamp 1636968456
transform 1 0 2484 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_27
timestamp 1636968456
transform 1 0 3588 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_39
timestamp 1636968456
transform 1 0 4692 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_209_51
timestamp 1
transform 1 0 5796 0 -1 116416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_55
timestamp 1
transform 1 0 6164 0 -1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_209_57
timestamp 1636968456
transform 1 0 6348 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_209_69
timestamp 1
transform 1 0 7452 0 -1 116416
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1122
timestamp 1636968456
transform 1 0 104328 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1134
timestamp 1636968456
transform 1 0 105432 0 -1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_209_1146
timestamp 1636968456
transform 1 0 106536 0 -1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_209_1158
timestamp 1
transform 1 0 107640 0 -1 116416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_209_1166
timestamp 1
transform 1 0 108376 0 -1 116416
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_210_3
timestamp 1636968456
transform 1 0 1380 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_15
timestamp 1636968456
transform 1 0 2484 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_210_27
timestamp 1
transform 1 0 3588 0 1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_210_29
timestamp 1636968456
transform 1 0 3772 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_41
timestamp 1636968456
transform 1 0 4876 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_53
timestamp 1636968456
transform 1 0 5980 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_210_65
timestamp 1
transform 1 0 7084 0 1 116416
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1122
timestamp 1636968456
transform 1 0 104328 0 1 116416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1134
timestamp 1636968456
transform 1 0 105432 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_210_1146
timestamp 1
transform 1 0 106536 0 1 116416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_210_1148
timestamp 1636968456
transform 1 0 106720 0 1 116416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_210_1160
timestamp 1
transform 1 0 107824 0 1 116416
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_211_3
timestamp 1636968456
transform 1 0 1380 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_15
timestamp 1636968456
transform 1 0 2484 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_27
timestamp 1636968456
transform 1 0 3588 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_39
timestamp 1636968456
transform 1 0 4692 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_211_51
timestamp 1
transform 1 0 5796 0 -1 117504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_211_55
timestamp 1
transform 1 0 6164 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_211_57
timestamp 1
transform 1 0 6348 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_211_65
timestamp 1
transform 1 0 7084 0 -1 117504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1122
timestamp 1636968456
transform 1 0 104328 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1134
timestamp 1636968456
transform 1 0 105432 0 -1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_211_1146
timestamp 1636968456
transform 1 0 106536 0 -1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_211_1158
timestamp 1
transform 1 0 107640 0 -1 117504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_211_1166
timestamp 1
transform 1 0 108376 0 -1 117504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_212_3
timestamp 1636968456
transform 1 0 1380 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_15
timestamp 1636968456
transform 1 0 2484 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_212_27
timestamp 1
transform 1 0 3588 0 1 117504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_212_29
timestamp 1636968456
transform 1 0 3772 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_41
timestamp 1636968456
transform 1 0 4876 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_212_53
timestamp 1
transform 1 0 5980 0 1 117504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1122
timestamp 1636968456
transform 1 0 104328 0 1 117504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1134
timestamp 1636968456
transform 1 0 105432 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_212_1146
timestamp 1
transform 1 0 106536 0 1 117504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_212_1148
timestamp 1636968456
transform 1 0 106720 0 1 117504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_212_1160
timestamp 1
transform 1 0 107824 0 1 117504
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_213_3
timestamp 1636968456
transform 1 0 1380 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_15
timestamp 1636968456
transform 1 0 2484 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_27
timestamp 1636968456
transform 1 0 3588 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_39
timestamp 1636968456
transform 1 0 4692 0 -1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_213_51
timestamp 1
transform 1 0 5796 0 -1 118592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_213_55
timestamp 1
transform 1 0 6164 0 -1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_213_57
timestamp 1636968456
transform 1 0 6348 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1122
timestamp 1636968456
transform 1 0 104328 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1134
timestamp 1636968456
transform 1 0 105432 0 -1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_213_1146
timestamp 1636968456
transform 1 0 106536 0 -1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_213_1158
timestamp 1
transform 1 0 107640 0 -1 118592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_213_1166
timestamp 1
transform 1 0 108376 0 -1 118592
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_214_3
timestamp 1636968456
transform 1 0 1380 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_15
timestamp 1636968456
transform 1 0 2484 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_214_27
timestamp 1
transform 1 0 3588 0 1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_214_29
timestamp 1636968456
transform 1 0 3772 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_41
timestamp 1636968456
transform 1 0 4876 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_53
timestamp 1636968456
transform 1 0 5980 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_214_65
timestamp 1
transform 1 0 7084 0 1 118592
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1122
timestamp 1636968456
transform 1 0 104328 0 1 118592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1134
timestamp 1636968456
transform 1 0 105432 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_214_1146
timestamp 1
transform 1 0 106536 0 1 118592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_214_1148
timestamp 1636968456
transform 1 0 106720 0 1 118592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_214_1160
timestamp 1
transform 1 0 107824 0 1 118592
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_215_3
timestamp 1636968456
transform 1 0 1380 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_15
timestamp 1636968456
transform 1 0 2484 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_27
timestamp 1636968456
transform 1 0 3588 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_39
timestamp 1636968456
transform 1 0 4692 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_215_51
timestamp 1
transform 1 0 5796 0 -1 119680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_215_55
timestamp 1
transform 1 0 6164 0 -1 119680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_215_57
timestamp 1636968456
transform 1 0 6348 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_215_69
timestamp 1
transform 1 0 7452 0 -1 119680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1122
timestamp 1636968456
transform 1 0 104328 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1134
timestamp 1636968456
transform 1 0 105432 0 -1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_215_1146
timestamp 1636968456
transform 1 0 106536 0 -1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_215_1158
timestamp 1
transform 1 0 107640 0 -1 119680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_215_1166
timestamp 1
transform 1 0 108376 0 -1 119680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_216_3
timestamp 1636968456
transform 1 0 1380 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_15
timestamp 1636968456
transform 1 0 2484 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_216_27
timestamp 1
transform 1 0 3588 0 1 119680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_216_29
timestamp 1636968456
transform 1 0 3772 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_41
timestamp 1636968456
transform 1 0 4876 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_53
timestamp 1636968456
transform 1 0 5980 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_216_65
timestamp 1
transform 1 0 7084 0 1 119680
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_216_1122
timestamp 1636968456
transform 1 0 104328 0 1 119680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_216_1134
timestamp 1636968456
transform 1 0 105432 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_216_1146
timestamp 1
transform 1 0 106536 0 1 119680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_216_1148
timestamp 1636968456
transform 1 0 106720 0 1 119680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_216_1160
timestamp 1
transform 1 0 107824 0 1 119680
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_217_3
timestamp 1636968456
transform 1 0 1380 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_15
timestamp 1636968456
transform 1 0 2484 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_27
timestamp 1636968456
transform 1 0 3588 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_39
timestamp 1636968456
transform 1 0 4692 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_217_51
timestamp 1
transform 1 0 5796 0 -1 120768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_217_55
timestamp 1
transform 1 0 6164 0 -1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_217_57
timestamp 1636968456
transform 1 0 6348 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_217_69
timestamp 1
transform 1 0 7452 0 -1 120768
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1122
timestamp 1636968456
transform 1 0 104328 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1134
timestamp 1636968456
transform 1 0 105432 0 -1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_217_1146
timestamp 1636968456
transform 1 0 106536 0 -1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_217_1158
timestamp 1
transform 1 0 107640 0 -1 120768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_217_1166
timestamp 1
transform 1 0 108376 0 -1 120768
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_218_3
timestamp 1636968456
transform 1 0 1380 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_15
timestamp 1636968456
transform 1 0 2484 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_218_27
timestamp 1
transform 1 0 3588 0 1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_218_29
timestamp 1636968456
transform 1 0 3772 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_41
timestamp 1636968456
transform 1 0 4876 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_53
timestamp 1636968456
transform 1 0 5980 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_218_65
timestamp 1
transform 1 0 7084 0 1 120768
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1122
timestamp 1636968456
transform 1 0 104328 0 1 120768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1134
timestamp 1636968456
transform 1 0 105432 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_218_1146
timestamp 1
transform 1 0 106536 0 1 120768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_218_1148
timestamp 1636968456
transform 1 0 106720 0 1 120768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_218_1160
timestamp 1
transform 1 0 107824 0 1 120768
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_219_3
timestamp 1636968456
transform 1 0 1380 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_15
timestamp 1636968456
transform 1 0 2484 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_27
timestamp 1636968456
transform 1 0 3588 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_39
timestamp 1636968456
transform 1 0 4692 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_219_51
timestamp 1
transform 1 0 5796 0 -1 121856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_219_55
timestamp 1
transform 1 0 6164 0 -1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_219_57
timestamp 1636968456
transform 1 0 6348 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_219_69
timestamp 1
transform 1 0 7452 0 -1 121856
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1122
timestamp 1636968456
transform 1 0 104328 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1134
timestamp 1636968456
transform 1 0 105432 0 -1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_219_1146
timestamp 1636968456
transform 1 0 106536 0 -1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_219_1158
timestamp 1
transform 1 0 107640 0 -1 121856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_219_1166
timestamp 1
transform 1 0 108376 0 -1 121856
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_220_3
timestamp 1636968456
transform 1 0 1380 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_15
timestamp 1636968456
transform 1 0 2484 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_220_27
timestamp 1
transform 1 0 3588 0 1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_220_29
timestamp 1636968456
transform 1 0 3772 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_41
timestamp 1636968456
transform 1 0 4876 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_53
timestamp 1636968456
transform 1 0 5980 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_220_65
timestamp 1
transform 1 0 7084 0 1 121856
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1122
timestamp 1636968456
transform 1 0 104328 0 1 121856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1134
timestamp 1636968456
transform 1 0 105432 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_220_1146
timestamp 1
transform 1 0 106536 0 1 121856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_220_1148
timestamp 1636968456
transform 1 0 106720 0 1 121856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_220_1160
timestamp 1
transform 1 0 107824 0 1 121856
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_221_3
timestamp 1636968456
transform 1 0 1380 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_15
timestamp 1636968456
transform 1 0 2484 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_27
timestamp 1636968456
transform 1 0 3588 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_39
timestamp 1636968456
transform 1 0 4692 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_221_51
timestamp 1
transform 1 0 5796 0 -1 122944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_221_55
timestamp 1
transform 1 0 6164 0 -1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_221_57
timestamp 1636968456
transform 1 0 6348 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_221_69
timestamp 1
transform 1 0 7452 0 -1 122944
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1122
timestamp 1636968456
transform 1 0 104328 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1134
timestamp 1636968456
transform 1 0 105432 0 -1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_221_1146
timestamp 1636968456
transform 1 0 106536 0 -1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_221_1158
timestamp 1
transform 1 0 107640 0 -1 122944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_221_1166
timestamp 1
transform 1 0 108376 0 -1 122944
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_222_3
timestamp 1636968456
transform 1 0 1380 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_15
timestamp 1636968456
transform 1 0 2484 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_222_27
timestamp 1
transform 1 0 3588 0 1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_222_29
timestamp 1636968456
transform 1 0 3772 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_41
timestamp 1636968456
transform 1 0 4876 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_53
timestamp 1636968456
transform 1 0 5980 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_222_65
timestamp 1
transform 1 0 7084 0 1 122944
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1122
timestamp 1636968456
transform 1 0 104328 0 1 122944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1134
timestamp 1636968456
transform 1 0 105432 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_222_1146
timestamp 1
transform 1 0 106536 0 1 122944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_222_1148
timestamp 1636968456
transform 1 0 106720 0 1 122944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_222_1160
timestamp 1
transform 1 0 107824 0 1 122944
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_223_3
timestamp 1636968456
transform 1 0 1380 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_15
timestamp 1636968456
transform 1 0 2484 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_27
timestamp 1636968456
transform 1 0 3588 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_39
timestamp 1636968456
transform 1 0 4692 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_223_51
timestamp 1
transform 1 0 5796 0 -1 124032
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_223_55
timestamp 1
transform 1 0 6164 0 -1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_223_57
timestamp 1636968456
transform 1 0 6348 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_223_69
timestamp 1
transform 1 0 7452 0 -1 124032
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1122
timestamp 1636968456
transform 1 0 104328 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1134
timestamp 1636968456
transform 1 0 105432 0 -1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_223_1146
timestamp 1636968456
transform 1 0 106536 0 -1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_223_1158
timestamp 1
transform 1 0 107640 0 -1 124032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_223_1166
timestamp 1
transform 1 0 108376 0 -1 124032
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_224_3
timestamp 1636968456
transform 1 0 1380 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_15
timestamp 1636968456
transform 1 0 2484 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_224_27
timestamp 1
transform 1 0 3588 0 1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_224_29
timestamp 1636968456
transform 1 0 3772 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_41
timestamp 1636968456
transform 1 0 4876 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_53
timestamp 1636968456
transform 1 0 5980 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_224_65
timestamp 1
transform 1 0 7084 0 1 124032
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1122
timestamp 1636968456
transform 1 0 104328 0 1 124032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1134
timestamp 1636968456
transform 1 0 105432 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_224_1146
timestamp 1
transform 1 0 106536 0 1 124032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_224_1148
timestamp 1636968456
transform 1 0 106720 0 1 124032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_224_1160
timestamp 1
transform 1 0 107824 0 1 124032
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_225_3
timestamp 1636968456
transform 1 0 1380 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_15
timestamp 1636968456
transform 1 0 2484 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_27
timestamp 1636968456
transform 1 0 3588 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_39
timestamp 1636968456
transform 1 0 4692 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_225_51
timestamp 1
transform 1 0 5796 0 -1 125120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_225_55
timestamp 1
transform 1 0 6164 0 -1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_225_57
timestamp 1636968456
transform 1 0 6348 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_225_69
timestamp 1
transform 1 0 7452 0 -1 125120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1122
timestamp 1636968456
transform 1 0 104328 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1134
timestamp 1636968456
transform 1 0 105432 0 -1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_225_1146
timestamp 1636968456
transform 1 0 106536 0 -1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_225_1158
timestamp 1
transform 1 0 107640 0 -1 125120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_225_1166
timestamp 1
transform 1 0 108376 0 -1 125120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_226_3
timestamp 1636968456
transform 1 0 1380 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_15
timestamp 1636968456
transform 1 0 2484 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_226_27
timestamp 1
transform 1 0 3588 0 1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_226_29
timestamp 1636968456
transform 1 0 3772 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_41
timestamp 1636968456
transform 1 0 4876 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_53
timestamp 1636968456
transform 1 0 5980 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_226_65
timestamp 1
transform 1 0 7084 0 1 125120
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1122
timestamp 1636968456
transform 1 0 104328 0 1 125120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1134
timestamp 1636968456
transform 1 0 105432 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_226_1146
timestamp 1
transform 1 0 106536 0 1 125120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_226_1148
timestamp 1636968456
transform 1 0 106720 0 1 125120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_226_1160
timestamp 1
transform 1 0 107824 0 1 125120
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_227_3
timestamp 1636968456
transform 1 0 1380 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_15
timestamp 1636968456
transform 1 0 2484 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_27
timestamp 1636968456
transform 1 0 3588 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_39
timestamp 1636968456
transform 1 0 4692 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_227_51
timestamp 1
transform 1 0 5796 0 -1 126208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_227_55
timestamp 1
transform 1 0 6164 0 -1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_227_57
timestamp 1636968456
transform 1 0 6348 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_227_69
timestamp 1
transform 1 0 7452 0 -1 126208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1122
timestamp 1636968456
transform 1 0 104328 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1134
timestamp 1636968456
transform 1 0 105432 0 -1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_227_1146
timestamp 1636968456
transform 1 0 106536 0 -1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_227_1158
timestamp 1
transform 1 0 107640 0 -1 126208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_227_1166
timestamp 1
transform 1 0 108376 0 -1 126208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_228_3
timestamp 1636968456
transform 1 0 1380 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_15
timestamp 1636968456
transform 1 0 2484 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_228_27
timestamp 1
transform 1 0 3588 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_29
timestamp 1636968456
transform 1 0 3772 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_41
timestamp 1636968456
transform 1 0 4876 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_53
timestamp 1636968456
transform 1 0 5980 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_228_65
timestamp 1
transform 1 0 7084 0 1 126208
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1122
timestamp 1636968456
transform 1 0 104328 0 1 126208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1134
timestamp 1636968456
transform 1 0 105432 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_228_1146
timestamp 1
transform 1 0 106536 0 1 126208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_228_1148
timestamp 1636968456
transform 1 0 106720 0 1 126208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_228_1160
timestamp 1
transform 1 0 107824 0 1 126208
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_229_3
timestamp 1636968456
transform 1 0 1380 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_15
timestamp 1636968456
transform 1 0 2484 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_27
timestamp 1636968456
transform 1 0 3588 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_39
timestamp 1636968456
transform 1 0 4692 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_229_51
timestamp 1
transform 1 0 5796 0 -1 127296
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_229_55
timestamp 1
transform 1 0 6164 0 -1 127296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_229_57
timestamp 1636968456
transform 1 0 6348 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_229_69
timestamp 1
transform 1 0 7452 0 -1 127296
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1122
timestamp 1636968456
transform 1 0 104328 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1134
timestamp 1636968456
transform 1 0 105432 0 -1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_229_1146
timestamp 1636968456
transform 1 0 106536 0 -1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_229_1158
timestamp 1
transform 1 0 107640 0 -1 127296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_229_1166
timestamp 1
transform 1 0 108376 0 -1 127296
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_230_3
timestamp 1636968456
transform 1 0 1380 0 1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_230_15
timestamp 1636968456
transform 1 0 2484 0 1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_230_27
timestamp 1
transform 1 0 3588 0 1 127296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_230_29
timestamp 1636968456
transform 1 0 3772 0 1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_230_41
timestamp 1636968456
transform 1 0 4876 0 1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_230_53
timestamp 1636968456
transform 1 0 5980 0 1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_230_65
timestamp 1
transform 1 0 7084 0 1 127296
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_230_1122
timestamp 1636968456
transform 1 0 104328 0 1 127296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_230_1134
timestamp 1636968456
transform 1 0 105432 0 1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_230_1146
timestamp 1
transform 1 0 106536 0 1 127296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_230_1148
timestamp 1636968456
transform 1 0 106720 0 1 127296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_230_1160
timestamp 1
transform 1 0 107824 0 1 127296
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_231_3
timestamp 1636968456
transform 1 0 1380 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_15
timestamp 1636968456
transform 1 0 2484 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_27
timestamp 1636968456
transform 1 0 3588 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_39
timestamp 1636968456
transform 1 0 4692 0 -1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_231_51
timestamp 1
transform 1 0 5796 0 -1 128384
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_231_55
timestamp 1
transform 1 0 6164 0 -1 128384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_231_57
timestamp 1636968456
transform 1 0 6348 0 -1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_231_69
timestamp 1
transform 1 0 7452 0 -1 128384
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_231_1122
timestamp 1636968456
transform 1 0 104328 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_1134
timestamp 1636968456
transform 1 0 105432 0 -1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_231_1146
timestamp 1636968456
transform 1 0 106536 0 -1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_231_1158
timestamp 1
transform 1 0 107640 0 -1 128384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_231_1166
timestamp 1
transform 1 0 108376 0 -1 128384
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_232_3
timestamp 1636968456
transform 1 0 1380 0 1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_232_15
timestamp 1636968456
transform 1 0 2484 0 1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_232_27
timestamp 1
transform 1 0 3588 0 1 128384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_232_29
timestamp 1636968456
transform 1 0 3772 0 1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_232_41
timestamp 1636968456
transform 1 0 4876 0 1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_232_53
timestamp 1636968456
transform 1 0 5980 0 1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_232_65
timestamp 1
transform 1 0 7084 0 1 128384
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_232_1122
timestamp 1636968456
transform 1 0 104328 0 1 128384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_232_1134
timestamp 1636968456
transform 1 0 105432 0 1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_232_1146
timestamp 1
transform 1 0 106536 0 1 128384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_232_1148
timestamp 1636968456
transform 1 0 106720 0 1 128384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_232_1160
timestamp 1
transform 1 0 107824 0 1 128384
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_233_3
timestamp 1636968456
transform 1 0 1380 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_15
timestamp 1636968456
transform 1 0 2484 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_27
timestamp 1636968456
transform 1 0 3588 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_39
timestamp 1636968456
transform 1 0 4692 0 -1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_233_51
timestamp 1
transform 1 0 5796 0 -1 129472
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_233_55
timestamp 1
transform 1 0 6164 0 -1 129472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_233_57
timestamp 1636968456
transform 1 0 6348 0 -1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_233_69
timestamp 1
transform 1 0 7452 0 -1 129472
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_233_1122
timestamp 1636968456
transform 1 0 104328 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_1134
timestamp 1636968456
transform 1 0 105432 0 -1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_233_1146
timestamp 1636968456
transform 1 0 106536 0 -1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_233_1158
timestamp 1
transform 1 0 107640 0 -1 129472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_233_1166
timestamp 1
transform 1 0 108376 0 -1 129472
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_234_3
timestamp 1636968456
transform 1 0 1380 0 1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_234_15
timestamp 1636968456
transform 1 0 2484 0 1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_234_27
timestamp 1
transform 1 0 3588 0 1 129472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_234_29
timestamp 1636968456
transform 1 0 3772 0 1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_234_41
timestamp 1636968456
transform 1 0 4876 0 1 129472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_234_53
timestamp 1636968456
transform 1 0 5980 0 1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_234_65
timestamp 1
transform 1 0 7084 0 1 129472
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_234_1125
timestamp 1636968456
transform 1 0 104604 0 1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_234_1137
timestamp 1
transform 1 0 105708 0 1 129472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_234_1145
timestamp 1
transform 1 0 106444 0 1 129472
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_234_1148
timestamp 1636968456
transform 1 0 106720 0 1 129472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_234_1160
timestamp 1
transform 1 0 107824 0 1 129472
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_235_3
timestamp 1636968456
transform 1 0 1380 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_15
timestamp 1636968456
transform 1 0 2484 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_27
timestamp 1636968456
transform 1 0 3588 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_39
timestamp 1636968456
transform 1 0 4692 0 -1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_235_51
timestamp 1
transform 1 0 5796 0 -1 130560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_235_55
timestamp 1
transform 1 0 6164 0 -1 130560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_235_57
timestamp 1636968456
transform 1 0 6348 0 -1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_235_69
timestamp 1
transform 1 0 7452 0 -1 130560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_235_1122
timestamp 1636968456
transform 1 0 104328 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_1134
timestamp 1636968456
transform 1 0 105432 0 -1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_235_1146
timestamp 1636968456
transform 1 0 106536 0 -1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_235_1158
timestamp 1
transform 1 0 107640 0 -1 130560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_235_1166
timestamp 1
transform 1 0 108376 0 -1 130560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_236_3
timestamp 1636968456
transform 1 0 1380 0 1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_236_15
timestamp 1636968456
transform 1 0 2484 0 1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_236_27
timestamp 1
transform 1 0 3588 0 1 130560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_236_29
timestamp 1636968456
transform 1 0 3772 0 1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_236_41
timestamp 1636968456
transform 1 0 4876 0 1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_236_53
timestamp 1636968456
transform 1 0 5980 0 1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_236_65
timestamp 1
transform 1 0 7084 0 1 130560
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_236_1122
timestamp 1636968456
transform 1 0 104328 0 1 130560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_236_1134
timestamp 1636968456
transform 1 0 105432 0 1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_236_1146
timestamp 1
transform 1 0 106536 0 1 130560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_236_1148
timestamp 1636968456
transform 1 0 106720 0 1 130560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_236_1160
timestamp 1
transform 1 0 107824 0 1 130560
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_237_3
timestamp 1636968456
transform 1 0 1380 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_15
timestamp 1636968456
transform 1 0 2484 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_27
timestamp 1636968456
transform 1 0 3588 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_39
timestamp 1636968456
transform 1 0 4692 0 -1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_237_51
timestamp 1
transform 1 0 5796 0 -1 131648
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_237_55
timestamp 1
transform 1 0 6164 0 -1 131648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_237_57
timestamp 1636968456
transform 1 0 6348 0 -1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_237_69
timestamp 1
transform 1 0 7452 0 -1 131648
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_237_1122
timestamp 1636968456
transform 1 0 104328 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_1134
timestamp 1636968456
transform 1 0 105432 0 -1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_237_1146
timestamp 1636968456
transform 1 0 106536 0 -1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_237_1158
timestamp 1
transform 1 0 107640 0 -1 131648
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_237_1166
timestamp 1
transform 1 0 108376 0 -1 131648
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_238_3
timestamp 1636968456
transform 1 0 1380 0 1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_238_15
timestamp 1636968456
transform 1 0 2484 0 1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_238_27
timestamp 1
transform 1 0 3588 0 1 131648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_238_29
timestamp 1636968456
transform 1 0 3772 0 1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_238_41
timestamp 1636968456
transform 1 0 4876 0 1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_238_53
timestamp 1636968456
transform 1 0 5980 0 1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_238_65
timestamp 1
transform 1 0 7084 0 1 131648
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_238_1122
timestamp 1636968456
transform 1 0 104328 0 1 131648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_238_1134
timestamp 1636968456
transform 1 0 105432 0 1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_238_1146
timestamp 1
transform 1 0 106536 0 1 131648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_238_1148
timestamp 1636968456
transform 1 0 106720 0 1 131648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_238_1160
timestamp 1
transform 1 0 107824 0 1 131648
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_239_3
timestamp 1636968456
transform 1 0 1380 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_15
timestamp 1636968456
transform 1 0 2484 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_27
timestamp 1636968456
transform 1 0 3588 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_39
timestamp 1636968456
transform 1 0 4692 0 -1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_239_51
timestamp 1
transform 1 0 5796 0 -1 132736
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_239_55
timestamp 1
transform 1 0 6164 0 -1 132736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_239_57
timestamp 1636968456
transform 1 0 6348 0 -1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_239_69
timestamp 1
transform 1 0 7452 0 -1 132736
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_239_1122
timestamp 1636968456
transform 1 0 104328 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_1134
timestamp 1636968456
transform 1 0 105432 0 -1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_239_1146
timestamp 1636968456
transform 1 0 106536 0 -1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_239_1158
timestamp 1
transform 1 0 107640 0 -1 132736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_239_1166
timestamp 1
transform 1 0 108376 0 -1 132736
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_240_3
timestamp 1636968456
transform 1 0 1380 0 1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_240_15
timestamp 1636968456
transform 1 0 2484 0 1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_240_27
timestamp 1
transform 1 0 3588 0 1 132736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_240_29
timestamp 1636968456
transform 1 0 3772 0 1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_240_41
timestamp 1636968456
transform 1 0 4876 0 1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_240_53
timestamp 1636968456
transform 1 0 5980 0 1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_240_65
timestamp 1
transform 1 0 7084 0 1 132736
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_240_1122
timestamp 1636968456
transform 1 0 104328 0 1 132736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_240_1134
timestamp 1636968456
transform 1 0 105432 0 1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_240_1146
timestamp 1
transform 1 0 106536 0 1 132736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_240_1148
timestamp 1636968456
transform 1 0 106720 0 1 132736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_240_1160
timestamp 1
transform 1 0 107824 0 1 132736
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_241_3
timestamp 1636968456
transform 1 0 1380 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_15
timestamp 1636968456
transform 1 0 2484 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_27
timestamp 1636968456
transform 1 0 3588 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_39
timestamp 1636968456
transform 1 0 4692 0 -1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_241_51
timestamp 1
transform 1 0 5796 0 -1 133824
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_241_55
timestamp 1
transform 1 0 6164 0 -1 133824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_241_57
timestamp 1636968456
transform 1 0 6348 0 -1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_241_69
timestamp 1
transform 1 0 7452 0 -1 133824
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_241_1122
timestamp 1636968456
transform 1 0 104328 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_1134
timestamp 1636968456
transform 1 0 105432 0 -1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_241_1146
timestamp 1636968456
transform 1 0 106536 0 -1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_241_1158
timestamp 1
transform 1 0 107640 0 -1 133824
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_241_1166
timestamp 1
transform 1 0 108376 0 -1 133824
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_242_3
timestamp 1636968456
transform 1 0 1380 0 1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_242_15
timestamp 1636968456
transform 1 0 2484 0 1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_242_27
timestamp 1
transform 1 0 3588 0 1 133824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_242_29
timestamp 1636968456
transform 1 0 3772 0 1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_242_41
timestamp 1636968456
transform 1 0 4876 0 1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_242_53
timestamp 1636968456
transform 1 0 5980 0 1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_242_65
timestamp 1
transform 1 0 7084 0 1 133824
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_242_1122
timestamp 1636968456
transform 1 0 104328 0 1 133824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_242_1134
timestamp 1636968456
transform 1 0 105432 0 1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_242_1146
timestamp 1
transform 1 0 106536 0 1 133824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_242_1148
timestamp 1636968456
transform 1 0 106720 0 1 133824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_242_1160
timestamp 1
transform 1 0 107824 0 1 133824
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_243_3
timestamp 1636968456
transform 1 0 1380 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_15
timestamp 1636968456
transform 1 0 2484 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_27
timestamp 1636968456
transform 1 0 3588 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_39
timestamp 1636968456
transform 1 0 4692 0 -1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_243_51
timestamp 1
transform 1 0 5796 0 -1 134912
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_243_55
timestamp 1
transform 1 0 6164 0 -1 134912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_243_57
timestamp 1636968456
transform 1 0 6348 0 -1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_243_69
timestamp 1
transform 1 0 7452 0 -1 134912
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_243_1122
timestamp 1636968456
transform 1 0 104328 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_1134
timestamp 1636968456
transform 1 0 105432 0 -1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_243_1146
timestamp 1636968456
transform 1 0 106536 0 -1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_243_1158
timestamp 1
transform 1 0 107640 0 -1 134912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_243_1166
timestamp 1
transform 1 0 108376 0 -1 134912
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_244_3
timestamp 1636968456
transform 1 0 1380 0 1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_244_15
timestamp 1636968456
transform 1 0 2484 0 1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_244_27
timestamp 1
transform 1 0 3588 0 1 134912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_244_29
timestamp 1636968456
transform 1 0 3772 0 1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_244_41
timestamp 1636968456
transform 1 0 4876 0 1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_244_53
timestamp 1636968456
transform 1 0 5980 0 1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_244_65
timestamp 1
transform 1 0 7084 0 1 134912
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_244_1122
timestamp 1636968456
transform 1 0 104328 0 1 134912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_244_1134
timestamp 1636968456
transform 1 0 105432 0 1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_244_1146
timestamp 1
transform 1 0 106536 0 1 134912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_244_1148
timestamp 1636968456
transform 1 0 106720 0 1 134912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_244_1160
timestamp 1
transform 1 0 107824 0 1 134912
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_245_3
timestamp 1636968456
transform 1 0 1380 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_15
timestamp 1636968456
transform 1 0 2484 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_27
timestamp 1636968456
transform 1 0 3588 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_39
timestamp 1636968456
transform 1 0 4692 0 -1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_245_51
timestamp 1
transform 1 0 5796 0 -1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_245_55
timestamp 1
transform 1 0 6164 0 -1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_245_57
timestamp 1636968456
transform 1 0 6348 0 -1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_245_69
timestamp 1
transform 1 0 7452 0 -1 136000
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_245_1122
timestamp 1636968456
transform 1 0 104328 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_1134
timestamp 1636968456
transform 1 0 105432 0 -1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_245_1146
timestamp 1636968456
transform 1 0 106536 0 -1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_245_1158
timestamp 1
transform 1 0 107640 0 -1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_245_1166
timestamp 1
transform 1 0 108376 0 -1 136000
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_246_3
timestamp 1636968456
transform 1 0 1380 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_15
timestamp 1636968456
transform 1 0 2484 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_246_27
timestamp 1
transform 1 0 3588 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_29
timestamp 1636968456
transform 1 0 3772 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_41
timestamp 1636968456
transform 1 0 4876 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_53
timestamp 1
transform 1 0 5980 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_57
timestamp 1636968456
transform 1 0 6348 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_69
timestamp 1636968456
transform 1 0 7452 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_81
timestamp 1
transform 1 0 8556 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_85
timestamp 1636968456
transform 1 0 8924 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_97
timestamp 1636968456
transform 1 0 10028 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_109
timestamp 1
transform 1 0 11132 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_113
timestamp 1636968456
transform 1 0 11500 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_125
timestamp 1636968456
transform 1 0 12604 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_137
timestamp 1
transform 1 0 13708 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_141
timestamp 1636968456
transform 1 0 14076 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_153
timestamp 1636968456
transform 1 0 15180 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_165
timestamp 1
transform 1 0 16284 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_169
timestamp 1636968456
transform 1 0 16652 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_181
timestamp 1636968456
transform 1 0 17756 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_193
timestamp 1
transform 1 0 18860 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_197
timestamp 1636968456
transform 1 0 19228 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_209
timestamp 1636968456
transform 1 0 20332 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_221
timestamp 1
transform 1 0 21436 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_225
timestamp 1636968456
transform 1 0 21804 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_237
timestamp 1636968456
transform 1 0 22908 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_249
timestamp 1
transform 1 0 24012 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_253
timestamp 1636968456
transform 1 0 24380 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_265
timestamp 1636968456
transform 1 0 25484 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_277
timestamp 1
transform 1 0 26588 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_281
timestamp 1636968456
transform 1 0 26956 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_293
timestamp 1636968456
transform 1 0 28060 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_305
timestamp 1
transform 1 0 29164 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_309
timestamp 1636968456
transform 1 0 29532 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_321
timestamp 1636968456
transform 1 0 30636 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_333
timestamp 1
transform 1 0 31740 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_337
timestamp 1636968456
transform 1 0 32108 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_349
timestamp 1
transform 1 0 33212 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_246_357
timestamp 1
transform 1 0 33948 0 1 136000
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_246_363
timestamp 1
transform 1 0 34500 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_246_367
timestamp 1
transform 1 0 34868 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_246_374
timestamp 1
transform 1 0 35512 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_246_378
timestamp 1
transform 1 0 35880 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_246_385
timestamp 1
transform 1 0 36524 0 1 136000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_246_391
timestamp 1
transform 1 0 37076 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_393
timestamp 1636968456
transform 1 0 37260 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_405
timestamp 1636968456
transform 1 0 38364 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_417
timestamp 1
transform 1 0 39468 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_421
timestamp 1636968456
transform 1 0 39836 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_433
timestamp 1636968456
transform 1 0 40940 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_445
timestamp 1
transform 1 0 42044 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_246_449
timestamp 1
transform 1 0 42412 0 1 136000
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_246_461
timestamp 1636968456
transform 1 0 43516 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_473
timestamp 1
transform 1 0 44620 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_477
timestamp 1636968456
transform 1 0 44988 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_491
timestamp 1636968456
transform 1 0 46276 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_246_503
timestamp 1
transform 1 0 47380 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_511
timestamp 1636968456
transform 1 0 48116 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_523
timestamp 1
transform 1 0 49220 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_531
timestamp 1
transform 1 0 49956 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_539
timestamp 1636968456
transform 1 0 50692 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_551
timestamp 1
transform 1 0 51796 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_559
timestamp 1
transform 1 0 52532 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_561
timestamp 1636968456
transform 1 0 52716 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_573
timestamp 1636968456
transform 1 0 53820 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_585
timestamp 1
transform 1 0 54924 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_595
timestamp 1636968456
transform 1 0 55844 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_607
timestamp 1
transform 1 0 56948 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_615
timestamp 1
transform 1 0 57684 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_623
timestamp 1636968456
transform 1 0 58420 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_635
timestamp 1
transform 1 0 59524 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_643
timestamp 1
transform 1 0 60260 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_651
timestamp 1636968456
transform 1 0 60996 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_663
timestamp 1
transform 1 0 62100 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_671
timestamp 1
transform 1 0 62836 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_681
timestamp 1636968456
transform 1 0 63756 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_246_693
timestamp 1
transform 1 0 64860 0 1 136000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_246_699
timestamp 1
transform 1 0 65412 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_701
timestamp 1636968456
transform 1 0 65596 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_713
timestamp 1636968456
transform 1 0 66700 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_725
timestamp 1
transform 1 0 67804 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_246_729
timestamp 1
transform 1 0 68172 0 1 136000
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_246_735
timestamp 1636968456
transform 1 0 68724 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_747
timestamp 1
transform 1 0 69828 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_755
timestamp 1
transform 1 0 70564 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_757
timestamp 1636968456
transform 1 0 70748 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_246_769
timestamp 1
transform 1 0 71852 0 1 136000
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_246_781
timestamp 1
transform 1 0 72956 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_791
timestamp 1636968456
transform 1 0 73876 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_803
timestamp 1
transform 1 0 74980 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_811
timestamp 1
transform 1 0 75716 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_813
timestamp 1636968456
transform 1 0 75900 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_825
timestamp 1
transform 1 0 77004 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_246_834
timestamp 1
transform 1 0 77832 0 1 136000
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_246_841
timestamp 1636968456
transform 1 0 78476 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_853
timestamp 1636968456
transform 1 0 79580 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_865
timestamp 1
transform 1 0 80684 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_869
timestamp 1636968456
transform 1 0 81052 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_881
timestamp 1636968456
transform 1 0 82156 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_893
timestamp 1
transform 1 0 83260 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_897
timestamp 1636968456
transform 1 0 83628 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_909
timestamp 1636968456
transform 1 0 84732 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_921
timestamp 1
transform 1 0 85836 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_246_927
timestamp 1
transform 1 0 86388 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_246_935
timestamp 1
transform 1 0 87124 0 1 136000
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_246_939
timestamp 1636968456
transform 1 0 87492 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_246_951
timestamp 1
transform 1 0 88596 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_246_953
timestamp 1636968456
transform 1 0 88780 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_965
timestamp 1636968456
transform 1 0 89884 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_977
timestamp 1
transform 1 0 90988 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_981
timestamp 1636968456
transform 1 0 91356 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_993
timestamp 1636968456
transform 1 0 92460 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1005
timestamp 1
transform 1 0 93564 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1009
timestamp 1636968456
transform 1 0 93932 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_246_1021
timestamp 1
transform 1 0 95036 0 1 136000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_246_1029
timestamp 1
transform 1 0 95772 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_246_1032
timestamp 1
transform 1 0 96048 0 1 136000
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1037
timestamp 1636968456
transform 1 0 96508 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1049
timestamp 1636968456
transform 1 0 97612 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1061
timestamp 1
transform 1 0 98716 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1065
timestamp 1636968456
transform 1 0 99084 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1077
timestamp 1636968456
transform 1 0 100188 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1089
timestamp 1
transform 1 0 101292 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1093
timestamp 1636968456
transform 1 0 101660 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1105
timestamp 1636968456
transform 1 0 102764 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1117
timestamp 1
transform 1 0 103868 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1121
timestamp 1636968456
transform 1 0 104236 0 1 136000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1133
timestamp 1636968456
transform 1 0 105340 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_246_1145
timestamp 1
transform 1 0 106444 0 1 136000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_246_1149
timestamp 1636968456
transform 1 0 106812 0 1 136000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_246_1161
timestamp 1
transform 1 0 107916 0 1 136000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_246_1167
timestamp 1
transform 1 0 108468 0 1 136000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_3
timestamp 1636968456
transform 1 0 1380 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_15
timestamp 1636968456
transform 1 0 2484 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_27
timestamp 1636968456
transform 1 0 3588 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_39
timestamp 1636968456
transform 1 0 4692 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_247_51
timestamp 1
transform 1 0 5796 0 -1 137088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_247_55
timestamp 1
transform 1 0 6164 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_57
timestamp 1636968456
transform 1 0 6348 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_69
timestamp 1636968456
transform 1 0 7452 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_81
timestamp 1636968456
transform 1 0 8556 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_93
timestamp 1636968456
transform 1 0 9660 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_105
timestamp 1
transform 1 0 10764 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_111
timestamp 1
transform 1 0 11316 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_113
timestamp 1636968456
transform 1 0 11500 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_125
timestamp 1636968456
transform 1 0 12604 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_137
timestamp 1636968456
transform 1 0 13708 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_149
timestamp 1636968456
transform 1 0 14812 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_161
timestamp 1
transform 1 0 15916 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_167
timestamp 1
transform 1 0 16468 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_169
timestamp 1636968456
transform 1 0 16652 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_181
timestamp 1636968456
transform 1 0 17756 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_193
timestamp 1636968456
transform 1 0 18860 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_205
timestamp 1636968456
transform 1 0 19964 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_217
timestamp 1
transform 1 0 21068 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_223
timestamp 1
transform 1 0 21620 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_225
timestamp 1636968456
transform 1 0 21804 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_237
timestamp 1636968456
transform 1 0 22908 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_249
timestamp 1636968456
transform 1 0 24012 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_261
timestamp 1636968456
transform 1 0 25116 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_273
timestamp 1
transform 1 0 26220 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_279
timestamp 1
transform 1 0 26772 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_281
timestamp 1636968456
transform 1 0 26956 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_293
timestamp 1636968456
transform 1 0 28060 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_305
timestamp 1636968456
transform 1 0 29164 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_317
timestamp 1636968456
transform 1 0 30268 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_329
timestamp 1
transform 1 0 31372 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_335
timestamp 1
transform 1 0 31924 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_337
timestamp 1636968456
transform 1 0 32108 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_349
timestamp 1636968456
transform 1 0 33212 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_361
timestamp 1636968456
transform 1 0 34316 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_373
timestamp 1636968456
transform 1 0 35420 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_385
timestamp 1
transform 1 0 36524 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_391
timestamp 1
transform 1 0 37076 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_393
timestamp 1636968456
transform 1 0 37260 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_405
timestamp 1636968456
transform 1 0 38364 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_417
timestamp 1636968456
transform 1 0 39468 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_429
timestamp 1636968456
transform 1 0 40572 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_441
timestamp 1
transform 1 0 41676 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_447
timestamp 1
transform 1 0 42228 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_449
timestamp 1636968456
transform 1 0 42412 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_461
timestamp 1636968456
transform 1 0 43516 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_473
timestamp 1636968456
transform 1 0 44620 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_485
timestamp 1636968456
transform 1 0 45724 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_497
timestamp 1
transform 1 0 46828 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_503
timestamp 1
transform 1 0 47380 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_505
timestamp 1636968456
transform 1 0 47564 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_517
timestamp 1636968456
transform 1 0 48668 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_529
timestamp 1636968456
transform 1 0 49772 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_541
timestamp 1636968456
transform 1 0 50876 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_553
timestamp 1
transform 1 0 51980 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_559
timestamp 1
transform 1 0 52532 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_561
timestamp 1636968456
transform 1 0 52716 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_573
timestamp 1636968456
transform 1 0 53820 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_585
timestamp 1636968456
transform 1 0 54924 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_597
timestamp 1636968456
transform 1 0 56028 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_609
timestamp 1
transform 1 0 57132 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_615
timestamp 1
transform 1 0 57684 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_617
timestamp 1636968456
transform 1 0 57868 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_629
timestamp 1636968456
transform 1 0 58972 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_641
timestamp 1636968456
transform 1 0 60076 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_653
timestamp 1636968456
transform 1 0 61180 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_665
timestamp 1
transform 1 0 62284 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_671
timestamp 1
transform 1 0 62836 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_673
timestamp 1636968456
transform 1 0 63020 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_685
timestamp 1636968456
transform 1 0 64124 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_697
timestamp 1636968456
transform 1 0 65228 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_709
timestamp 1636968456
transform 1 0 66332 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_721
timestamp 1
transform 1 0 67436 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_727
timestamp 1
transform 1 0 67988 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_729
timestamp 1636968456
transform 1 0 68172 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_741
timestamp 1636968456
transform 1 0 69276 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_753
timestamp 1636968456
transform 1 0 70380 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_765
timestamp 1636968456
transform 1 0 71484 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_777
timestamp 1
transform 1 0 72588 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_783
timestamp 1
transform 1 0 73140 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_785
timestamp 1636968456
transform 1 0 73324 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_797
timestamp 1636968456
transform 1 0 74428 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_809
timestamp 1636968456
transform 1 0 75532 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_821
timestamp 1636968456
transform 1 0 76636 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_833
timestamp 1
transform 1 0 77740 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_839
timestamp 1
transform 1 0 78292 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_841
timestamp 1636968456
transform 1 0 78476 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_853
timestamp 1636968456
transform 1 0 79580 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_865
timestamp 1636968456
transform 1 0 80684 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_877
timestamp 1636968456
transform 1 0 81788 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_889
timestamp 1
transform 1 0 82892 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_895
timestamp 1
transform 1 0 83444 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_920
timestamp 1636968456
transform 1 0 85744 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_932
timestamp 1636968456
transform 1 0 86848 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_247_944
timestamp 1
transform 1 0 87952 0 -1 137088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_247_953
timestamp 1636968456
transform 1 0 88780 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_965
timestamp 1636968456
transform 1 0 89884 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_977
timestamp 1636968456
transform 1 0 90988 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_989
timestamp 1636968456
transform 1 0 92092 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_1001
timestamp 1
transform 1 0 93196 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_1007
timestamp 1
transform 1 0 93748 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1009
timestamp 1636968456
transform 1 0 93932 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1021
timestamp 1636968456
transform 1 0 95036 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1033
timestamp 1636968456
transform 1 0 96140 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1045
timestamp 1636968456
transform 1 0 97244 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_1057
timestamp 1
transform 1 0 98348 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_1063
timestamp 1
transform 1 0 98900 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1065
timestamp 1636968456
transform 1 0 99084 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1077
timestamp 1636968456
transform 1 0 100188 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1089
timestamp 1636968456
transform 1 0 101292 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1101
timestamp 1636968456
transform 1 0 102396 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_247_1113
timestamp 1
transform 1 0 103500 0 -1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_247_1119
timestamp 1
transform 1 0 104052 0 -1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1121
timestamp 1636968456
transform 1 0 104236 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1133
timestamp 1636968456
transform 1 0 105340 0 -1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_247_1145
timestamp 1636968456
transform 1 0 106444 0 -1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_247_1157
timestamp 1
transform 1 0 107548 0 -1 137088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_247_1165
timestamp 1
transform 1 0 108284 0 -1 137088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_248_3
timestamp 1636968456
transform 1 0 1380 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_15
timestamp 1636968456
transform 1 0 2484 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_248_27
timestamp 1
transform 1 0 3588 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_29
timestamp 1636968456
transform 1 0 3772 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_41
timestamp 1636968456
transform 1 0 4876 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_53
timestamp 1636968456
transform 1 0 5980 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_65
timestamp 1636968456
transform 1 0 7084 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_77
timestamp 1
transform 1 0 8188 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_83
timestamp 1
transform 1 0 8740 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_85
timestamp 1636968456
transform 1 0 8924 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_97
timestamp 1636968456
transform 1 0 10028 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_109
timestamp 1636968456
transform 1 0 11132 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_121
timestamp 1636968456
transform 1 0 12236 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_133
timestamp 1
transform 1 0 13340 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_139
timestamp 1
transform 1 0 13892 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_141
timestamp 1636968456
transform 1 0 14076 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_153
timestamp 1636968456
transform 1 0 15180 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_165
timestamp 1636968456
transform 1 0 16284 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_177
timestamp 1636968456
transform 1 0 17388 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_189
timestamp 1
transform 1 0 18492 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_195
timestamp 1
transform 1 0 19044 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_197
timestamp 1636968456
transform 1 0 19228 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_209
timestamp 1636968456
transform 1 0 20332 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_221
timestamp 1636968456
transform 1 0 21436 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_233
timestamp 1636968456
transform 1 0 22540 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_245
timestamp 1
transform 1 0 23644 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_251
timestamp 1
transform 1 0 24196 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_253
timestamp 1636968456
transform 1 0 24380 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_265
timestamp 1636968456
transform 1 0 25484 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_277
timestamp 1636968456
transform 1 0 26588 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_289
timestamp 1636968456
transform 1 0 27692 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_301
timestamp 1
transform 1 0 28796 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_307
timestamp 1
transform 1 0 29348 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_309
timestamp 1636968456
transform 1 0 29532 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_321
timestamp 1636968456
transform 1 0 30636 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_333
timestamp 1636968456
transform 1 0 31740 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_345
timestamp 1636968456
transform 1 0 32844 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_357
timestamp 1
transform 1 0 33948 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_363
timestamp 1
transform 1 0 34500 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_365
timestamp 1636968456
transform 1 0 34684 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_377
timestamp 1636968456
transform 1 0 35788 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_389
timestamp 1636968456
transform 1 0 36892 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_401
timestamp 1636968456
transform 1 0 37996 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_413
timestamp 1
transform 1 0 39100 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_419
timestamp 1
transform 1 0 39652 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_421
timestamp 1636968456
transform 1 0 39836 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_433
timestamp 1636968456
transform 1 0 40940 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_445
timestamp 1636968456
transform 1 0 42044 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_457
timestamp 1636968456
transform 1 0 43148 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_469
timestamp 1
transform 1 0 44252 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_475
timestamp 1
transform 1 0 44804 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_477
timestamp 1636968456
transform 1 0 44988 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_489
timestamp 1636968456
transform 1 0 46092 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_501
timestamp 1636968456
transform 1 0 47196 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_513
timestamp 1636968456
transform 1 0 48300 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_525
timestamp 1
transform 1 0 49404 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_531
timestamp 1
transform 1 0 49956 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_533
timestamp 1636968456
transform 1 0 50140 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_545
timestamp 1636968456
transform 1 0 51244 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_557
timestamp 1636968456
transform 1 0 52348 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_569
timestamp 1636968456
transform 1 0 53452 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_581
timestamp 1
transform 1 0 54556 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_587
timestamp 1
transform 1 0 55108 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_589
timestamp 1636968456
transform 1 0 55292 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_601
timestamp 1636968456
transform 1 0 56396 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_613
timestamp 1636968456
transform 1 0 57500 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_625
timestamp 1636968456
transform 1 0 58604 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_637
timestamp 1
transform 1 0 59708 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_643
timestamp 1
transform 1 0 60260 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_645
timestamp 1636968456
transform 1 0 60444 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_657
timestamp 1636968456
transform 1 0 61548 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_669
timestamp 1636968456
transform 1 0 62652 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_681
timestamp 1636968456
transform 1 0 63756 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_693
timestamp 1
transform 1 0 64860 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_699
timestamp 1
transform 1 0 65412 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_701
timestamp 1636968456
transform 1 0 65596 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_713
timestamp 1636968456
transform 1 0 66700 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_725
timestamp 1636968456
transform 1 0 67804 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_737
timestamp 1636968456
transform 1 0 68908 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_749
timestamp 1
transform 1 0 70012 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_755
timestamp 1
transform 1 0 70564 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_757
timestamp 1636968456
transform 1 0 70748 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_769
timestamp 1636968456
transform 1 0 71852 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_781
timestamp 1636968456
transform 1 0 72956 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_793
timestamp 1636968456
transform 1 0 74060 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_805
timestamp 1
transform 1 0 75164 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_811
timestamp 1
transform 1 0 75716 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_813
timestamp 1636968456
transform 1 0 75900 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_825
timestamp 1636968456
transform 1 0 77004 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_837
timestamp 1636968456
transform 1 0 78108 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_849
timestamp 1636968456
transform 1 0 79212 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_861
timestamp 1
transform 1 0 80316 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_867
timestamp 1
transform 1 0 80868 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_869
timestamp 1636968456
transform 1 0 81052 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_881
timestamp 1636968456
transform 1 0 82156 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_893
timestamp 1636968456
transform 1 0 83260 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_905
timestamp 1636968456
transform 1 0 84364 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_917
timestamp 1
transform 1 0 85468 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_923
timestamp 1
transform 1 0 86020 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_925
timestamp 1636968456
transform 1 0 86204 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_937
timestamp 1636968456
transform 1 0 87308 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_949
timestamp 1636968456
transform 1 0 88412 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_961
timestamp 1636968456
transform 1 0 89516 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_973
timestamp 1
transform 1 0 90620 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_979
timestamp 1
transform 1 0 91172 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_981
timestamp 1636968456
transform 1 0 91356 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_993
timestamp 1636968456
transform 1 0 92460 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1005
timestamp 1636968456
transform 1 0 93564 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1017
timestamp 1636968456
transform 1 0 94668 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_1029
timestamp 1
transform 1 0 95772 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_1035
timestamp 1
transform 1 0 96324 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1037
timestamp 1636968456
transform 1 0 96508 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1049
timestamp 1636968456
transform 1 0 97612 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1061
timestamp 1636968456
transform 1 0 98716 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1073
timestamp 1636968456
transform 1 0 99820 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_1085
timestamp 1
transform 1 0 100924 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_1091
timestamp 1
transform 1 0 101476 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1093
timestamp 1636968456
transform 1 0 101660 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1105
timestamp 1636968456
transform 1 0 102764 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1117
timestamp 1636968456
transform 1 0 103868 0 1 137088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1129
timestamp 1636968456
transform 1 0 104972 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_1141
timestamp 1
transform 1 0 106076 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_1147
timestamp 1
transform 1 0 106628 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_248_1149
timestamp 1636968456
transform 1 0 106812 0 1 137088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_248_1161
timestamp 1
transform 1 0 107916 0 1 137088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_248_1167
timestamp 1
transform 1 0 108468 0 1 137088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_3
timestamp 1636968456
transform 1 0 1380 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_15
timestamp 1636968456
transform 1 0 2484 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_27
timestamp 1636968456
transform 1 0 3588 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_39
timestamp 1636968456
transform 1 0 4692 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_249_51
timestamp 1
transform 1 0 5796 0 -1 138176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_249_55
timestamp 1
transform 1 0 6164 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_57
timestamp 1636968456
transform 1 0 6348 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_69
timestamp 1636968456
transform 1 0 7452 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_81
timestamp 1636968456
transform 1 0 8556 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_93
timestamp 1636968456
transform 1 0 9660 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_105
timestamp 1
transform 1 0 10764 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_111
timestamp 1
transform 1 0 11316 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_113
timestamp 1636968456
transform 1 0 11500 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_125
timestamp 1636968456
transform 1 0 12604 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_137
timestamp 1636968456
transform 1 0 13708 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_149
timestamp 1636968456
transform 1 0 14812 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_161
timestamp 1
transform 1 0 15916 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_167
timestamp 1
transform 1 0 16468 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_169
timestamp 1636968456
transform 1 0 16652 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_181
timestamp 1636968456
transform 1 0 17756 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_193
timestamp 1636968456
transform 1 0 18860 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_205
timestamp 1636968456
transform 1 0 19964 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_217
timestamp 1
transform 1 0 21068 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_223
timestamp 1
transform 1 0 21620 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_225
timestamp 1636968456
transform 1 0 21804 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_237
timestamp 1636968456
transform 1 0 22908 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_249
timestamp 1636968456
transform 1 0 24012 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_261
timestamp 1636968456
transform 1 0 25116 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_273
timestamp 1
transform 1 0 26220 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_279
timestamp 1
transform 1 0 26772 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_281
timestamp 1636968456
transform 1 0 26956 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_293
timestamp 1636968456
transform 1 0 28060 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_305
timestamp 1636968456
transform 1 0 29164 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_317
timestamp 1636968456
transform 1 0 30268 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_329
timestamp 1
transform 1 0 31372 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_335
timestamp 1
transform 1 0 31924 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_337
timestamp 1636968456
transform 1 0 32108 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_349
timestamp 1636968456
transform 1 0 33212 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_361
timestamp 1636968456
transform 1 0 34316 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_373
timestamp 1636968456
transform 1 0 35420 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_385
timestamp 1
transform 1 0 36524 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_391
timestamp 1
transform 1 0 37076 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_393
timestamp 1636968456
transform 1 0 37260 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_405
timestamp 1636968456
transform 1 0 38364 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_417
timestamp 1636968456
transform 1 0 39468 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_429
timestamp 1636968456
transform 1 0 40572 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_441
timestamp 1
transform 1 0 41676 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_447
timestamp 1
transform 1 0 42228 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_449
timestamp 1636968456
transform 1 0 42412 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_461
timestamp 1636968456
transform 1 0 43516 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_473
timestamp 1636968456
transform 1 0 44620 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_485
timestamp 1636968456
transform 1 0 45724 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_497
timestamp 1
transform 1 0 46828 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_503
timestamp 1
transform 1 0 47380 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_505
timestamp 1636968456
transform 1 0 47564 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_517
timestamp 1636968456
transform 1 0 48668 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_529
timestamp 1636968456
transform 1 0 49772 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_541
timestamp 1636968456
transform 1 0 50876 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_553
timestamp 1
transform 1 0 51980 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_559
timestamp 1
transform 1 0 52532 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_561
timestamp 1636968456
transform 1 0 52716 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_573
timestamp 1636968456
transform 1 0 53820 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_585
timestamp 1636968456
transform 1 0 54924 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_597
timestamp 1636968456
transform 1 0 56028 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_609
timestamp 1
transform 1 0 57132 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_615
timestamp 1
transform 1 0 57684 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_617
timestamp 1636968456
transform 1 0 57868 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_629
timestamp 1636968456
transform 1 0 58972 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_641
timestamp 1636968456
transform 1 0 60076 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_653
timestamp 1636968456
transform 1 0 61180 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_665
timestamp 1
transform 1 0 62284 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_671
timestamp 1
transform 1 0 62836 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_673
timestamp 1636968456
transform 1 0 63020 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_685
timestamp 1636968456
transform 1 0 64124 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_697
timestamp 1636968456
transform 1 0 65228 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_709
timestamp 1636968456
transform 1 0 66332 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_721
timestamp 1
transform 1 0 67436 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_727
timestamp 1
transform 1 0 67988 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_729
timestamp 1636968456
transform 1 0 68172 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_741
timestamp 1636968456
transform 1 0 69276 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_753
timestamp 1636968456
transform 1 0 70380 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_765
timestamp 1636968456
transform 1 0 71484 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_777
timestamp 1
transform 1 0 72588 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_783
timestamp 1
transform 1 0 73140 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_785
timestamp 1636968456
transform 1 0 73324 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_797
timestamp 1636968456
transform 1 0 74428 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_809
timestamp 1636968456
transform 1 0 75532 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_821
timestamp 1636968456
transform 1 0 76636 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_833
timestamp 1
transform 1 0 77740 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_839
timestamp 1
transform 1 0 78292 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_841
timestamp 1636968456
transform 1 0 78476 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_853
timestamp 1636968456
transform 1 0 79580 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_865
timestamp 1636968456
transform 1 0 80684 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_877
timestamp 1636968456
transform 1 0 81788 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_889
timestamp 1
transform 1 0 82892 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_895
timestamp 1
transform 1 0 83444 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_897
timestamp 1636968456
transform 1 0 83628 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_909
timestamp 1636968456
transform 1 0 84732 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_921
timestamp 1636968456
transform 1 0 85836 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_933
timestamp 1636968456
transform 1 0 86940 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_945
timestamp 1
transform 1 0 88044 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_951
timestamp 1
transform 1 0 88596 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_953
timestamp 1636968456
transform 1 0 88780 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_965
timestamp 1636968456
transform 1 0 89884 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_977
timestamp 1636968456
transform 1 0 90988 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_989
timestamp 1636968456
transform 1 0 92092 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_1001
timestamp 1
transform 1 0 93196 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_1007
timestamp 1
transform 1 0 93748 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1009
timestamp 1636968456
transform 1 0 93932 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1021
timestamp 1636968456
transform 1 0 95036 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1033
timestamp 1636968456
transform 1 0 96140 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1045
timestamp 1636968456
transform 1 0 97244 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_1057
timestamp 1
transform 1 0 98348 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_1063
timestamp 1
transform 1 0 98900 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1065
timestamp 1636968456
transform 1 0 99084 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1077
timestamp 1636968456
transform 1 0 100188 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1089
timestamp 1636968456
transform 1 0 101292 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1101
timestamp 1636968456
transform 1 0 102396 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_249_1113
timestamp 1
transform 1 0 103500 0 -1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_249_1119
timestamp 1
transform 1 0 104052 0 -1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1121
timestamp 1636968456
transform 1 0 104236 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1133
timestamp 1636968456
transform 1 0 105340 0 -1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_249_1145
timestamp 1636968456
transform 1 0 106444 0 -1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_249_1157
timestamp 1
transform 1 0 107548 0 -1 138176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_249_1165
timestamp 1
transform 1 0 108284 0 -1 138176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_250_3
timestamp 1636968456
transform 1 0 1380 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_15
timestamp 1636968456
transform 1 0 2484 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_250_27
timestamp 1
transform 1 0 3588 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_29
timestamp 1636968456
transform 1 0 3772 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_41
timestamp 1636968456
transform 1 0 4876 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_53
timestamp 1636968456
transform 1 0 5980 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_65
timestamp 1636968456
transform 1 0 7084 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_77
timestamp 1
transform 1 0 8188 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_83
timestamp 1
transform 1 0 8740 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_85
timestamp 1636968456
transform 1 0 8924 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_97
timestamp 1636968456
transform 1 0 10028 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_109
timestamp 1636968456
transform 1 0 11132 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_121
timestamp 1636968456
transform 1 0 12236 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_133
timestamp 1
transform 1 0 13340 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_139
timestamp 1
transform 1 0 13892 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_141
timestamp 1636968456
transform 1 0 14076 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_153
timestamp 1636968456
transform 1 0 15180 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_165
timestamp 1636968456
transform 1 0 16284 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_177
timestamp 1636968456
transform 1 0 17388 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_189
timestamp 1
transform 1 0 18492 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_195
timestamp 1
transform 1 0 19044 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_197
timestamp 1636968456
transform 1 0 19228 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_209
timestamp 1636968456
transform 1 0 20332 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_221
timestamp 1636968456
transform 1 0 21436 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_233
timestamp 1636968456
transform 1 0 22540 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_245
timestamp 1
transform 1 0 23644 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_251
timestamp 1
transform 1 0 24196 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_253
timestamp 1636968456
transform 1 0 24380 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_265
timestamp 1636968456
transform 1 0 25484 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_277
timestamp 1636968456
transform 1 0 26588 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_289
timestamp 1636968456
transform 1 0 27692 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_301
timestamp 1
transform 1 0 28796 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_307
timestamp 1
transform 1 0 29348 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_309
timestamp 1636968456
transform 1 0 29532 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_321
timestamp 1636968456
transform 1 0 30636 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_333
timestamp 1636968456
transform 1 0 31740 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_345
timestamp 1636968456
transform 1 0 32844 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_357
timestamp 1
transform 1 0 33948 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_363
timestamp 1
transform 1 0 34500 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_365
timestamp 1636968456
transform 1 0 34684 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_377
timestamp 1636968456
transform 1 0 35788 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_389
timestamp 1636968456
transform 1 0 36892 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_401
timestamp 1636968456
transform 1 0 37996 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_413
timestamp 1
transform 1 0 39100 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_419
timestamp 1
transform 1 0 39652 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_421
timestamp 1636968456
transform 1 0 39836 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_433
timestamp 1636968456
transform 1 0 40940 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_445
timestamp 1636968456
transform 1 0 42044 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_457
timestamp 1636968456
transform 1 0 43148 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_469
timestamp 1
transform 1 0 44252 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_475
timestamp 1
transform 1 0 44804 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_477
timestamp 1636968456
transform 1 0 44988 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_489
timestamp 1636968456
transform 1 0 46092 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_501
timestamp 1636968456
transform 1 0 47196 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_513
timestamp 1636968456
transform 1 0 48300 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_525
timestamp 1
transform 1 0 49404 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_531
timestamp 1
transform 1 0 49956 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_533
timestamp 1636968456
transform 1 0 50140 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_545
timestamp 1636968456
transform 1 0 51244 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_557
timestamp 1636968456
transform 1 0 52348 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_569
timestamp 1636968456
transform 1 0 53452 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_581
timestamp 1
transform 1 0 54556 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_587
timestamp 1
transform 1 0 55108 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_589
timestamp 1636968456
transform 1 0 55292 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_601
timestamp 1636968456
transform 1 0 56396 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_613
timestamp 1636968456
transform 1 0 57500 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_625
timestamp 1636968456
transform 1 0 58604 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_637
timestamp 1
transform 1 0 59708 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_643
timestamp 1
transform 1 0 60260 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_645
timestamp 1636968456
transform 1 0 60444 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_657
timestamp 1636968456
transform 1 0 61548 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_669
timestamp 1636968456
transform 1 0 62652 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_681
timestamp 1636968456
transform 1 0 63756 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_693
timestamp 1
transform 1 0 64860 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_699
timestamp 1
transform 1 0 65412 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_701
timestamp 1636968456
transform 1 0 65596 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_713
timestamp 1636968456
transform 1 0 66700 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_725
timestamp 1636968456
transform 1 0 67804 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_737
timestamp 1636968456
transform 1 0 68908 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_749
timestamp 1
transform 1 0 70012 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_755
timestamp 1
transform 1 0 70564 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_757
timestamp 1636968456
transform 1 0 70748 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_769
timestamp 1636968456
transform 1 0 71852 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_781
timestamp 1636968456
transform 1 0 72956 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_793
timestamp 1636968456
transform 1 0 74060 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_805
timestamp 1
transform 1 0 75164 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_811
timestamp 1
transform 1 0 75716 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_813
timestamp 1636968456
transform 1 0 75900 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_825
timestamp 1636968456
transform 1 0 77004 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_837
timestamp 1636968456
transform 1 0 78108 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_849
timestamp 1636968456
transform 1 0 79212 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_861
timestamp 1
transform 1 0 80316 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_867
timestamp 1
transform 1 0 80868 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_869
timestamp 1636968456
transform 1 0 81052 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_881
timestamp 1636968456
transform 1 0 82156 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_893
timestamp 1636968456
transform 1 0 83260 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_905
timestamp 1636968456
transform 1 0 84364 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_917
timestamp 1
transform 1 0 85468 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_923
timestamp 1
transform 1 0 86020 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_925
timestamp 1636968456
transform 1 0 86204 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_937
timestamp 1636968456
transform 1 0 87308 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_949
timestamp 1636968456
transform 1 0 88412 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_961
timestamp 1636968456
transform 1 0 89516 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_973
timestamp 1
transform 1 0 90620 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_979
timestamp 1
transform 1 0 91172 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_981
timestamp 1636968456
transform 1 0 91356 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_993
timestamp 1636968456
transform 1 0 92460 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1005
timestamp 1636968456
transform 1 0 93564 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1017
timestamp 1636968456
transform 1 0 94668 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_1029
timestamp 1
transform 1 0 95772 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_1035
timestamp 1
transform 1 0 96324 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1037
timestamp 1636968456
transform 1 0 96508 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1049
timestamp 1636968456
transform 1 0 97612 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1061
timestamp 1636968456
transform 1 0 98716 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1073
timestamp 1636968456
transform 1 0 99820 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_1085
timestamp 1
transform 1 0 100924 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_1091
timestamp 1
transform 1 0 101476 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1093
timestamp 1636968456
transform 1 0 101660 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1105
timestamp 1636968456
transform 1 0 102764 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1117
timestamp 1636968456
transform 1 0 103868 0 1 138176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1129
timestamp 1636968456
transform 1 0 104972 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_1141
timestamp 1
transform 1 0 106076 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_1147
timestamp 1
transform 1 0 106628 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_250_1149
timestamp 1636968456
transform 1 0 106812 0 1 138176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_250_1161
timestamp 1
transform 1 0 107916 0 1 138176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_250_1167
timestamp 1
transform 1 0 108468 0 1 138176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_3
timestamp 1636968456
transform 1 0 1380 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_15
timestamp 1636968456
transform 1 0 2484 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_27
timestamp 1636968456
transform 1 0 3588 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_39
timestamp 1636968456
transform 1 0 4692 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_251_51
timestamp 1
transform 1 0 5796 0 -1 139264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_251_55
timestamp 1
transform 1 0 6164 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_57
timestamp 1636968456
transform 1 0 6348 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_69
timestamp 1636968456
transform 1 0 7452 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_81
timestamp 1636968456
transform 1 0 8556 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_93
timestamp 1636968456
transform 1 0 9660 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_105
timestamp 1
transform 1 0 10764 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_111
timestamp 1
transform 1 0 11316 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_113
timestamp 1636968456
transform 1 0 11500 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_125
timestamp 1636968456
transform 1 0 12604 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_137
timestamp 1636968456
transform 1 0 13708 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_149
timestamp 1636968456
transform 1 0 14812 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_161
timestamp 1
transform 1 0 15916 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_167
timestamp 1
transform 1 0 16468 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_169
timestamp 1636968456
transform 1 0 16652 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_181
timestamp 1636968456
transform 1 0 17756 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_193
timestamp 1636968456
transform 1 0 18860 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_205
timestamp 1636968456
transform 1 0 19964 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_217
timestamp 1
transform 1 0 21068 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_223
timestamp 1
transform 1 0 21620 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_225
timestamp 1636968456
transform 1 0 21804 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_237
timestamp 1636968456
transform 1 0 22908 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_249
timestamp 1636968456
transform 1 0 24012 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_261
timestamp 1636968456
transform 1 0 25116 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_273
timestamp 1
transform 1 0 26220 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_279
timestamp 1
transform 1 0 26772 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_281
timestamp 1636968456
transform 1 0 26956 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_293
timestamp 1636968456
transform 1 0 28060 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_305
timestamp 1636968456
transform 1 0 29164 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_317
timestamp 1636968456
transform 1 0 30268 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_329
timestamp 1
transform 1 0 31372 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_335
timestamp 1
transform 1 0 31924 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_337
timestamp 1636968456
transform 1 0 32108 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_349
timestamp 1636968456
transform 1 0 33212 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_361
timestamp 1636968456
transform 1 0 34316 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_373
timestamp 1636968456
transform 1 0 35420 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_385
timestamp 1
transform 1 0 36524 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_391
timestamp 1
transform 1 0 37076 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_393
timestamp 1636968456
transform 1 0 37260 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_405
timestamp 1636968456
transform 1 0 38364 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_417
timestamp 1636968456
transform 1 0 39468 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_429
timestamp 1636968456
transform 1 0 40572 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_441
timestamp 1
transform 1 0 41676 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_447
timestamp 1
transform 1 0 42228 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_449
timestamp 1636968456
transform 1 0 42412 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_461
timestamp 1636968456
transform 1 0 43516 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_473
timestamp 1636968456
transform 1 0 44620 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_485
timestamp 1636968456
transform 1 0 45724 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_497
timestamp 1
transform 1 0 46828 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_503
timestamp 1
transform 1 0 47380 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_505
timestamp 1636968456
transform 1 0 47564 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_517
timestamp 1636968456
transform 1 0 48668 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_529
timestamp 1636968456
transform 1 0 49772 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_541
timestamp 1636968456
transform 1 0 50876 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_553
timestamp 1
transform 1 0 51980 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_559
timestamp 1
transform 1 0 52532 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_561
timestamp 1636968456
transform 1 0 52716 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_573
timestamp 1636968456
transform 1 0 53820 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_585
timestamp 1636968456
transform 1 0 54924 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_597
timestamp 1636968456
transform 1 0 56028 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_609
timestamp 1
transform 1 0 57132 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_615
timestamp 1
transform 1 0 57684 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_617
timestamp 1636968456
transform 1 0 57868 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_629
timestamp 1636968456
transform 1 0 58972 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_641
timestamp 1636968456
transform 1 0 60076 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_653
timestamp 1636968456
transform 1 0 61180 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_665
timestamp 1
transform 1 0 62284 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_671
timestamp 1
transform 1 0 62836 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_673
timestamp 1636968456
transform 1 0 63020 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_685
timestamp 1636968456
transform 1 0 64124 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_697
timestamp 1636968456
transform 1 0 65228 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_709
timestamp 1636968456
transform 1 0 66332 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_721
timestamp 1
transform 1 0 67436 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_727
timestamp 1
transform 1 0 67988 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_729
timestamp 1636968456
transform 1 0 68172 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_741
timestamp 1636968456
transform 1 0 69276 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_753
timestamp 1636968456
transform 1 0 70380 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_765
timestamp 1636968456
transform 1 0 71484 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_777
timestamp 1
transform 1 0 72588 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_783
timestamp 1
transform 1 0 73140 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_785
timestamp 1636968456
transform 1 0 73324 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_797
timestamp 1636968456
transform 1 0 74428 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_809
timestamp 1636968456
transform 1 0 75532 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_821
timestamp 1636968456
transform 1 0 76636 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_833
timestamp 1
transform 1 0 77740 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_839
timestamp 1
transform 1 0 78292 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_841
timestamp 1636968456
transform 1 0 78476 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_853
timestamp 1636968456
transform 1 0 79580 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_865
timestamp 1636968456
transform 1 0 80684 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_877
timestamp 1636968456
transform 1 0 81788 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_889
timestamp 1
transform 1 0 82892 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_895
timestamp 1
transform 1 0 83444 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_897
timestamp 1636968456
transform 1 0 83628 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_909
timestamp 1636968456
transform 1 0 84732 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_921
timestamp 1636968456
transform 1 0 85836 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_933
timestamp 1636968456
transform 1 0 86940 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_945
timestamp 1
transform 1 0 88044 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_951
timestamp 1
transform 1 0 88596 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_953
timestamp 1636968456
transform 1 0 88780 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_965
timestamp 1636968456
transform 1 0 89884 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_977
timestamp 1636968456
transform 1 0 90988 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_989
timestamp 1636968456
transform 1 0 92092 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_1001
timestamp 1
transform 1 0 93196 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_1007
timestamp 1
transform 1 0 93748 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1009
timestamp 1636968456
transform 1 0 93932 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1021
timestamp 1636968456
transform 1 0 95036 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1033
timestamp 1636968456
transform 1 0 96140 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1045
timestamp 1636968456
transform 1 0 97244 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_1057
timestamp 1
transform 1 0 98348 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_1063
timestamp 1
transform 1 0 98900 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1065
timestamp 1636968456
transform 1 0 99084 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1077
timestamp 1636968456
transform 1 0 100188 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1089
timestamp 1636968456
transform 1 0 101292 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1101
timestamp 1636968456
transform 1 0 102396 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_251_1113
timestamp 1
transform 1 0 103500 0 -1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_251_1119
timestamp 1
transform 1 0 104052 0 -1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1121
timestamp 1636968456
transform 1 0 104236 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1133
timestamp 1636968456
transform 1 0 105340 0 -1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_251_1145
timestamp 1636968456
transform 1 0 106444 0 -1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_251_1157
timestamp 1
transform 1 0 107548 0 -1 139264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_251_1165
timestamp 1
transform 1 0 108284 0 -1 139264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_252_3
timestamp 1636968456
transform 1 0 1380 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_15
timestamp 1636968456
transform 1 0 2484 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_252_27
timestamp 1
transform 1 0 3588 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_29
timestamp 1636968456
transform 1 0 3772 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_41
timestamp 1636968456
transform 1 0 4876 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_53
timestamp 1636968456
transform 1 0 5980 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_65
timestamp 1636968456
transform 1 0 7084 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_77
timestamp 1
transform 1 0 8188 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_83
timestamp 1
transform 1 0 8740 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_85
timestamp 1636968456
transform 1 0 8924 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_97
timestamp 1636968456
transform 1 0 10028 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_109
timestamp 1636968456
transform 1 0 11132 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_121
timestamp 1636968456
transform 1 0 12236 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_133
timestamp 1
transform 1 0 13340 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_139
timestamp 1
transform 1 0 13892 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_141
timestamp 1636968456
transform 1 0 14076 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_153
timestamp 1636968456
transform 1 0 15180 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_165
timestamp 1636968456
transform 1 0 16284 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_177
timestamp 1636968456
transform 1 0 17388 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_189
timestamp 1
transform 1 0 18492 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_195
timestamp 1
transform 1 0 19044 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_197
timestamp 1636968456
transform 1 0 19228 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_209
timestamp 1636968456
transform 1 0 20332 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_221
timestamp 1636968456
transform 1 0 21436 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_233
timestamp 1636968456
transform 1 0 22540 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_245
timestamp 1
transform 1 0 23644 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_251
timestamp 1
transform 1 0 24196 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_253
timestamp 1636968456
transform 1 0 24380 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_265
timestamp 1636968456
transform 1 0 25484 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_277
timestamp 1636968456
transform 1 0 26588 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_289
timestamp 1636968456
transform 1 0 27692 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_301
timestamp 1
transform 1 0 28796 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_307
timestamp 1
transform 1 0 29348 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_309
timestamp 1636968456
transform 1 0 29532 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_321
timestamp 1636968456
transform 1 0 30636 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_333
timestamp 1636968456
transform 1 0 31740 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_345
timestamp 1636968456
transform 1 0 32844 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_357
timestamp 1
transform 1 0 33948 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_363
timestamp 1
transform 1 0 34500 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_365
timestamp 1636968456
transform 1 0 34684 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_377
timestamp 1636968456
transform 1 0 35788 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_389
timestamp 1636968456
transform 1 0 36892 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_401
timestamp 1636968456
transform 1 0 37996 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_413
timestamp 1
transform 1 0 39100 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_419
timestamp 1
transform 1 0 39652 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_421
timestamp 1636968456
transform 1 0 39836 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_433
timestamp 1636968456
transform 1 0 40940 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_445
timestamp 1636968456
transform 1 0 42044 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_457
timestamp 1636968456
transform 1 0 43148 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_469
timestamp 1
transform 1 0 44252 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_475
timestamp 1
transform 1 0 44804 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_477
timestamp 1636968456
transform 1 0 44988 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_489
timestamp 1636968456
transform 1 0 46092 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_501
timestamp 1636968456
transform 1 0 47196 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_513
timestamp 1636968456
transform 1 0 48300 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_525
timestamp 1
transform 1 0 49404 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_531
timestamp 1
transform 1 0 49956 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_533
timestamp 1636968456
transform 1 0 50140 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_545
timestamp 1636968456
transform 1 0 51244 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_557
timestamp 1636968456
transform 1 0 52348 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_569
timestamp 1636968456
transform 1 0 53452 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_581
timestamp 1
transform 1 0 54556 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_587
timestamp 1
transform 1 0 55108 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_589
timestamp 1636968456
transform 1 0 55292 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_601
timestamp 1636968456
transform 1 0 56396 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_613
timestamp 1636968456
transform 1 0 57500 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_625
timestamp 1636968456
transform 1 0 58604 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_637
timestamp 1
transform 1 0 59708 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_643
timestamp 1
transform 1 0 60260 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_645
timestamp 1636968456
transform 1 0 60444 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_657
timestamp 1636968456
transform 1 0 61548 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_669
timestamp 1636968456
transform 1 0 62652 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_681
timestamp 1636968456
transform 1 0 63756 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_693
timestamp 1
transform 1 0 64860 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_699
timestamp 1
transform 1 0 65412 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_701
timestamp 1636968456
transform 1 0 65596 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_713
timestamp 1636968456
transform 1 0 66700 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_725
timestamp 1636968456
transform 1 0 67804 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_737
timestamp 1636968456
transform 1 0 68908 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_749
timestamp 1
transform 1 0 70012 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_755
timestamp 1
transform 1 0 70564 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_757
timestamp 1636968456
transform 1 0 70748 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_769
timestamp 1636968456
transform 1 0 71852 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_781
timestamp 1636968456
transform 1 0 72956 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_793
timestamp 1636968456
transform 1 0 74060 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_805
timestamp 1
transform 1 0 75164 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_811
timestamp 1
transform 1 0 75716 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_813
timestamp 1636968456
transform 1 0 75900 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_825
timestamp 1636968456
transform 1 0 77004 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_837
timestamp 1636968456
transform 1 0 78108 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_849
timestamp 1636968456
transform 1 0 79212 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_861
timestamp 1
transform 1 0 80316 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_867
timestamp 1
transform 1 0 80868 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_869
timestamp 1636968456
transform 1 0 81052 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_881
timestamp 1636968456
transform 1 0 82156 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_893
timestamp 1636968456
transform 1 0 83260 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_905
timestamp 1636968456
transform 1 0 84364 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_917
timestamp 1
transform 1 0 85468 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_923
timestamp 1
transform 1 0 86020 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_925
timestamp 1636968456
transform 1 0 86204 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_937
timestamp 1636968456
transform 1 0 87308 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_949
timestamp 1636968456
transform 1 0 88412 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_961
timestamp 1636968456
transform 1 0 89516 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_973
timestamp 1
transform 1 0 90620 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_979
timestamp 1
transform 1 0 91172 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_981
timestamp 1636968456
transform 1 0 91356 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_993
timestamp 1636968456
transform 1 0 92460 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1005
timestamp 1636968456
transform 1 0 93564 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1017
timestamp 1636968456
transform 1 0 94668 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_1029
timestamp 1
transform 1 0 95772 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_1035
timestamp 1
transform 1 0 96324 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1037
timestamp 1636968456
transform 1 0 96508 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1049
timestamp 1636968456
transform 1 0 97612 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1061
timestamp 1636968456
transform 1 0 98716 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1073
timestamp 1636968456
transform 1 0 99820 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_1085
timestamp 1
transform 1 0 100924 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_1091
timestamp 1
transform 1 0 101476 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1093
timestamp 1636968456
transform 1 0 101660 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1105
timestamp 1636968456
transform 1 0 102764 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1117
timestamp 1636968456
transform 1 0 103868 0 1 139264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1129
timestamp 1636968456
transform 1 0 104972 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_1141
timestamp 1
transform 1 0 106076 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_1147
timestamp 1
transform 1 0 106628 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_252_1149
timestamp 1636968456
transform 1 0 106812 0 1 139264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_252_1161
timestamp 1
transform 1 0 107916 0 1 139264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_252_1167
timestamp 1
transform 1 0 108468 0 1 139264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_3
timestamp 1636968456
transform 1 0 1380 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_15
timestamp 1636968456
transform 1 0 2484 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_27
timestamp 1636968456
transform 1 0 3588 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_39
timestamp 1636968456
transform 1 0 4692 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_253_51
timestamp 1
transform 1 0 5796 0 -1 140352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_253_55
timestamp 1
transform 1 0 6164 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_57
timestamp 1636968456
transform 1 0 6348 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_69
timestamp 1636968456
transform 1 0 7452 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_81
timestamp 1636968456
transform 1 0 8556 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_93
timestamp 1636968456
transform 1 0 9660 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_105
timestamp 1
transform 1 0 10764 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_111
timestamp 1
transform 1 0 11316 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_113
timestamp 1636968456
transform 1 0 11500 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_125
timestamp 1636968456
transform 1 0 12604 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_137
timestamp 1636968456
transform 1 0 13708 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_149
timestamp 1636968456
transform 1 0 14812 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_161
timestamp 1
transform 1 0 15916 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_167
timestamp 1
transform 1 0 16468 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_169
timestamp 1636968456
transform 1 0 16652 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_181
timestamp 1636968456
transform 1 0 17756 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_193
timestamp 1636968456
transform 1 0 18860 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_205
timestamp 1636968456
transform 1 0 19964 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_217
timestamp 1
transform 1 0 21068 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_223
timestamp 1
transform 1 0 21620 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_225
timestamp 1636968456
transform 1 0 21804 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_237
timestamp 1636968456
transform 1 0 22908 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_249
timestamp 1636968456
transform 1 0 24012 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_261
timestamp 1636968456
transform 1 0 25116 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_273
timestamp 1
transform 1 0 26220 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_279
timestamp 1
transform 1 0 26772 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_281
timestamp 1636968456
transform 1 0 26956 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_293
timestamp 1636968456
transform 1 0 28060 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_305
timestamp 1636968456
transform 1 0 29164 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_317
timestamp 1636968456
transform 1 0 30268 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_329
timestamp 1
transform 1 0 31372 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_335
timestamp 1
transform 1 0 31924 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_337
timestamp 1636968456
transform 1 0 32108 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_349
timestamp 1636968456
transform 1 0 33212 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_361
timestamp 1636968456
transform 1 0 34316 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_373
timestamp 1636968456
transform 1 0 35420 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_385
timestamp 1
transform 1 0 36524 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_391
timestamp 1
transform 1 0 37076 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_393
timestamp 1636968456
transform 1 0 37260 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_405
timestamp 1636968456
transform 1 0 38364 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_417
timestamp 1636968456
transform 1 0 39468 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_429
timestamp 1636968456
transform 1 0 40572 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_441
timestamp 1
transform 1 0 41676 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_447
timestamp 1
transform 1 0 42228 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_449
timestamp 1636968456
transform 1 0 42412 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_461
timestamp 1636968456
transform 1 0 43516 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_473
timestamp 1636968456
transform 1 0 44620 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_485
timestamp 1636968456
transform 1 0 45724 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_497
timestamp 1
transform 1 0 46828 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_503
timestamp 1
transform 1 0 47380 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_505
timestamp 1636968456
transform 1 0 47564 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_517
timestamp 1636968456
transform 1 0 48668 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_529
timestamp 1636968456
transform 1 0 49772 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_541
timestamp 1636968456
transform 1 0 50876 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_553
timestamp 1
transform 1 0 51980 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_559
timestamp 1
transform 1 0 52532 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_561
timestamp 1636968456
transform 1 0 52716 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_573
timestamp 1636968456
transform 1 0 53820 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_585
timestamp 1636968456
transform 1 0 54924 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_597
timestamp 1636968456
transform 1 0 56028 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_609
timestamp 1
transform 1 0 57132 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_615
timestamp 1
transform 1 0 57684 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_617
timestamp 1636968456
transform 1 0 57868 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_629
timestamp 1636968456
transform 1 0 58972 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_641
timestamp 1636968456
transform 1 0 60076 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_653
timestamp 1636968456
transform 1 0 61180 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_665
timestamp 1
transform 1 0 62284 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_671
timestamp 1
transform 1 0 62836 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_673
timestamp 1636968456
transform 1 0 63020 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_685
timestamp 1636968456
transform 1 0 64124 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_697
timestamp 1636968456
transform 1 0 65228 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_709
timestamp 1636968456
transform 1 0 66332 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_721
timestamp 1
transform 1 0 67436 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_727
timestamp 1
transform 1 0 67988 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_729
timestamp 1636968456
transform 1 0 68172 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_741
timestamp 1636968456
transform 1 0 69276 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_753
timestamp 1636968456
transform 1 0 70380 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_765
timestamp 1636968456
transform 1 0 71484 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_777
timestamp 1
transform 1 0 72588 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_783
timestamp 1
transform 1 0 73140 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_785
timestamp 1636968456
transform 1 0 73324 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_797
timestamp 1636968456
transform 1 0 74428 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_809
timestamp 1636968456
transform 1 0 75532 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_821
timestamp 1636968456
transform 1 0 76636 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_833
timestamp 1
transform 1 0 77740 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_839
timestamp 1
transform 1 0 78292 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_841
timestamp 1636968456
transform 1 0 78476 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_853
timestamp 1636968456
transform 1 0 79580 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_865
timestamp 1636968456
transform 1 0 80684 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_877
timestamp 1636968456
transform 1 0 81788 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_889
timestamp 1
transform 1 0 82892 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_895
timestamp 1
transform 1 0 83444 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_897
timestamp 1636968456
transform 1 0 83628 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_909
timestamp 1636968456
transform 1 0 84732 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_921
timestamp 1636968456
transform 1 0 85836 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_933
timestamp 1636968456
transform 1 0 86940 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_945
timestamp 1
transform 1 0 88044 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_951
timestamp 1
transform 1 0 88596 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_953
timestamp 1636968456
transform 1 0 88780 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_965
timestamp 1636968456
transform 1 0 89884 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_977
timestamp 1636968456
transform 1 0 90988 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_989
timestamp 1636968456
transform 1 0 92092 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_1001
timestamp 1
transform 1 0 93196 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_1007
timestamp 1
transform 1 0 93748 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1009
timestamp 1636968456
transform 1 0 93932 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1021
timestamp 1636968456
transform 1 0 95036 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1033
timestamp 1636968456
transform 1 0 96140 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1045
timestamp 1636968456
transform 1 0 97244 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_1057
timestamp 1
transform 1 0 98348 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_1063
timestamp 1
transform 1 0 98900 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1065
timestamp 1636968456
transform 1 0 99084 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1077
timestamp 1636968456
transform 1 0 100188 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1089
timestamp 1636968456
transform 1 0 101292 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1101
timestamp 1636968456
transform 1 0 102396 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_253_1113
timestamp 1
transform 1 0 103500 0 -1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_253_1119
timestamp 1
transform 1 0 104052 0 -1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1121
timestamp 1636968456
transform 1 0 104236 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1133
timestamp 1636968456
transform 1 0 105340 0 -1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_253_1145
timestamp 1636968456
transform 1 0 106444 0 -1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_253_1157
timestamp 1
transform 1 0 107548 0 -1 140352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_253_1165
timestamp 1
transform 1 0 108284 0 -1 140352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_254_3
timestamp 1636968456
transform 1 0 1380 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_15
timestamp 1636968456
transform 1 0 2484 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_254_27
timestamp 1
transform 1 0 3588 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_29
timestamp 1636968456
transform 1 0 3772 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_41
timestamp 1636968456
transform 1 0 4876 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_53
timestamp 1636968456
transform 1 0 5980 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_65
timestamp 1636968456
transform 1 0 7084 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_77
timestamp 1
transform 1 0 8188 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_83
timestamp 1
transform 1 0 8740 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_85
timestamp 1636968456
transform 1 0 8924 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_97
timestamp 1636968456
transform 1 0 10028 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_109
timestamp 1636968456
transform 1 0 11132 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_121
timestamp 1636968456
transform 1 0 12236 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_133
timestamp 1
transform 1 0 13340 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_139
timestamp 1
transform 1 0 13892 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_141
timestamp 1636968456
transform 1 0 14076 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_153
timestamp 1636968456
transform 1 0 15180 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_165
timestamp 1636968456
transform 1 0 16284 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_177
timestamp 1636968456
transform 1 0 17388 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_189
timestamp 1
transform 1 0 18492 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_195
timestamp 1
transform 1 0 19044 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_197
timestamp 1636968456
transform 1 0 19228 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_209
timestamp 1636968456
transform 1 0 20332 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_221
timestamp 1636968456
transform 1 0 21436 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_233
timestamp 1636968456
transform 1 0 22540 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_245
timestamp 1
transform 1 0 23644 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_251
timestamp 1
transform 1 0 24196 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_253
timestamp 1636968456
transform 1 0 24380 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_265
timestamp 1636968456
transform 1 0 25484 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_277
timestamp 1636968456
transform 1 0 26588 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_289
timestamp 1636968456
transform 1 0 27692 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_301
timestamp 1
transform 1 0 28796 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_307
timestamp 1
transform 1 0 29348 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_309
timestamp 1636968456
transform 1 0 29532 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_321
timestamp 1636968456
transform 1 0 30636 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_333
timestamp 1636968456
transform 1 0 31740 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_345
timestamp 1636968456
transform 1 0 32844 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_357
timestamp 1
transform 1 0 33948 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_363
timestamp 1
transform 1 0 34500 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_365
timestamp 1636968456
transform 1 0 34684 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_377
timestamp 1636968456
transform 1 0 35788 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_389
timestamp 1636968456
transform 1 0 36892 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_401
timestamp 1636968456
transform 1 0 37996 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_413
timestamp 1
transform 1 0 39100 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_419
timestamp 1
transform 1 0 39652 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_421
timestamp 1636968456
transform 1 0 39836 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_433
timestamp 1636968456
transform 1 0 40940 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_445
timestamp 1636968456
transform 1 0 42044 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_457
timestamp 1636968456
transform 1 0 43148 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_469
timestamp 1
transform 1 0 44252 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_475
timestamp 1
transform 1 0 44804 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_477
timestamp 1636968456
transform 1 0 44988 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_489
timestamp 1636968456
transform 1 0 46092 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_501
timestamp 1636968456
transform 1 0 47196 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_513
timestamp 1636968456
transform 1 0 48300 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_525
timestamp 1
transform 1 0 49404 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_531
timestamp 1
transform 1 0 49956 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_533
timestamp 1636968456
transform 1 0 50140 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_545
timestamp 1636968456
transform 1 0 51244 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_557
timestamp 1636968456
transform 1 0 52348 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_569
timestamp 1636968456
transform 1 0 53452 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_581
timestamp 1
transform 1 0 54556 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_587
timestamp 1
transform 1 0 55108 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_589
timestamp 1636968456
transform 1 0 55292 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_601
timestamp 1636968456
transform 1 0 56396 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_613
timestamp 1636968456
transform 1 0 57500 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_625
timestamp 1636968456
transform 1 0 58604 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_637
timestamp 1
transform 1 0 59708 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_643
timestamp 1
transform 1 0 60260 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_645
timestamp 1636968456
transform 1 0 60444 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_657
timestamp 1636968456
transform 1 0 61548 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_669
timestamp 1636968456
transform 1 0 62652 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_681
timestamp 1636968456
transform 1 0 63756 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_693
timestamp 1
transform 1 0 64860 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_699
timestamp 1
transform 1 0 65412 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_701
timestamp 1636968456
transform 1 0 65596 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_713
timestamp 1636968456
transform 1 0 66700 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_725
timestamp 1636968456
transform 1 0 67804 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_737
timestamp 1636968456
transform 1 0 68908 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_749
timestamp 1
transform 1 0 70012 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_755
timestamp 1
transform 1 0 70564 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_757
timestamp 1636968456
transform 1 0 70748 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_769
timestamp 1636968456
transform 1 0 71852 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_781
timestamp 1636968456
transform 1 0 72956 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_793
timestamp 1636968456
transform 1 0 74060 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_805
timestamp 1
transform 1 0 75164 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_811
timestamp 1
transform 1 0 75716 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_813
timestamp 1636968456
transform 1 0 75900 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_825
timestamp 1636968456
transform 1 0 77004 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_837
timestamp 1636968456
transform 1 0 78108 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_849
timestamp 1636968456
transform 1 0 79212 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_861
timestamp 1
transform 1 0 80316 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_867
timestamp 1
transform 1 0 80868 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_869
timestamp 1636968456
transform 1 0 81052 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_881
timestamp 1636968456
transform 1 0 82156 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_893
timestamp 1636968456
transform 1 0 83260 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_905
timestamp 1636968456
transform 1 0 84364 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_917
timestamp 1
transform 1 0 85468 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_923
timestamp 1
transform 1 0 86020 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_925
timestamp 1636968456
transform 1 0 86204 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_937
timestamp 1636968456
transform 1 0 87308 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_949
timestamp 1636968456
transform 1 0 88412 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_961
timestamp 1636968456
transform 1 0 89516 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_973
timestamp 1
transform 1 0 90620 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_979
timestamp 1
transform 1 0 91172 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_981
timestamp 1636968456
transform 1 0 91356 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_993
timestamp 1636968456
transform 1 0 92460 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1005
timestamp 1636968456
transform 1 0 93564 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1017
timestamp 1636968456
transform 1 0 94668 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_1029
timestamp 1
transform 1 0 95772 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_1035
timestamp 1
transform 1 0 96324 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1037
timestamp 1636968456
transform 1 0 96508 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1049
timestamp 1636968456
transform 1 0 97612 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1061
timestamp 1636968456
transform 1 0 98716 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1073
timestamp 1636968456
transform 1 0 99820 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_1085
timestamp 1
transform 1 0 100924 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_1091
timestamp 1
transform 1 0 101476 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1093
timestamp 1636968456
transform 1 0 101660 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1105
timestamp 1636968456
transform 1 0 102764 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1117
timestamp 1636968456
transform 1 0 103868 0 1 140352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1129
timestamp 1636968456
transform 1 0 104972 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_1141
timestamp 1
transform 1 0 106076 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_1147
timestamp 1
transform 1 0 106628 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_254_1149
timestamp 1636968456
transform 1 0 106812 0 1 140352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_254_1161
timestamp 1
transform 1 0 107916 0 1 140352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_254_1167
timestamp 1
transform 1 0 108468 0 1 140352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_3
timestamp 1636968456
transform 1 0 1380 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_15
timestamp 1636968456
transform 1 0 2484 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_27
timestamp 1636968456
transform 1 0 3588 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_39
timestamp 1636968456
transform 1 0 4692 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_255_51
timestamp 1
transform 1 0 5796 0 -1 141440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_255_55
timestamp 1
transform 1 0 6164 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_57
timestamp 1636968456
transform 1 0 6348 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_69
timestamp 1636968456
transform 1 0 7452 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_81
timestamp 1636968456
transform 1 0 8556 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_93
timestamp 1636968456
transform 1 0 9660 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_105
timestamp 1
transform 1 0 10764 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_111
timestamp 1
transform 1 0 11316 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_113
timestamp 1636968456
transform 1 0 11500 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_125
timestamp 1636968456
transform 1 0 12604 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_137
timestamp 1636968456
transform 1 0 13708 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_149
timestamp 1636968456
transform 1 0 14812 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_161
timestamp 1
transform 1 0 15916 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_167
timestamp 1
transform 1 0 16468 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_169
timestamp 1636968456
transform 1 0 16652 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_181
timestamp 1636968456
transform 1 0 17756 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_193
timestamp 1636968456
transform 1 0 18860 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_205
timestamp 1636968456
transform 1 0 19964 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_217
timestamp 1
transform 1 0 21068 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_223
timestamp 1
transform 1 0 21620 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_225
timestamp 1636968456
transform 1 0 21804 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_237
timestamp 1636968456
transform 1 0 22908 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_249
timestamp 1636968456
transform 1 0 24012 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_261
timestamp 1636968456
transform 1 0 25116 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_273
timestamp 1
transform 1 0 26220 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_279
timestamp 1
transform 1 0 26772 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_281
timestamp 1636968456
transform 1 0 26956 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_293
timestamp 1636968456
transform 1 0 28060 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_305
timestamp 1636968456
transform 1 0 29164 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_317
timestamp 1636968456
transform 1 0 30268 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_329
timestamp 1
transform 1 0 31372 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_335
timestamp 1
transform 1 0 31924 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_337
timestamp 1636968456
transform 1 0 32108 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_349
timestamp 1636968456
transform 1 0 33212 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_361
timestamp 1636968456
transform 1 0 34316 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_373
timestamp 1636968456
transform 1 0 35420 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_385
timestamp 1
transform 1 0 36524 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_391
timestamp 1
transform 1 0 37076 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_393
timestamp 1636968456
transform 1 0 37260 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_405
timestamp 1636968456
transform 1 0 38364 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_417
timestamp 1636968456
transform 1 0 39468 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_429
timestamp 1636968456
transform 1 0 40572 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_441
timestamp 1
transform 1 0 41676 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_447
timestamp 1
transform 1 0 42228 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_449
timestamp 1636968456
transform 1 0 42412 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_461
timestamp 1636968456
transform 1 0 43516 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_473
timestamp 1636968456
transform 1 0 44620 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_485
timestamp 1636968456
transform 1 0 45724 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_497
timestamp 1
transform 1 0 46828 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_503
timestamp 1
transform 1 0 47380 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_505
timestamp 1636968456
transform 1 0 47564 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_517
timestamp 1636968456
transform 1 0 48668 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_529
timestamp 1636968456
transform 1 0 49772 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_541
timestamp 1636968456
transform 1 0 50876 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_553
timestamp 1
transform 1 0 51980 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_559
timestamp 1
transform 1 0 52532 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_561
timestamp 1636968456
transform 1 0 52716 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_573
timestamp 1636968456
transform 1 0 53820 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_585
timestamp 1636968456
transform 1 0 54924 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_597
timestamp 1636968456
transform 1 0 56028 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_609
timestamp 1
transform 1 0 57132 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_615
timestamp 1
transform 1 0 57684 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_617
timestamp 1636968456
transform 1 0 57868 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_629
timestamp 1636968456
transform 1 0 58972 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_641
timestamp 1636968456
transform 1 0 60076 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_653
timestamp 1636968456
transform 1 0 61180 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_665
timestamp 1
transform 1 0 62284 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_671
timestamp 1
transform 1 0 62836 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_673
timestamp 1636968456
transform 1 0 63020 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_685
timestamp 1636968456
transform 1 0 64124 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_697
timestamp 1636968456
transform 1 0 65228 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_709
timestamp 1636968456
transform 1 0 66332 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_721
timestamp 1
transform 1 0 67436 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_727
timestamp 1
transform 1 0 67988 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_729
timestamp 1636968456
transform 1 0 68172 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_741
timestamp 1636968456
transform 1 0 69276 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_753
timestamp 1636968456
transform 1 0 70380 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_765
timestamp 1636968456
transform 1 0 71484 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_777
timestamp 1
transform 1 0 72588 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_783
timestamp 1
transform 1 0 73140 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_785
timestamp 1636968456
transform 1 0 73324 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_797
timestamp 1636968456
transform 1 0 74428 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_809
timestamp 1636968456
transform 1 0 75532 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_821
timestamp 1636968456
transform 1 0 76636 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_833
timestamp 1
transform 1 0 77740 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_839
timestamp 1
transform 1 0 78292 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_841
timestamp 1636968456
transform 1 0 78476 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_853
timestamp 1636968456
transform 1 0 79580 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_865
timestamp 1636968456
transform 1 0 80684 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_877
timestamp 1636968456
transform 1 0 81788 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_889
timestamp 1
transform 1 0 82892 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_895
timestamp 1
transform 1 0 83444 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_897
timestamp 1636968456
transform 1 0 83628 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_909
timestamp 1636968456
transform 1 0 84732 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_921
timestamp 1636968456
transform 1 0 85836 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_933
timestamp 1636968456
transform 1 0 86940 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_945
timestamp 1
transform 1 0 88044 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_951
timestamp 1
transform 1 0 88596 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_953
timestamp 1636968456
transform 1 0 88780 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_965
timestamp 1636968456
transform 1 0 89884 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_977
timestamp 1636968456
transform 1 0 90988 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_989
timestamp 1636968456
transform 1 0 92092 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_1001
timestamp 1
transform 1 0 93196 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_1007
timestamp 1
transform 1 0 93748 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1009
timestamp 1636968456
transform 1 0 93932 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1021
timestamp 1636968456
transform 1 0 95036 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1033
timestamp 1636968456
transform 1 0 96140 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1045
timestamp 1636968456
transform 1 0 97244 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_1057
timestamp 1
transform 1 0 98348 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_1063
timestamp 1
transform 1 0 98900 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1065
timestamp 1636968456
transform 1 0 99084 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1077
timestamp 1636968456
transform 1 0 100188 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1089
timestamp 1636968456
transform 1 0 101292 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1101
timestamp 1636968456
transform 1 0 102396 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_255_1113
timestamp 1
transform 1 0 103500 0 -1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_255_1119
timestamp 1
transform 1 0 104052 0 -1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1121
timestamp 1636968456
transform 1 0 104236 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1133
timestamp 1636968456
transform 1 0 105340 0 -1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_255_1145
timestamp 1636968456
transform 1 0 106444 0 -1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_255_1157
timestamp 1
transform 1 0 107548 0 -1 141440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_255_1165
timestamp 1
transform 1 0 108284 0 -1 141440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_256_3
timestamp 1636968456
transform 1 0 1380 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_15
timestamp 1636968456
transform 1 0 2484 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_256_27
timestamp 1
transform 1 0 3588 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_29
timestamp 1636968456
transform 1 0 3772 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_41
timestamp 1636968456
transform 1 0 4876 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_53
timestamp 1636968456
transform 1 0 5980 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_65
timestamp 1636968456
transform 1 0 7084 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_77
timestamp 1
transform 1 0 8188 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_83
timestamp 1
transform 1 0 8740 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_85
timestamp 1636968456
transform 1 0 8924 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_97
timestamp 1636968456
transform 1 0 10028 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_109
timestamp 1636968456
transform 1 0 11132 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_121
timestamp 1636968456
transform 1 0 12236 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_133
timestamp 1
transform 1 0 13340 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_139
timestamp 1
transform 1 0 13892 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_141
timestamp 1636968456
transform 1 0 14076 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_153
timestamp 1636968456
transform 1 0 15180 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_165
timestamp 1636968456
transform 1 0 16284 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_177
timestamp 1636968456
transform 1 0 17388 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_189
timestamp 1
transform 1 0 18492 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_195
timestamp 1
transform 1 0 19044 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_197
timestamp 1636968456
transform 1 0 19228 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_209
timestamp 1636968456
transform 1 0 20332 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_221
timestamp 1636968456
transform 1 0 21436 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_233
timestamp 1636968456
transform 1 0 22540 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_245
timestamp 1
transform 1 0 23644 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_251
timestamp 1
transform 1 0 24196 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_253
timestamp 1636968456
transform 1 0 24380 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_265
timestamp 1636968456
transform 1 0 25484 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_277
timestamp 1636968456
transform 1 0 26588 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_289
timestamp 1636968456
transform 1 0 27692 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_301
timestamp 1
transform 1 0 28796 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_307
timestamp 1
transform 1 0 29348 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_309
timestamp 1636968456
transform 1 0 29532 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_321
timestamp 1636968456
transform 1 0 30636 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_333
timestamp 1636968456
transform 1 0 31740 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_345
timestamp 1636968456
transform 1 0 32844 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_357
timestamp 1
transform 1 0 33948 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_363
timestamp 1
transform 1 0 34500 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_365
timestamp 1636968456
transform 1 0 34684 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_377
timestamp 1636968456
transform 1 0 35788 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_389
timestamp 1636968456
transform 1 0 36892 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_401
timestamp 1636968456
transform 1 0 37996 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_413
timestamp 1
transform 1 0 39100 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_419
timestamp 1
transform 1 0 39652 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_421
timestamp 1636968456
transform 1 0 39836 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_433
timestamp 1636968456
transform 1 0 40940 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_445
timestamp 1636968456
transform 1 0 42044 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_457
timestamp 1636968456
transform 1 0 43148 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_469
timestamp 1
transform 1 0 44252 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_475
timestamp 1
transform 1 0 44804 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_477
timestamp 1636968456
transform 1 0 44988 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_489
timestamp 1636968456
transform 1 0 46092 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_501
timestamp 1636968456
transform 1 0 47196 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_513
timestamp 1636968456
transform 1 0 48300 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_525
timestamp 1
transform 1 0 49404 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_531
timestamp 1
transform 1 0 49956 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_533
timestamp 1636968456
transform 1 0 50140 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_545
timestamp 1636968456
transform 1 0 51244 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_557
timestamp 1636968456
transform 1 0 52348 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_569
timestamp 1636968456
transform 1 0 53452 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_581
timestamp 1
transform 1 0 54556 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_587
timestamp 1
transform 1 0 55108 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_589
timestamp 1636968456
transform 1 0 55292 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_601
timestamp 1636968456
transform 1 0 56396 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_613
timestamp 1636968456
transform 1 0 57500 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_625
timestamp 1636968456
transform 1 0 58604 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_637
timestamp 1
transform 1 0 59708 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_643
timestamp 1
transform 1 0 60260 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_645
timestamp 1636968456
transform 1 0 60444 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_657
timestamp 1636968456
transform 1 0 61548 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_669
timestamp 1636968456
transform 1 0 62652 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_681
timestamp 1636968456
transform 1 0 63756 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_693
timestamp 1
transform 1 0 64860 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_699
timestamp 1
transform 1 0 65412 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_701
timestamp 1636968456
transform 1 0 65596 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_713
timestamp 1636968456
transform 1 0 66700 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_725
timestamp 1636968456
transform 1 0 67804 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_737
timestamp 1636968456
transform 1 0 68908 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_749
timestamp 1
transform 1 0 70012 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_755
timestamp 1
transform 1 0 70564 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_757
timestamp 1636968456
transform 1 0 70748 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_769
timestamp 1636968456
transform 1 0 71852 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_781
timestamp 1636968456
transform 1 0 72956 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_793
timestamp 1636968456
transform 1 0 74060 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_805
timestamp 1
transform 1 0 75164 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_811
timestamp 1
transform 1 0 75716 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_813
timestamp 1636968456
transform 1 0 75900 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_825
timestamp 1636968456
transform 1 0 77004 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_837
timestamp 1636968456
transform 1 0 78108 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_849
timestamp 1636968456
transform 1 0 79212 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_861
timestamp 1
transform 1 0 80316 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_867
timestamp 1
transform 1 0 80868 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_869
timestamp 1636968456
transform 1 0 81052 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_881
timestamp 1636968456
transform 1 0 82156 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_893
timestamp 1636968456
transform 1 0 83260 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_905
timestamp 1636968456
transform 1 0 84364 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_917
timestamp 1
transform 1 0 85468 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_923
timestamp 1
transform 1 0 86020 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_925
timestamp 1636968456
transform 1 0 86204 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_937
timestamp 1636968456
transform 1 0 87308 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_949
timestamp 1636968456
transform 1 0 88412 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_961
timestamp 1636968456
transform 1 0 89516 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_973
timestamp 1
transform 1 0 90620 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_979
timestamp 1
transform 1 0 91172 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_981
timestamp 1636968456
transform 1 0 91356 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_993
timestamp 1636968456
transform 1 0 92460 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1005
timestamp 1636968456
transform 1 0 93564 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1017
timestamp 1636968456
transform 1 0 94668 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_1029
timestamp 1
transform 1 0 95772 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_1035
timestamp 1
transform 1 0 96324 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1037
timestamp 1636968456
transform 1 0 96508 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1049
timestamp 1636968456
transform 1 0 97612 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1061
timestamp 1636968456
transform 1 0 98716 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1073
timestamp 1636968456
transform 1 0 99820 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_1085
timestamp 1
transform 1 0 100924 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_1091
timestamp 1
transform 1 0 101476 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1093
timestamp 1636968456
transform 1 0 101660 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1105
timestamp 1636968456
transform 1 0 102764 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1117
timestamp 1636968456
transform 1 0 103868 0 1 141440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1129
timestamp 1636968456
transform 1 0 104972 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_1141
timestamp 1
transform 1 0 106076 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_1147
timestamp 1
transform 1 0 106628 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_256_1149
timestamp 1636968456
transform 1 0 106812 0 1 141440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_256_1161
timestamp 1
transform 1 0 107916 0 1 141440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_256_1167
timestamp 1
transform 1 0 108468 0 1 141440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_3
timestamp 1636968456
transform 1 0 1380 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_15
timestamp 1636968456
transform 1 0 2484 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_27
timestamp 1636968456
transform 1 0 3588 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_39
timestamp 1636968456
transform 1 0 4692 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_257_51
timestamp 1
transform 1 0 5796 0 -1 142528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_257_55
timestamp 1
transform 1 0 6164 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_57
timestamp 1636968456
transform 1 0 6348 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_69
timestamp 1636968456
transform 1 0 7452 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_81
timestamp 1636968456
transform 1 0 8556 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_93
timestamp 1636968456
transform 1 0 9660 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_105
timestamp 1
transform 1 0 10764 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_111
timestamp 1
transform 1 0 11316 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_113
timestamp 1636968456
transform 1 0 11500 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_125
timestamp 1636968456
transform 1 0 12604 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_137
timestamp 1636968456
transform 1 0 13708 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_149
timestamp 1636968456
transform 1 0 14812 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_161
timestamp 1
transform 1 0 15916 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_167
timestamp 1
transform 1 0 16468 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_169
timestamp 1636968456
transform 1 0 16652 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_181
timestamp 1636968456
transform 1 0 17756 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_193
timestamp 1636968456
transform 1 0 18860 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_205
timestamp 1636968456
transform 1 0 19964 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_217
timestamp 1
transform 1 0 21068 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_223
timestamp 1
transform 1 0 21620 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_225
timestamp 1636968456
transform 1 0 21804 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_237
timestamp 1636968456
transform 1 0 22908 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_249
timestamp 1636968456
transform 1 0 24012 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_261
timestamp 1636968456
transform 1 0 25116 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_273
timestamp 1
transform 1 0 26220 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_279
timestamp 1
transform 1 0 26772 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_281
timestamp 1636968456
transform 1 0 26956 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_293
timestamp 1636968456
transform 1 0 28060 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_305
timestamp 1636968456
transform 1 0 29164 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_317
timestamp 1636968456
transform 1 0 30268 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_329
timestamp 1
transform 1 0 31372 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_335
timestamp 1
transform 1 0 31924 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_337
timestamp 1636968456
transform 1 0 32108 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_349
timestamp 1636968456
transform 1 0 33212 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_361
timestamp 1636968456
transform 1 0 34316 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_373
timestamp 1636968456
transform 1 0 35420 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_385
timestamp 1
transform 1 0 36524 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_391
timestamp 1
transform 1 0 37076 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_393
timestamp 1636968456
transform 1 0 37260 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_405
timestamp 1636968456
transform 1 0 38364 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_417
timestamp 1636968456
transform 1 0 39468 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_429
timestamp 1636968456
transform 1 0 40572 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_441
timestamp 1
transform 1 0 41676 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_447
timestamp 1
transform 1 0 42228 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_449
timestamp 1636968456
transform 1 0 42412 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_461
timestamp 1636968456
transform 1 0 43516 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_473
timestamp 1636968456
transform 1 0 44620 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_485
timestamp 1636968456
transform 1 0 45724 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_497
timestamp 1
transform 1 0 46828 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_503
timestamp 1
transform 1 0 47380 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_505
timestamp 1636968456
transform 1 0 47564 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_517
timestamp 1636968456
transform 1 0 48668 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_529
timestamp 1636968456
transform 1 0 49772 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_541
timestamp 1636968456
transform 1 0 50876 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_553
timestamp 1
transform 1 0 51980 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_559
timestamp 1
transform 1 0 52532 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_561
timestamp 1636968456
transform 1 0 52716 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_573
timestamp 1636968456
transform 1 0 53820 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_585
timestamp 1636968456
transform 1 0 54924 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_597
timestamp 1636968456
transform 1 0 56028 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_609
timestamp 1
transform 1 0 57132 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_615
timestamp 1
transform 1 0 57684 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_617
timestamp 1636968456
transform 1 0 57868 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_629
timestamp 1636968456
transform 1 0 58972 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_641
timestamp 1636968456
transform 1 0 60076 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_653
timestamp 1636968456
transform 1 0 61180 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_665
timestamp 1
transform 1 0 62284 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_671
timestamp 1
transform 1 0 62836 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_673
timestamp 1636968456
transform 1 0 63020 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_685
timestamp 1636968456
transform 1 0 64124 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_697
timestamp 1636968456
transform 1 0 65228 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_709
timestamp 1636968456
transform 1 0 66332 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_721
timestamp 1
transform 1 0 67436 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_727
timestamp 1
transform 1 0 67988 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_729
timestamp 1636968456
transform 1 0 68172 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_741
timestamp 1636968456
transform 1 0 69276 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_753
timestamp 1636968456
transform 1 0 70380 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_765
timestamp 1636968456
transform 1 0 71484 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_777
timestamp 1
transform 1 0 72588 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_783
timestamp 1
transform 1 0 73140 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_785
timestamp 1636968456
transform 1 0 73324 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_797
timestamp 1636968456
transform 1 0 74428 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_809
timestamp 1636968456
transform 1 0 75532 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_821
timestamp 1636968456
transform 1 0 76636 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_833
timestamp 1
transform 1 0 77740 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_839
timestamp 1
transform 1 0 78292 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_841
timestamp 1636968456
transform 1 0 78476 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_853
timestamp 1636968456
transform 1 0 79580 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_865
timestamp 1636968456
transform 1 0 80684 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_877
timestamp 1636968456
transform 1 0 81788 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_889
timestamp 1
transform 1 0 82892 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_895
timestamp 1
transform 1 0 83444 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_897
timestamp 1636968456
transform 1 0 83628 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_909
timestamp 1636968456
transform 1 0 84732 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_921
timestamp 1636968456
transform 1 0 85836 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_933
timestamp 1636968456
transform 1 0 86940 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_945
timestamp 1
transform 1 0 88044 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_951
timestamp 1
transform 1 0 88596 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_953
timestamp 1636968456
transform 1 0 88780 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_965
timestamp 1636968456
transform 1 0 89884 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_977
timestamp 1636968456
transform 1 0 90988 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_989
timestamp 1636968456
transform 1 0 92092 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_1001
timestamp 1
transform 1 0 93196 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_1007
timestamp 1
transform 1 0 93748 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1009
timestamp 1636968456
transform 1 0 93932 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1021
timestamp 1636968456
transform 1 0 95036 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1033
timestamp 1636968456
transform 1 0 96140 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1045
timestamp 1636968456
transform 1 0 97244 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_1057
timestamp 1
transform 1 0 98348 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_1063
timestamp 1
transform 1 0 98900 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1065
timestamp 1636968456
transform 1 0 99084 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1077
timestamp 1636968456
transform 1 0 100188 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1089
timestamp 1636968456
transform 1 0 101292 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1101
timestamp 1636968456
transform 1 0 102396 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_257_1113
timestamp 1
transform 1 0 103500 0 -1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_257_1119
timestamp 1
transform 1 0 104052 0 -1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1121
timestamp 1636968456
transform 1 0 104236 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1133
timestamp 1636968456
transform 1 0 105340 0 -1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_257_1145
timestamp 1636968456
transform 1 0 106444 0 -1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_257_1157
timestamp 1
transform 1 0 107548 0 -1 142528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_257_1165
timestamp 1
transform 1 0 108284 0 -1 142528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_258_3
timestamp 1636968456
transform 1 0 1380 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_15
timestamp 1636968456
transform 1 0 2484 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_258_27
timestamp 1
transform 1 0 3588 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_29
timestamp 1636968456
transform 1 0 3772 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_41
timestamp 1636968456
transform 1 0 4876 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_53
timestamp 1636968456
transform 1 0 5980 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_65
timestamp 1636968456
transform 1 0 7084 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_77
timestamp 1
transform 1 0 8188 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_83
timestamp 1
transform 1 0 8740 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_85
timestamp 1636968456
transform 1 0 8924 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_97
timestamp 1636968456
transform 1 0 10028 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_109
timestamp 1636968456
transform 1 0 11132 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_121
timestamp 1636968456
transform 1 0 12236 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_133
timestamp 1
transform 1 0 13340 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_139
timestamp 1
transform 1 0 13892 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_141
timestamp 1636968456
transform 1 0 14076 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_153
timestamp 1636968456
transform 1 0 15180 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_165
timestamp 1636968456
transform 1 0 16284 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_177
timestamp 1636968456
transform 1 0 17388 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_189
timestamp 1
transform 1 0 18492 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_195
timestamp 1
transform 1 0 19044 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_197
timestamp 1636968456
transform 1 0 19228 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_209
timestamp 1636968456
transform 1 0 20332 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_221
timestamp 1636968456
transform 1 0 21436 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_233
timestamp 1636968456
transform 1 0 22540 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_245
timestamp 1
transform 1 0 23644 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_251
timestamp 1
transform 1 0 24196 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_253
timestamp 1636968456
transform 1 0 24380 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_265
timestamp 1636968456
transform 1 0 25484 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_277
timestamp 1636968456
transform 1 0 26588 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_289
timestamp 1636968456
transform 1 0 27692 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_301
timestamp 1
transform 1 0 28796 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_307
timestamp 1
transform 1 0 29348 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_309
timestamp 1636968456
transform 1 0 29532 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_321
timestamp 1636968456
transform 1 0 30636 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_333
timestamp 1636968456
transform 1 0 31740 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_345
timestamp 1636968456
transform 1 0 32844 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_357
timestamp 1
transform 1 0 33948 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_363
timestamp 1
transform 1 0 34500 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_365
timestamp 1636968456
transform 1 0 34684 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_377
timestamp 1636968456
transform 1 0 35788 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_389
timestamp 1636968456
transform 1 0 36892 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_401
timestamp 1636968456
transform 1 0 37996 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_413
timestamp 1
transform 1 0 39100 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_419
timestamp 1
transform 1 0 39652 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_421
timestamp 1636968456
transform 1 0 39836 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_433
timestamp 1636968456
transform 1 0 40940 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_445
timestamp 1636968456
transform 1 0 42044 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_457
timestamp 1636968456
transform 1 0 43148 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_469
timestamp 1
transform 1 0 44252 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_475
timestamp 1
transform 1 0 44804 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_477
timestamp 1636968456
transform 1 0 44988 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_489
timestamp 1636968456
transform 1 0 46092 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_501
timestamp 1636968456
transform 1 0 47196 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_513
timestamp 1636968456
transform 1 0 48300 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_525
timestamp 1
transform 1 0 49404 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_531
timestamp 1
transform 1 0 49956 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_533
timestamp 1636968456
transform 1 0 50140 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_545
timestamp 1636968456
transform 1 0 51244 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_557
timestamp 1636968456
transform 1 0 52348 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_569
timestamp 1636968456
transform 1 0 53452 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_581
timestamp 1
transform 1 0 54556 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_587
timestamp 1
transform 1 0 55108 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_589
timestamp 1636968456
transform 1 0 55292 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_601
timestamp 1636968456
transform 1 0 56396 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_613
timestamp 1636968456
transform 1 0 57500 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_625
timestamp 1636968456
transform 1 0 58604 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_637
timestamp 1
transform 1 0 59708 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_643
timestamp 1
transform 1 0 60260 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_645
timestamp 1636968456
transform 1 0 60444 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_657
timestamp 1636968456
transform 1 0 61548 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_669
timestamp 1636968456
transform 1 0 62652 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_681
timestamp 1636968456
transform 1 0 63756 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_693
timestamp 1
transform 1 0 64860 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_699
timestamp 1
transform 1 0 65412 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_701
timestamp 1636968456
transform 1 0 65596 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_713
timestamp 1636968456
transform 1 0 66700 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_725
timestamp 1636968456
transform 1 0 67804 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_737
timestamp 1636968456
transform 1 0 68908 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_749
timestamp 1
transform 1 0 70012 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_755
timestamp 1
transform 1 0 70564 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_757
timestamp 1636968456
transform 1 0 70748 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_769
timestamp 1636968456
transform 1 0 71852 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_781
timestamp 1636968456
transform 1 0 72956 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_793
timestamp 1636968456
transform 1 0 74060 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_805
timestamp 1
transform 1 0 75164 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_811
timestamp 1
transform 1 0 75716 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_813
timestamp 1636968456
transform 1 0 75900 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_825
timestamp 1636968456
transform 1 0 77004 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_837
timestamp 1636968456
transform 1 0 78108 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_849
timestamp 1636968456
transform 1 0 79212 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_861
timestamp 1
transform 1 0 80316 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_867
timestamp 1
transform 1 0 80868 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_869
timestamp 1636968456
transform 1 0 81052 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_881
timestamp 1636968456
transform 1 0 82156 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_893
timestamp 1636968456
transform 1 0 83260 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_905
timestamp 1636968456
transform 1 0 84364 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_917
timestamp 1
transform 1 0 85468 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_923
timestamp 1
transform 1 0 86020 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_925
timestamp 1636968456
transform 1 0 86204 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_937
timestamp 1636968456
transform 1 0 87308 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_949
timestamp 1636968456
transform 1 0 88412 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_961
timestamp 1636968456
transform 1 0 89516 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_973
timestamp 1
transform 1 0 90620 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_979
timestamp 1
transform 1 0 91172 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_981
timestamp 1636968456
transform 1 0 91356 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_993
timestamp 1636968456
transform 1 0 92460 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1005
timestamp 1636968456
transform 1 0 93564 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1017
timestamp 1636968456
transform 1 0 94668 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_1029
timestamp 1
transform 1 0 95772 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_1035
timestamp 1
transform 1 0 96324 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1037
timestamp 1636968456
transform 1 0 96508 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1049
timestamp 1636968456
transform 1 0 97612 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1061
timestamp 1636968456
transform 1 0 98716 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1073
timestamp 1636968456
transform 1 0 99820 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_1085
timestamp 1
transform 1 0 100924 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_1091
timestamp 1
transform 1 0 101476 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1093
timestamp 1636968456
transform 1 0 101660 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1105
timestamp 1636968456
transform 1 0 102764 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1117
timestamp 1636968456
transform 1 0 103868 0 1 142528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1129
timestamp 1636968456
transform 1 0 104972 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_1141
timestamp 1
transform 1 0 106076 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_1147
timestamp 1
transform 1 0 106628 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_258_1149
timestamp 1636968456
transform 1 0 106812 0 1 142528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_258_1161
timestamp 1
transform 1 0 107916 0 1 142528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_258_1167
timestamp 1
transform 1 0 108468 0 1 142528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_3
timestamp 1636968456
transform 1 0 1380 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_15
timestamp 1636968456
transform 1 0 2484 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_27
timestamp 1636968456
transform 1 0 3588 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_39
timestamp 1636968456
transform 1 0 4692 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_259_51
timestamp 1
transform 1 0 5796 0 -1 143616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_259_55
timestamp 1
transform 1 0 6164 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_57
timestamp 1636968456
transform 1 0 6348 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_69
timestamp 1636968456
transform 1 0 7452 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_81
timestamp 1636968456
transform 1 0 8556 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_93
timestamp 1636968456
transform 1 0 9660 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_105
timestamp 1
transform 1 0 10764 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_111
timestamp 1
transform 1 0 11316 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_113
timestamp 1636968456
transform 1 0 11500 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_125
timestamp 1636968456
transform 1 0 12604 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_137
timestamp 1636968456
transform 1 0 13708 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_149
timestamp 1636968456
transform 1 0 14812 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_161
timestamp 1
transform 1 0 15916 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_167
timestamp 1
transform 1 0 16468 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_169
timestamp 1636968456
transform 1 0 16652 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_181
timestamp 1636968456
transform 1 0 17756 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_193
timestamp 1636968456
transform 1 0 18860 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_205
timestamp 1636968456
transform 1 0 19964 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_217
timestamp 1
transform 1 0 21068 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_223
timestamp 1
transform 1 0 21620 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_225
timestamp 1636968456
transform 1 0 21804 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_237
timestamp 1636968456
transform 1 0 22908 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_249
timestamp 1636968456
transform 1 0 24012 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_261
timestamp 1636968456
transform 1 0 25116 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_273
timestamp 1
transform 1 0 26220 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_279
timestamp 1
transform 1 0 26772 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_281
timestamp 1636968456
transform 1 0 26956 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_293
timestamp 1636968456
transform 1 0 28060 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_305
timestamp 1636968456
transform 1 0 29164 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_317
timestamp 1636968456
transform 1 0 30268 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_329
timestamp 1
transform 1 0 31372 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_335
timestamp 1
transform 1 0 31924 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_337
timestamp 1636968456
transform 1 0 32108 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_349
timestamp 1636968456
transform 1 0 33212 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_361
timestamp 1636968456
transform 1 0 34316 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_373
timestamp 1636968456
transform 1 0 35420 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_385
timestamp 1
transform 1 0 36524 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_391
timestamp 1
transform 1 0 37076 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_393
timestamp 1636968456
transform 1 0 37260 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_405
timestamp 1636968456
transform 1 0 38364 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_417
timestamp 1636968456
transform 1 0 39468 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_429
timestamp 1636968456
transform 1 0 40572 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_441
timestamp 1
transform 1 0 41676 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_447
timestamp 1
transform 1 0 42228 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_449
timestamp 1636968456
transform 1 0 42412 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_461
timestamp 1636968456
transform 1 0 43516 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_473
timestamp 1636968456
transform 1 0 44620 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_485
timestamp 1636968456
transform 1 0 45724 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_497
timestamp 1
transform 1 0 46828 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_503
timestamp 1
transform 1 0 47380 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_505
timestamp 1636968456
transform 1 0 47564 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_517
timestamp 1636968456
transform 1 0 48668 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_529
timestamp 1636968456
transform 1 0 49772 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_541
timestamp 1636968456
transform 1 0 50876 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_553
timestamp 1
transform 1 0 51980 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_559
timestamp 1
transform 1 0 52532 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_561
timestamp 1636968456
transform 1 0 52716 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_573
timestamp 1636968456
transform 1 0 53820 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_585
timestamp 1636968456
transform 1 0 54924 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_597
timestamp 1636968456
transform 1 0 56028 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_609
timestamp 1
transform 1 0 57132 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_615
timestamp 1
transform 1 0 57684 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_617
timestamp 1636968456
transform 1 0 57868 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_629
timestamp 1636968456
transform 1 0 58972 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_641
timestamp 1636968456
transform 1 0 60076 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_653
timestamp 1636968456
transform 1 0 61180 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_665
timestamp 1
transform 1 0 62284 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_671
timestamp 1
transform 1 0 62836 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_673
timestamp 1636968456
transform 1 0 63020 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_685
timestamp 1636968456
transform 1 0 64124 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_697
timestamp 1636968456
transform 1 0 65228 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_709
timestamp 1636968456
transform 1 0 66332 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_721
timestamp 1
transform 1 0 67436 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_727
timestamp 1
transform 1 0 67988 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_729
timestamp 1636968456
transform 1 0 68172 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_741
timestamp 1636968456
transform 1 0 69276 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_753
timestamp 1636968456
transform 1 0 70380 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_765
timestamp 1636968456
transform 1 0 71484 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_777
timestamp 1
transform 1 0 72588 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_783
timestamp 1
transform 1 0 73140 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_785
timestamp 1636968456
transform 1 0 73324 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_797
timestamp 1636968456
transform 1 0 74428 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_809
timestamp 1636968456
transform 1 0 75532 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_821
timestamp 1636968456
transform 1 0 76636 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_833
timestamp 1
transform 1 0 77740 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_839
timestamp 1
transform 1 0 78292 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_841
timestamp 1636968456
transform 1 0 78476 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_853
timestamp 1636968456
transform 1 0 79580 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_865
timestamp 1636968456
transform 1 0 80684 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_877
timestamp 1636968456
transform 1 0 81788 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_889
timestamp 1
transform 1 0 82892 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_895
timestamp 1
transform 1 0 83444 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_897
timestamp 1636968456
transform 1 0 83628 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_909
timestamp 1636968456
transform 1 0 84732 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_921
timestamp 1636968456
transform 1 0 85836 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_933
timestamp 1636968456
transform 1 0 86940 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_945
timestamp 1
transform 1 0 88044 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_951
timestamp 1
transform 1 0 88596 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_953
timestamp 1636968456
transform 1 0 88780 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_965
timestamp 1636968456
transform 1 0 89884 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_977
timestamp 1636968456
transform 1 0 90988 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_989
timestamp 1636968456
transform 1 0 92092 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_1001
timestamp 1
transform 1 0 93196 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_1007
timestamp 1
transform 1 0 93748 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1009
timestamp 1636968456
transform 1 0 93932 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1021
timestamp 1636968456
transform 1 0 95036 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1033
timestamp 1636968456
transform 1 0 96140 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1045
timestamp 1636968456
transform 1 0 97244 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_1057
timestamp 1
transform 1 0 98348 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_1063
timestamp 1
transform 1 0 98900 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1065
timestamp 1636968456
transform 1 0 99084 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1077
timestamp 1636968456
transform 1 0 100188 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1089
timestamp 1636968456
transform 1 0 101292 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1101
timestamp 1636968456
transform 1 0 102396 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_259_1113
timestamp 1
transform 1 0 103500 0 -1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_259_1119
timestamp 1
transform 1 0 104052 0 -1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1121
timestamp 1636968456
transform 1 0 104236 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1133
timestamp 1636968456
transform 1 0 105340 0 -1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_259_1145
timestamp 1636968456
transform 1 0 106444 0 -1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_259_1157
timestamp 1
transform 1 0 107548 0 -1 143616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_259_1165
timestamp 1
transform 1 0 108284 0 -1 143616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_260_3
timestamp 1636968456
transform 1 0 1380 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_15
timestamp 1636968456
transform 1 0 2484 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_260_27
timestamp 1
transform 1 0 3588 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_29
timestamp 1636968456
transform 1 0 3772 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_41
timestamp 1636968456
transform 1 0 4876 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_53
timestamp 1636968456
transform 1 0 5980 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_65
timestamp 1636968456
transform 1 0 7084 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_77
timestamp 1
transform 1 0 8188 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_83
timestamp 1
transform 1 0 8740 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_85
timestamp 1636968456
transform 1 0 8924 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_97
timestamp 1636968456
transform 1 0 10028 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_109
timestamp 1636968456
transform 1 0 11132 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_121
timestamp 1636968456
transform 1 0 12236 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_133
timestamp 1
transform 1 0 13340 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_139
timestamp 1
transform 1 0 13892 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_141
timestamp 1636968456
transform 1 0 14076 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_153
timestamp 1636968456
transform 1 0 15180 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_165
timestamp 1636968456
transform 1 0 16284 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_177
timestamp 1636968456
transform 1 0 17388 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_189
timestamp 1
transform 1 0 18492 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_195
timestamp 1
transform 1 0 19044 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_197
timestamp 1636968456
transform 1 0 19228 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_209
timestamp 1636968456
transform 1 0 20332 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_221
timestamp 1636968456
transform 1 0 21436 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_233
timestamp 1636968456
transform 1 0 22540 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_245
timestamp 1
transform 1 0 23644 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_251
timestamp 1
transform 1 0 24196 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_253
timestamp 1636968456
transform 1 0 24380 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_265
timestamp 1636968456
transform 1 0 25484 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_277
timestamp 1636968456
transform 1 0 26588 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_289
timestamp 1636968456
transform 1 0 27692 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_301
timestamp 1
transform 1 0 28796 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_307
timestamp 1
transform 1 0 29348 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_309
timestamp 1636968456
transform 1 0 29532 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_321
timestamp 1636968456
transform 1 0 30636 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_333
timestamp 1636968456
transform 1 0 31740 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_345
timestamp 1636968456
transform 1 0 32844 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_357
timestamp 1
transform 1 0 33948 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_363
timestamp 1
transform 1 0 34500 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_365
timestamp 1636968456
transform 1 0 34684 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_377
timestamp 1636968456
transform 1 0 35788 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_389
timestamp 1636968456
transform 1 0 36892 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_401
timestamp 1636968456
transform 1 0 37996 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_413
timestamp 1
transform 1 0 39100 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_419
timestamp 1
transform 1 0 39652 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_421
timestamp 1636968456
transform 1 0 39836 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_433
timestamp 1636968456
transform 1 0 40940 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_445
timestamp 1636968456
transform 1 0 42044 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_457
timestamp 1636968456
transform 1 0 43148 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_469
timestamp 1
transform 1 0 44252 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_475
timestamp 1
transform 1 0 44804 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_477
timestamp 1636968456
transform 1 0 44988 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_489
timestamp 1636968456
transform 1 0 46092 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_501
timestamp 1636968456
transform 1 0 47196 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_513
timestamp 1636968456
transform 1 0 48300 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_525
timestamp 1
transform 1 0 49404 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_531
timestamp 1
transform 1 0 49956 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_533
timestamp 1636968456
transform 1 0 50140 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_545
timestamp 1636968456
transform 1 0 51244 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_557
timestamp 1636968456
transform 1 0 52348 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_569
timestamp 1636968456
transform 1 0 53452 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_581
timestamp 1
transform 1 0 54556 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_587
timestamp 1
transform 1 0 55108 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_589
timestamp 1636968456
transform 1 0 55292 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_601
timestamp 1636968456
transform 1 0 56396 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_613
timestamp 1636968456
transform 1 0 57500 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_625
timestamp 1636968456
transform 1 0 58604 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_637
timestamp 1
transform 1 0 59708 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_643
timestamp 1
transform 1 0 60260 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_645
timestamp 1636968456
transform 1 0 60444 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_657
timestamp 1636968456
transform 1 0 61548 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_669
timestamp 1636968456
transform 1 0 62652 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_681
timestamp 1636968456
transform 1 0 63756 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_693
timestamp 1
transform 1 0 64860 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_699
timestamp 1
transform 1 0 65412 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_701
timestamp 1636968456
transform 1 0 65596 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_713
timestamp 1636968456
transform 1 0 66700 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_725
timestamp 1636968456
transform 1 0 67804 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_737
timestamp 1636968456
transform 1 0 68908 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_749
timestamp 1
transform 1 0 70012 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_755
timestamp 1
transform 1 0 70564 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_757
timestamp 1636968456
transform 1 0 70748 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_769
timestamp 1636968456
transform 1 0 71852 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_781
timestamp 1636968456
transform 1 0 72956 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_793
timestamp 1636968456
transform 1 0 74060 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_805
timestamp 1
transform 1 0 75164 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_811
timestamp 1
transform 1 0 75716 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_813
timestamp 1636968456
transform 1 0 75900 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_825
timestamp 1636968456
transform 1 0 77004 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_837
timestamp 1636968456
transform 1 0 78108 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_849
timestamp 1636968456
transform 1 0 79212 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_861
timestamp 1
transform 1 0 80316 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_867
timestamp 1
transform 1 0 80868 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_869
timestamp 1636968456
transform 1 0 81052 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_881
timestamp 1636968456
transform 1 0 82156 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_893
timestamp 1636968456
transform 1 0 83260 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_905
timestamp 1636968456
transform 1 0 84364 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_917
timestamp 1
transform 1 0 85468 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_923
timestamp 1
transform 1 0 86020 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_925
timestamp 1636968456
transform 1 0 86204 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_937
timestamp 1636968456
transform 1 0 87308 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_949
timestamp 1636968456
transform 1 0 88412 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_961
timestamp 1636968456
transform 1 0 89516 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_973
timestamp 1
transform 1 0 90620 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_979
timestamp 1
transform 1 0 91172 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_981
timestamp 1636968456
transform 1 0 91356 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_993
timestamp 1636968456
transform 1 0 92460 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1005
timestamp 1636968456
transform 1 0 93564 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1017
timestamp 1636968456
transform 1 0 94668 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_1029
timestamp 1
transform 1 0 95772 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_1035
timestamp 1
transform 1 0 96324 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1037
timestamp 1636968456
transform 1 0 96508 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1049
timestamp 1636968456
transform 1 0 97612 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1061
timestamp 1636968456
transform 1 0 98716 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1073
timestamp 1636968456
transform 1 0 99820 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_1085
timestamp 1
transform 1 0 100924 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_1091
timestamp 1
transform 1 0 101476 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1093
timestamp 1636968456
transform 1 0 101660 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1105
timestamp 1636968456
transform 1 0 102764 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1117
timestamp 1636968456
transform 1 0 103868 0 1 143616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1129
timestamp 1636968456
transform 1 0 104972 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_1141
timestamp 1
transform 1 0 106076 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_1147
timestamp 1
transform 1 0 106628 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_260_1149
timestamp 1636968456
transform 1 0 106812 0 1 143616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_260_1161
timestamp 1
transform 1 0 107916 0 1 143616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_260_1167
timestamp 1
transform 1 0 108468 0 1 143616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_3
timestamp 1636968456
transform 1 0 1380 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_15
timestamp 1636968456
transform 1 0 2484 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_27
timestamp 1636968456
transform 1 0 3588 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_39
timestamp 1636968456
transform 1 0 4692 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_261_51
timestamp 1
transform 1 0 5796 0 -1 144704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_261_55
timestamp 1
transform 1 0 6164 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_57
timestamp 1636968456
transform 1 0 6348 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_69
timestamp 1636968456
transform 1 0 7452 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_81
timestamp 1636968456
transform 1 0 8556 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_93
timestamp 1636968456
transform 1 0 9660 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_105
timestamp 1
transform 1 0 10764 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_111
timestamp 1
transform 1 0 11316 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_113
timestamp 1636968456
transform 1 0 11500 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_125
timestamp 1636968456
transform 1 0 12604 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_137
timestamp 1636968456
transform 1 0 13708 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_149
timestamp 1636968456
transform 1 0 14812 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_161
timestamp 1
transform 1 0 15916 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_167
timestamp 1
transform 1 0 16468 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_169
timestamp 1636968456
transform 1 0 16652 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_181
timestamp 1636968456
transform 1 0 17756 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_193
timestamp 1636968456
transform 1 0 18860 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_205
timestamp 1636968456
transform 1 0 19964 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_217
timestamp 1
transform 1 0 21068 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_223
timestamp 1
transform 1 0 21620 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_225
timestamp 1636968456
transform 1 0 21804 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_237
timestamp 1636968456
transform 1 0 22908 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_249
timestamp 1636968456
transform 1 0 24012 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_261
timestamp 1636968456
transform 1 0 25116 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_273
timestamp 1
transform 1 0 26220 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_279
timestamp 1
transform 1 0 26772 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_281
timestamp 1636968456
transform 1 0 26956 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_293
timestamp 1636968456
transform 1 0 28060 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_305
timestamp 1636968456
transform 1 0 29164 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_317
timestamp 1636968456
transform 1 0 30268 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_329
timestamp 1
transform 1 0 31372 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_335
timestamp 1
transform 1 0 31924 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_337
timestamp 1636968456
transform 1 0 32108 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_349
timestamp 1636968456
transform 1 0 33212 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_361
timestamp 1636968456
transform 1 0 34316 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_373
timestamp 1636968456
transform 1 0 35420 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_385
timestamp 1
transform 1 0 36524 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_391
timestamp 1
transform 1 0 37076 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_393
timestamp 1636968456
transform 1 0 37260 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_405
timestamp 1636968456
transform 1 0 38364 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_417
timestamp 1636968456
transform 1 0 39468 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_429
timestamp 1636968456
transform 1 0 40572 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_441
timestamp 1
transform 1 0 41676 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_447
timestamp 1
transform 1 0 42228 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_449
timestamp 1636968456
transform 1 0 42412 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_461
timestamp 1636968456
transform 1 0 43516 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_473
timestamp 1636968456
transform 1 0 44620 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_485
timestamp 1636968456
transform 1 0 45724 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_497
timestamp 1
transform 1 0 46828 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_503
timestamp 1
transform 1 0 47380 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_505
timestamp 1636968456
transform 1 0 47564 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_517
timestamp 1636968456
transform 1 0 48668 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_529
timestamp 1636968456
transform 1 0 49772 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_541
timestamp 1636968456
transform 1 0 50876 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_553
timestamp 1
transform 1 0 51980 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_559
timestamp 1
transform 1 0 52532 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_561
timestamp 1636968456
transform 1 0 52716 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_573
timestamp 1636968456
transform 1 0 53820 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_585
timestamp 1636968456
transform 1 0 54924 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_597
timestamp 1636968456
transform 1 0 56028 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_609
timestamp 1
transform 1 0 57132 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_615
timestamp 1
transform 1 0 57684 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_617
timestamp 1636968456
transform 1 0 57868 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_629
timestamp 1636968456
transform 1 0 58972 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_641
timestamp 1636968456
transform 1 0 60076 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_653
timestamp 1636968456
transform 1 0 61180 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_665
timestamp 1
transform 1 0 62284 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_671
timestamp 1
transform 1 0 62836 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_673
timestamp 1636968456
transform 1 0 63020 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_685
timestamp 1636968456
transform 1 0 64124 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_697
timestamp 1636968456
transform 1 0 65228 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_709
timestamp 1636968456
transform 1 0 66332 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_721
timestamp 1
transform 1 0 67436 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_727
timestamp 1
transform 1 0 67988 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_729
timestamp 1636968456
transform 1 0 68172 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_741
timestamp 1636968456
transform 1 0 69276 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_753
timestamp 1636968456
transform 1 0 70380 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_765
timestamp 1636968456
transform 1 0 71484 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_777
timestamp 1
transform 1 0 72588 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_783
timestamp 1
transform 1 0 73140 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_785
timestamp 1636968456
transform 1 0 73324 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_797
timestamp 1636968456
transform 1 0 74428 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_809
timestamp 1636968456
transform 1 0 75532 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_821
timestamp 1636968456
transform 1 0 76636 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_833
timestamp 1
transform 1 0 77740 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_839
timestamp 1
transform 1 0 78292 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_841
timestamp 1636968456
transform 1 0 78476 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_853
timestamp 1636968456
transform 1 0 79580 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_865
timestamp 1636968456
transform 1 0 80684 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_877
timestamp 1636968456
transform 1 0 81788 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_889
timestamp 1
transform 1 0 82892 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_895
timestamp 1
transform 1 0 83444 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_897
timestamp 1636968456
transform 1 0 83628 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_909
timestamp 1636968456
transform 1 0 84732 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_921
timestamp 1636968456
transform 1 0 85836 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_933
timestamp 1636968456
transform 1 0 86940 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_945
timestamp 1
transform 1 0 88044 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_951
timestamp 1
transform 1 0 88596 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_953
timestamp 1636968456
transform 1 0 88780 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_965
timestamp 1636968456
transform 1 0 89884 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_977
timestamp 1636968456
transform 1 0 90988 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_989
timestamp 1636968456
transform 1 0 92092 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_1001
timestamp 1
transform 1 0 93196 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_1007
timestamp 1
transform 1 0 93748 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1009
timestamp 1636968456
transform 1 0 93932 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1021
timestamp 1636968456
transform 1 0 95036 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1033
timestamp 1636968456
transform 1 0 96140 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1045
timestamp 1636968456
transform 1 0 97244 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_1057
timestamp 1
transform 1 0 98348 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_1063
timestamp 1
transform 1 0 98900 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1065
timestamp 1636968456
transform 1 0 99084 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1077
timestamp 1636968456
transform 1 0 100188 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1089
timestamp 1636968456
transform 1 0 101292 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1101
timestamp 1636968456
transform 1 0 102396 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_261_1113
timestamp 1
transform 1 0 103500 0 -1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_261_1119
timestamp 1
transform 1 0 104052 0 -1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1121
timestamp 1636968456
transform 1 0 104236 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1133
timestamp 1636968456
transform 1 0 105340 0 -1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_261_1145
timestamp 1636968456
transform 1 0 106444 0 -1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_261_1157
timestamp 1
transform 1 0 107548 0 -1 144704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_261_1165
timestamp 1
transform 1 0 108284 0 -1 144704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_262_3
timestamp 1636968456
transform 1 0 1380 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_15
timestamp 1636968456
transform 1 0 2484 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_262_27
timestamp 1
transform 1 0 3588 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_29
timestamp 1636968456
transform 1 0 3772 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_41
timestamp 1636968456
transform 1 0 4876 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_53
timestamp 1636968456
transform 1 0 5980 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_65
timestamp 1636968456
transform 1 0 7084 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_77
timestamp 1
transform 1 0 8188 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_83
timestamp 1
transform 1 0 8740 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_85
timestamp 1636968456
transform 1 0 8924 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_97
timestamp 1636968456
transform 1 0 10028 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_109
timestamp 1636968456
transform 1 0 11132 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_121
timestamp 1636968456
transform 1 0 12236 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_133
timestamp 1
transform 1 0 13340 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_139
timestamp 1
transform 1 0 13892 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_141
timestamp 1636968456
transform 1 0 14076 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_153
timestamp 1636968456
transform 1 0 15180 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_165
timestamp 1636968456
transform 1 0 16284 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_177
timestamp 1636968456
transform 1 0 17388 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_189
timestamp 1
transform 1 0 18492 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_195
timestamp 1
transform 1 0 19044 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_197
timestamp 1636968456
transform 1 0 19228 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_209
timestamp 1636968456
transform 1 0 20332 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_221
timestamp 1636968456
transform 1 0 21436 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_233
timestamp 1636968456
transform 1 0 22540 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_245
timestamp 1
transform 1 0 23644 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_251
timestamp 1
transform 1 0 24196 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_253
timestamp 1636968456
transform 1 0 24380 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_265
timestamp 1636968456
transform 1 0 25484 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_277
timestamp 1636968456
transform 1 0 26588 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_289
timestamp 1636968456
transform 1 0 27692 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_301
timestamp 1
transform 1 0 28796 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_307
timestamp 1
transform 1 0 29348 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_309
timestamp 1636968456
transform 1 0 29532 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_321
timestamp 1636968456
transform 1 0 30636 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_333
timestamp 1636968456
transform 1 0 31740 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_345
timestamp 1636968456
transform 1 0 32844 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_357
timestamp 1
transform 1 0 33948 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_363
timestamp 1
transform 1 0 34500 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_365
timestamp 1636968456
transform 1 0 34684 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_377
timestamp 1636968456
transform 1 0 35788 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_389
timestamp 1636968456
transform 1 0 36892 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_401
timestamp 1636968456
transform 1 0 37996 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_413
timestamp 1
transform 1 0 39100 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_419
timestamp 1
transform 1 0 39652 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_421
timestamp 1636968456
transform 1 0 39836 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_433
timestamp 1636968456
transform 1 0 40940 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_445
timestamp 1636968456
transform 1 0 42044 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_457
timestamp 1636968456
transform 1 0 43148 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_469
timestamp 1
transform 1 0 44252 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_475
timestamp 1
transform 1 0 44804 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_477
timestamp 1636968456
transform 1 0 44988 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_489
timestamp 1636968456
transform 1 0 46092 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_501
timestamp 1636968456
transform 1 0 47196 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_513
timestamp 1636968456
transform 1 0 48300 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_525
timestamp 1
transform 1 0 49404 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_531
timestamp 1
transform 1 0 49956 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_533
timestamp 1636968456
transform 1 0 50140 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_545
timestamp 1636968456
transform 1 0 51244 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_557
timestamp 1636968456
transform 1 0 52348 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_569
timestamp 1636968456
transform 1 0 53452 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_581
timestamp 1
transform 1 0 54556 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_587
timestamp 1
transform 1 0 55108 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_589
timestamp 1636968456
transform 1 0 55292 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_601
timestamp 1636968456
transform 1 0 56396 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_613
timestamp 1636968456
transform 1 0 57500 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_625
timestamp 1636968456
transform 1 0 58604 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_637
timestamp 1
transform 1 0 59708 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_643
timestamp 1
transform 1 0 60260 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_645
timestamp 1636968456
transform 1 0 60444 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_657
timestamp 1636968456
transform 1 0 61548 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_669
timestamp 1636968456
transform 1 0 62652 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_681
timestamp 1636968456
transform 1 0 63756 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_693
timestamp 1
transform 1 0 64860 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_699
timestamp 1
transform 1 0 65412 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_701
timestamp 1636968456
transform 1 0 65596 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_713
timestamp 1636968456
transform 1 0 66700 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_725
timestamp 1636968456
transform 1 0 67804 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_737
timestamp 1636968456
transform 1 0 68908 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_749
timestamp 1
transform 1 0 70012 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_755
timestamp 1
transform 1 0 70564 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_757
timestamp 1636968456
transform 1 0 70748 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_769
timestamp 1636968456
transform 1 0 71852 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_781
timestamp 1636968456
transform 1 0 72956 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_793
timestamp 1636968456
transform 1 0 74060 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_805
timestamp 1
transform 1 0 75164 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_811
timestamp 1
transform 1 0 75716 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_813
timestamp 1636968456
transform 1 0 75900 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_825
timestamp 1636968456
transform 1 0 77004 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_837
timestamp 1636968456
transform 1 0 78108 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_849
timestamp 1636968456
transform 1 0 79212 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_861
timestamp 1
transform 1 0 80316 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_867
timestamp 1
transform 1 0 80868 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_869
timestamp 1636968456
transform 1 0 81052 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_881
timestamp 1636968456
transform 1 0 82156 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_893
timestamp 1636968456
transform 1 0 83260 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_905
timestamp 1636968456
transform 1 0 84364 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_917
timestamp 1
transform 1 0 85468 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_923
timestamp 1
transform 1 0 86020 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_925
timestamp 1636968456
transform 1 0 86204 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_937
timestamp 1636968456
transform 1 0 87308 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_949
timestamp 1636968456
transform 1 0 88412 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_961
timestamp 1636968456
transform 1 0 89516 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_973
timestamp 1
transform 1 0 90620 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_979
timestamp 1
transform 1 0 91172 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_981
timestamp 1636968456
transform 1 0 91356 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_993
timestamp 1636968456
transform 1 0 92460 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1005
timestamp 1636968456
transform 1 0 93564 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1017
timestamp 1636968456
transform 1 0 94668 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_1029
timestamp 1
transform 1 0 95772 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_1035
timestamp 1
transform 1 0 96324 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1037
timestamp 1636968456
transform 1 0 96508 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1049
timestamp 1636968456
transform 1 0 97612 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1061
timestamp 1636968456
transform 1 0 98716 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1073
timestamp 1636968456
transform 1 0 99820 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_1085
timestamp 1
transform 1 0 100924 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_1091
timestamp 1
transform 1 0 101476 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1093
timestamp 1636968456
transform 1 0 101660 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1105
timestamp 1636968456
transform 1 0 102764 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1117
timestamp 1636968456
transform 1 0 103868 0 1 144704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1129
timestamp 1636968456
transform 1 0 104972 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_1141
timestamp 1
transform 1 0 106076 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_1147
timestamp 1
transform 1 0 106628 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_262_1149
timestamp 1636968456
transform 1 0 106812 0 1 144704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_262_1161
timestamp 1
transform 1 0 107916 0 1 144704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_262_1167
timestamp 1
transform 1 0 108468 0 1 144704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_3
timestamp 1636968456
transform 1 0 1380 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_15
timestamp 1636968456
transform 1 0 2484 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_27
timestamp 1636968456
transform 1 0 3588 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_39
timestamp 1636968456
transform 1 0 4692 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_263_51
timestamp 1
transform 1 0 5796 0 -1 145792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_263_55
timestamp 1
transform 1 0 6164 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_57
timestamp 1636968456
transform 1 0 6348 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_69
timestamp 1636968456
transform 1 0 7452 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_81
timestamp 1636968456
transform 1 0 8556 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_93
timestamp 1636968456
transform 1 0 9660 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_105
timestamp 1
transform 1 0 10764 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_111
timestamp 1
transform 1 0 11316 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_113
timestamp 1636968456
transform 1 0 11500 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_125
timestamp 1636968456
transform 1 0 12604 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_137
timestamp 1636968456
transform 1 0 13708 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_149
timestamp 1636968456
transform 1 0 14812 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_161
timestamp 1
transform 1 0 15916 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_167
timestamp 1
transform 1 0 16468 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_169
timestamp 1636968456
transform 1 0 16652 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_181
timestamp 1636968456
transform 1 0 17756 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_193
timestamp 1636968456
transform 1 0 18860 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_205
timestamp 1636968456
transform 1 0 19964 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_217
timestamp 1
transform 1 0 21068 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_223
timestamp 1
transform 1 0 21620 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_225
timestamp 1636968456
transform 1 0 21804 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_237
timestamp 1636968456
transform 1 0 22908 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_249
timestamp 1636968456
transform 1 0 24012 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_261
timestamp 1636968456
transform 1 0 25116 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_273
timestamp 1
transform 1 0 26220 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_279
timestamp 1
transform 1 0 26772 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_281
timestamp 1636968456
transform 1 0 26956 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_293
timestamp 1636968456
transform 1 0 28060 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_305
timestamp 1636968456
transform 1 0 29164 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_317
timestamp 1636968456
transform 1 0 30268 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_329
timestamp 1
transform 1 0 31372 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_335
timestamp 1
transform 1 0 31924 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_337
timestamp 1636968456
transform 1 0 32108 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_349
timestamp 1636968456
transform 1 0 33212 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_361
timestamp 1636968456
transform 1 0 34316 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_373
timestamp 1636968456
transform 1 0 35420 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_385
timestamp 1
transform 1 0 36524 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_391
timestamp 1
transform 1 0 37076 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_393
timestamp 1636968456
transform 1 0 37260 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_405
timestamp 1636968456
transform 1 0 38364 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_417
timestamp 1636968456
transform 1 0 39468 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_429
timestamp 1636968456
transform 1 0 40572 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_441
timestamp 1
transform 1 0 41676 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_447
timestamp 1
transform 1 0 42228 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_449
timestamp 1636968456
transform 1 0 42412 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_461
timestamp 1636968456
transform 1 0 43516 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_473
timestamp 1636968456
transform 1 0 44620 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_485
timestamp 1636968456
transform 1 0 45724 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_497
timestamp 1
transform 1 0 46828 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_503
timestamp 1
transform 1 0 47380 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_505
timestamp 1636968456
transform 1 0 47564 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_517
timestamp 1636968456
transform 1 0 48668 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_529
timestamp 1636968456
transform 1 0 49772 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_541
timestamp 1636968456
transform 1 0 50876 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_553
timestamp 1
transform 1 0 51980 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_559
timestamp 1
transform 1 0 52532 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_561
timestamp 1636968456
transform 1 0 52716 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_573
timestamp 1636968456
transform 1 0 53820 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_585
timestamp 1636968456
transform 1 0 54924 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_597
timestamp 1636968456
transform 1 0 56028 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_609
timestamp 1
transform 1 0 57132 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_615
timestamp 1
transform 1 0 57684 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_617
timestamp 1636968456
transform 1 0 57868 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_629
timestamp 1636968456
transform 1 0 58972 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_641
timestamp 1636968456
transform 1 0 60076 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_653
timestamp 1636968456
transform 1 0 61180 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_665
timestamp 1
transform 1 0 62284 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_671
timestamp 1
transform 1 0 62836 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_673
timestamp 1636968456
transform 1 0 63020 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_685
timestamp 1636968456
transform 1 0 64124 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_697
timestamp 1636968456
transform 1 0 65228 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_709
timestamp 1636968456
transform 1 0 66332 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_721
timestamp 1
transform 1 0 67436 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_727
timestamp 1
transform 1 0 67988 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_729
timestamp 1636968456
transform 1 0 68172 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_741
timestamp 1636968456
transform 1 0 69276 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_753
timestamp 1636968456
transform 1 0 70380 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_765
timestamp 1636968456
transform 1 0 71484 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_777
timestamp 1
transform 1 0 72588 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_783
timestamp 1
transform 1 0 73140 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_785
timestamp 1636968456
transform 1 0 73324 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_797
timestamp 1636968456
transform 1 0 74428 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_809
timestamp 1636968456
transform 1 0 75532 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_821
timestamp 1636968456
transform 1 0 76636 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_833
timestamp 1
transform 1 0 77740 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_839
timestamp 1
transform 1 0 78292 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_841
timestamp 1636968456
transform 1 0 78476 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_853
timestamp 1636968456
transform 1 0 79580 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_865
timestamp 1636968456
transform 1 0 80684 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_877
timestamp 1636968456
transform 1 0 81788 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_889
timestamp 1
transform 1 0 82892 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_895
timestamp 1
transform 1 0 83444 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_897
timestamp 1636968456
transform 1 0 83628 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_909
timestamp 1636968456
transform 1 0 84732 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_921
timestamp 1636968456
transform 1 0 85836 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_933
timestamp 1636968456
transform 1 0 86940 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_945
timestamp 1
transform 1 0 88044 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_951
timestamp 1
transform 1 0 88596 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_953
timestamp 1636968456
transform 1 0 88780 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_965
timestamp 1636968456
transform 1 0 89884 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_977
timestamp 1636968456
transform 1 0 90988 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_989
timestamp 1636968456
transform 1 0 92092 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_1001
timestamp 1
transform 1 0 93196 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_1007
timestamp 1
transform 1 0 93748 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1009
timestamp 1636968456
transform 1 0 93932 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1021
timestamp 1636968456
transform 1 0 95036 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1033
timestamp 1636968456
transform 1 0 96140 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1045
timestamp 1636968456
transform 1 0 97244 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_1057
timestamp 1
transform 1 0 98348 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_1063
timestamp 1
transform 1 0 98900 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1065
timestamp 1636968456
transform 1 0 99084 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1077
timestamp 1636968456
transform 1 0 100188 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1089
timestamp 1636968456
transform 1 0 101292 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1101
timestamp 1636968456
transform 1 0 102396 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_263_1113
timestamp 1
transform 1 0 103500 0 -1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_263_1119
timestamp 1
transform 1 0 104052 0 -1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1121
timestamp 1636968456
transform 1 0 104236 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1133
timestamp 1636968456
transform 1 0 105340 0 -1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_263_1145
timestamp 1636968456
transform 1 0 106444 0 -1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_263_1157
timestamp 1
transform 1 0 107548 0 -1 145792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_263_1165
timestamp 1
transform 1 0 108284 0 -1 145792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_264_3
timestamp 1636968456
transform 1 0 1380 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_15
timestamp 1636968456
transform 1 0 2484 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_264_27
timestamp 1
transform 1 0 3588 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_29
timestamp 1636968456
transform 1 0 3772 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_41
timestamp 1636968456
transform 1 0 4876 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_53
timestamp 1636968456
transform 1 0 5980 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_65
timestamp 1636968456
transform 1 0 7084 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_77
timestamp 1
transform 1 0 8188 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_83
timestamp 1
transform 1 0 8740 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_85
timestamp 1636968456
transform 1 0 8924 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_97
timestamp 1636968456
transform 1 0 10028 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_109
timestamp 1636968456
transform 1 0 11132 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_121
timestamp 1636968456
transform 1 0 12236 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_133
timestamp 1
transform 1 0 13340 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_139
timestamp 1
transform 1 0 13892 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_141
timestamp 1636968456
transform 1 0 14076 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_153
timestamp 1636968456
transform 1 0 15180 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_165
timestamp 1636968456
transform 1 0 16284 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_177
timestamp 1636968456
transform 1 0 17388 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_189
timestamp 1
transform 1 0 18492 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_195
timestamp 1
transform 1 0 19044 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_197
timestamp 1636968456
transform 1 0 19228 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_209
timestamp 1636968456
transform 1 0 20332 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_221
timestamp 1636968456
transform 1 0 21436 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_233
timestamp 1636968456
transform 1 0 22540 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_245
timestamp 1
transform 1 0 23644 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_251
timestamp 1
transform 1 0 24196 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_253
timestamp 1636968456
transform 1 0 24380 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_265
timestamp 1636968456
transform 1 0 25484 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_277
timestamp 1636968456
transform 1 0 26588 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_289
timestamp 1636968456
transform 1 0 27692 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_301
timestamp 1
transform 1 0 28796 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_307
timestamp 1
transform 1 0 29348 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_309
timestamp 1636968456
transform 1 0 29532 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_321
timestamp 1636968456
transform 1 0 30636 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_333
timestamp 1636968456
transform 1 0 31740 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_345
timestamp 1636968456
transform 1 0 32844 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_357
timestamp 1
transform 1 0 33948 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_363
timestamp 1
transform 1 0 34500 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_365
timestamp 1636968456
transform 1 0 34684 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_377
timestamp 1636968456
transform 1 0 35788 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_389
timestamp 1636968456
transform 1 0 36892 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_401
timestamp 1636968456
transform 1 0 37996 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_413
timestamp 1
transform 1 0 39100 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_419
timestamp 1
transform 1 0 39652 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_421
timestamp 1636968456
transform 1 0 39836 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_433
timestamp 1636968456
transform 1 0 40940 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_445
timestamp 1636968456
transform 1 0 42044 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_457
timestamp 1636968456
transform 1 0 43148 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_469
timestamp 1
transform 1 0 44252 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_475
timestamp 1
transform 1 0 44804 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_477
timestamp 1636968456
transform 1 0 44988 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_489
timestamp 1636968456
transform 1 0 46092 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_501
timestamp 1636968456
transform 1 0 47196 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_513
timestamp 1636968456
transform 1 0 48300 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_525
timestamp 1
transform 1 0 49404 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_531
timestamp 1
transform 1 0 49956 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_533
timestamp 1636968456
transform 1 0 50140 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_545
timestamp 1636968456
transform 1 0 51244 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_557
timestamp 1636968456
transform 1 0 52348 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_569
timestamp 1636968456
transform 1 0 53452 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_581
timestamp 1
transform 1 0 54556 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_587
timestamp 1
transform 1 0 55108 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_589
timestamp 1636968456
transform 1 0 55292 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_601
timestamp 1636968456
transform 1 0 56396 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_613
timestamp 1636968456
transform 1 0 57500 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_625
timestamp 1636968456
transform 1 0 58604 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_637
timestamp 1
transform 1 0 59708 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_643
timestamp 1
transform 1 0 60260 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_645
timestamp 1636968456
transform 1 0 60444 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_657
timestamp 1636968456
transform 1 0 61548 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_669
timestamp 1636968456
transform 1 0 62652 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_681
timestamp 1636968456
transform 1 0 63756 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_693
timestamp 1
transform 1 0 64860 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_699
timestamp 1
transform 1 0 65412 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_701
timestamp 1636968456
transform 1 0 65596 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_713
timestamp 1636968456
transform 1 0 66700 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_725
timestamp 1636968456
transform 1 0 67804 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_737
timestamp 1636968456
transform 1 0 68908 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_749
timestamp 1
transform 1 0 70012 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_755
timestamp 1
transform 1 0 70564 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_757
timestamp 1636968456
transform 1 0 70748 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_769
timestamp 1636968456
transform 1 0 71852 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_781
timestamp 1636968456
transform 1 0 72956 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_793
timestamp 1636968456
transform 1 0 74060 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_805
timestamp 1
transform 1 0 75164 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_811
timestamp 1
transform 1 0 75716 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_813
timestamp 1636968456
transform 1 0 75900 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_825
timestamp 1636968456
transform 1 0 77004 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_837
timestamp 1636968456
transform 1 0 78108 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_849
timestamp 1636968456
transform 1 0 79212 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_861
timestamp 1
transform 1 0 80316 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_867
timestamp 1
transform 1 0 80868 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_869
timestamp 1636968456
transform 1 0 81052 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_881
timestamp 1636968456
transform 1 0 82156 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_893
timestamp 1636968456
transform 1 0 83260 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_905
timestamp 1636968456
transform 1 0 84364 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_917
timestamp 1
transform 1 0 85468 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_923
timestamp 1
transform 1 0 86020 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_925
timestamp 1636968456
transform 1 0 86204 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_937
timestamp 1636968456
transform 1 0 87308 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_949
timestamp 1636968456
transform 1 0 88412 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_961
timestamp 1636968456
transform 1 0 89516 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_973
timestamp 1
transform 1 0 90620 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_979
timestamp 1
transform 1 0 91172 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_981
timestamp 1636968456
transform 1 0 91356 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_993
timestamp 1636968456
transform 1 0 92460 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1005
timestamp 1636968456
transform 1 0 93564 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1017
timestamp 1636968456
transform 1 0 94668 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_1029
timestamp 1
transform 1 0 95772 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_1035
timestamp 1
transform 1 0 96324 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1037
timestamp 1636968456
transform 1 0 96508 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1049
timestamp 1636968456
transform 1 0 97612 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1061
timestamp 1636968456
transform 1 0 98716 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1073
timestamp 1636968456
transform 1 0 99820 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_1085
timestamp 1
transform 1 0 100924 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_1091
timestamp 1
transform 1 0 101476 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1093
timestamp 1636968456
transform 1 0 101660 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1105
timestamp 1636968456
transform 1 0 102764 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1117
timestamp 1636968456
transform 1 0 103868 0 1 145792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1129
timestamp 1636968456
transform 1 0 104972 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_1141
timestamp 1
transform 1 0 106076 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_1147
timestamp 1
transform 1 0 106628 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_264_1149
timestamp 1636968456
transform 1 0 106812 0 1 145792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_264_1161
timestamp 1
transform 1 0 107916 0 1 145792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_264_1167
timestamp 1
transform 1 0 108468 0 1 145792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_3
timestamp 1636968456
transform 1 0 1380 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_15
timestamp 1636968456
transform 1 0 2484 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_27
timestamp 1636968456
transform 1 0 3588 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_39
timestamp 1636968456
transform 1 0 4692 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_265_51
timestamp 1
transform 1 0 5796 0 -1 146880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_265_55
timestamp 1
transform 1 0 6164 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_57
timestamp 1636968456
transform 1 0 6348 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_69
timestamp 1636968456
transform 1 0 7452 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_81
timestamp 1636968456
transform 1 0 8556 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_93
timestamp 1636968456
transform 1 0 9660 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_105
timestamp 1
transform 1 0 10764 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_111
timestamp 1
transform 1 0 11316 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_113
timestamp 1636968456
transform 1 0 11500 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_125
timestamp 1636968456
transform 1 0 12604 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_137
timestamp 1636968456
transform 1 0 13708 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_149
timestamp 1636968456
transform 1 0 14812 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_161
timestamp 1
transform 1 0 15916 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_167
timestamp 1
transform 1 0 16468 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_169
timestamp 1636968456
transform 1 0 16652 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_181
timestamp 1636968456
transform 1 0 17756 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_193
timestamp 1636968456
transform 1 0 18860 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_205
timestamp 1636968456
transform 1 0 19964 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_217
timestamp 1
transform 1 0 21068 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_223
timestamp 1
transform 1 0 21620 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_225
timestamp 1636968456
transform 1 0 21804 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_237
timestamp 1636968456
transform 1 0 22908 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_249
timestamp 1636968456
transform 1 0 24012 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_261
timestamp 1636968456
transform 1 0 25116 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_273
timestamp 1
transform 1 0 26220 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_279
timestamp 1
transform 1 0 26772 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_281
timestamp 1636968456
transform 1 0 26956 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_293
timestamp 1636968456
transform 1 0 28060 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_305
timestamp 1636968456
transform 1 0 29164 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_317
timestamp 1636968456
transform 1 0 30268 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_329
timestamp 1
transform 1 0 31372 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_335
timestamp 1
transform 1 0 31924 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_337
timestamp 1636968456
transform 1 0 32108 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_349
timestamp 1636968456
transform 1 0 33212 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_361
timestamp 1636968456
transform 1 0 34316 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_373
timestamp 1636968456
transform 1 0 35420 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_385
timestamp 1
transform 1 0 36524 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_391
timestamp 1
transform 1 0 37076 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_393
timestamp 1636968456
transform 1 0 37260 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_405
timestamp 1636968456
transform 1 0 38364 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_417
timestamp 1636968456
transform 1 0 39468 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_429
timestamp 1636968456
transform 1 0 40572 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_441
timestamp 1
transform 1 0 41676 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_447
timestamp 1
transform 1 0 42228 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_449
timestamp 1636968456
transform 1 0 42412 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_461
timestamp 1636968456
transform 1 0 43516 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_473
timestamp 1636968456
transform 1 0 44620 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_485
timestamp 1636968456
transform 1 0 45724 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_497
timestamp 1
transform 1 0 46828 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_503
timestamp 1
transform 1 0 47380 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_505
timestamp 1636968456
transform 1 0 47564 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_517
timestamp 1636968456
transform 1 0 48668 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_529
timestamp 1636968456
transform 1 0 49772 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_541
timestamp 1636968456
transform 1 0 50876 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_553
timestamp 1
transform 1 0 51980 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_559
timestamp 1
transform 1 0 52532 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_561
timestamp 1636968456
transform 1 0 52716 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_573
timestamp 1636968456
transform 1 0 53820 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_585
timestamp 1636968456
transform 1 0 54924 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_597
timestamp 1636968456
transform 1 0 56028 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_609
timestamp 1
transform 1 0 57132 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_615
timestamp 1
transform 1 0 57684 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_617
timestamp 1636968456
transform 1 0 57868 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_629
timestamp 1636968456
transform 1 0 58972 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_641
timestamp 1636968456
transform 1 0 60076 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_653
timestamp 1636968456
transform 1 0 61180 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_665
timestamp 1
transform 1 0 62284 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_671
timestamp 1
transform 1 0 62836 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_673
timestamp 1636968456
transform 1 0 63020 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_685
timestamp 1636968456
transform 1 0 64124 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_697
timestamp 1636968456
transform 1 0 65228 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_709
timestamp 1636968456
transform 1 0 66332 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_721
timestamp 1
transform 1 0 67436 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_727
timestamp 1
transform 1 0 67988 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_729
timestamp 1636968456
transform 1 0 68172 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_741
timestamp 1636968456
transform 1 0 69276 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_753
timestamp 1636968456
transform 1 0 70380 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_765
timestamp 1636968456
transform 1 0 71484 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_777
timestamp 1
transform 1 0 72588 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_783
timestamp 1
transform 1 0 73140 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_785
timestamp 1636968456
transform 1 0 73324 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_797
timestamp 1636968456
transform 1 0 74428 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_809
timestamp 1636968456
transform 1 0 75532 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_821
timestamp 1636968456
transform 1 0 76636 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_833
timestamp 1
transform 1 0 77740 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_839
timestamp 1
transform 1 0 78292 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_841
timestamp 1636968456
transform 1 0 78476 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_853
timestamp 1636968456
transform 1 0 79580 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_865
timestamp 1636968456
transform 1 0 80684 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_877
timestamp 1636968456
transform 1 0 81788 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_889
timestamp 1
transform 1 0 82892 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_895
timestamp 1
transform 1 0 83444 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_897
timestamp 1636968456
transform 1 0 83628 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_909
timestamp 1636968456
transform 1 0 84732 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_921
timestamp 1636968456
transform 1 0 85836 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_933
timestamp 1636968456
transform 1 0 86940 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_945
timestamp 1
transform 1 0 88044 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_951
timestamp 1
transform 1 0 88596 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_953
timestamp 1636968456
transform 1 0 88780 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_965
timestamp 1636968456
transform 1 0 89884 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_977
timestamp 1636968456
transform 1 0 90988 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_989
timestamp 1636968456
transform 1 0 92092 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_1001
timestamp 1
transform 1 0 93196 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_1007
timestamp 1
transform 1 0 93748 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1009
timestamp 1636968456
transform 1 0 93932 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1021
timestamp 1636968456
transform 1 0 95036 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1033
timestamp 1636968456
transform 1 0 96140 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1045
timestamp 1636968456
transform 1 0 97244 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_1057
timestamp 1
transform 1 0 98348 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_1063
timestamp 1
transform 1 0 98900 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1065
timestamp 1636968456
transform 1 0 99084 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1077
timestamp 1636968456
transform 1 0 100188 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1089
timestamp 1636968456
transform 1 0 101292 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1101
timestamp 1636968456
transform 1 0 102396 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_265_1113
timestamp 1
transform 1 0 103500 0 -1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_265_1119
timestamp 1
transform 1 0 104052 0 -1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1121
timestamp 1636968456
transform 1 0 104236 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1133
timestamp 1636968456
transform 1 0 105340 0 -1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_265_1145
timestamp 1636968456
transform 1 0 106444 0 -1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_265_1157
timestamp 1
transform 1 0 107548 0 -1 146880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_265_1165
timestamp 1
transform 1 0 108284 0 -1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_3
timestamp 1636968456
transform 1 0 1380 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_15
timestamp 1636968456
transform 1 0 2484 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_266_27
timestamp 1
transform 1 0 3588 0 1 146880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_266_29
timestamp 1636968456
transform 1 0 3772 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_41
timestamp 1636968456
transform 1 0 4876 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_53
timestamp 1
transform 1 0 5980 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_57
timestamp 1636968456
transform 1 0 6348 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_69
timestamp 1636968456
transform 1 0 7452 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_81
timestamp 1
transform 1 0 8556 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_85
timestamp 1636968456
transform 1 0 8924 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_97
timestamp 1636968456
transform 1 0 10028 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_109
timestamp 1
transform 1 0 11132 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_113
timestamp 1636968456
transform 1 0 11500 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_125
timestamp 1636968456
transform 1 0 12604 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_137
timestamp 1
transform 1 0 13708 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_141
timestamp 1636968456
transform 1 0 14076 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_153
timestamp 1636968456
transform 1 0 15180 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_165
timestamp 1
transform 1 0 16284 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_169
timestamp 1636968456
transform 1 0 16652 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_181
timestamp 1636968456
transform 1 0 17756 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_193
timestamp 1
transform 1 0 18860 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_197
timestamp 1636968456
transform 1 0 19228 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_209
timestamp 1636968456
transform 1 0 20332 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_221
timestamp 1
transform 1 0 21436 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_225
timestamp 1636968456
transform 1 0 21804 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_237
timestamp 1636968456
transform 1 0 22908 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_249
timestamp 1
transform 1 0 24012 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_253
timestamp 1636968456
transform 1 0 24380 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_265
timestamp 1636968456
transform 1 0 25484 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_277
timestamp 1
transform 1 0 26588 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_281
timestamp 1636968456
transform 1 0 26956 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_293
timestamp 1636968456
transform 1 0 28060 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_305
timestamp 1
transform 1 0 29164 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_309
timestamp 1636968456
transform 1 0 29532 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_321
timestamp 1636968456
transform 1 0 30636 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_333
timestamp 1
transform 1 0 31740 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_337
timestamp 1636968456
transform 1 0 32108 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_349
timestamp 1636968456
transform 1 0 33212 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_361
timestamp 1
transform 1 0 34316 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_365
timestamp 1636968456
transform 1 0 34684 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_377
timestamp 1636968456
transform 1 0 35788 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_389
timestamp 1
transform 1 0 36892 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_393
timestamp 1636968456
transform 1 0 37260 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_405
timestamp 1636968456
transform 1 0 38364 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_417
timestamp 1
transform 1 0 39468 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_421
timestamp 1636968456
transform 1 0 39836 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_433
timestamp 1636968456
transform 1 0 40940 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_445
timestamp 1
transform 1 0 42044 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_449
timestamp 1636968456
transform 1 0 42412 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_461
timestamp 1636968456
transform 1 0 43516 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_473
timestamp 1
transform 1 0 44620 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_477
timestamp 1636968456
transform 1 0 44988 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_489
timestamp 1636968456
transform 1 0 46092 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_501
timestamp 1
transform 1 0 47196 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_505
timestamp 1636968456
transform 1 0 47564 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_517
timestamp 1636968456
transform 1 0 48668 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_529
timestamp 1
transform 1 0 49772 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_533
timestamp 1636968456
transform 1 0 50140 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_545
timestamp 1636968456
transform 1 0 51244 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_557
timestamp 1
transform 1 0 52348 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_561
timestamp 1636968456
transform 1 0 52716 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_573
timestamp 1636968456
transform 1 0 53820 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_585
timestamp 1
transform 1 0 54924 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_589
timestamp 1636968456
transform 1 0 55292 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_601
timestamp 1636968456
transform 1 0 56396 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_613
timestamp 1
transform 1 0 57500 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_617
timestamp 1636968456
transform 1 0 57868 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_629
timestamp 1636968456
transform 1 0 58972 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_641
timestamp 1
transform 1 0 60076 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_645
timestamp 1636968456
transform 1 0 60444 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_657
timestamp 1636968456
transform 1 0 61548 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_669
timestamp 1
transform 1 0 62652 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_673
timestamp 1636968456
transform 1 0 63020 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_685
timestamp 1636968456
transform 1 0 64124 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_697
timestamp 1
transform 1 0 65228 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_701
timestamp 1636968456
transform 1 0 65596 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_713
timestamp 1636968456
transform 1 0 66700 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_725
timestamp 1
transform 1 0 67804 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_729
timestamp 1636968456
transform 1 0 68172 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_741
timestamp 1636968456
transform 1 0 69276 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_753
timestamp 1
transform 1 0 70380 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_757
timestamp 1636968456
transform 1 0 70748 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_769
timestamp 1636968456
transform 1 0 71852 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_781
timestamp 1
transform 1 0 72956 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_785
timestamp 1636968456
transform 1 0 73324 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_797
timestamp 1636968456
transform 1 0 74428 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_809
timestamp 1
transform 1 0 75532 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_813
timestamp 1636968456
transform 1 0 75900 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_825
timestamp 1636968456
transform 1 0 77004 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_837
timestamp 1
transform 1 0 78108 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_841
timestamp 1636968456
transform 1 0 78476 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_853
timestamp 1636968456
transform 1 0 79580 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_865
timestamp 1
transform 1 0 80684 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_869
timestamp 1636968456
transform 1 0 81052 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_881
timestamp 1636968456
transform 1 0 82156 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_893
timestamp 1
transform 1 0 83260 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_897
timestamp 1636968456
transform 1 0 83628 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_909
timestamp 1636968456
transform 1 0 84732 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_921
timestamp 1
transform 1 0 85836 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_925
timestamp 1636968456
transform 1 0 86204 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_937
timestamp 1636968456
transform 1 0 87308 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_949
timestamp 1
transform 1 0 88412 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_953
timestamp 1636968456
transform 1 0 88780 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_965
timestamp 1636968456
transform 1 0 89884 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_977
timestamp 1
transform 1 0 90988 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_981
timestamp 1636968456
transform 1 0 91356 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_993
timestamp 1636968456
transform 1 0 92460 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1005
timestamp 1
transform 1 0 93564 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1009
timestamp 1636968456
transform 1 0 93932 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1021
timestamp 1636968456
transform 1 0 95036 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1033
timestamp 1
transform 1 0 96140 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1037
timestamp 1636968456
transform 1 0 96508 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1049
timestamp 1636968456
transform 1 0 97612 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1061
timestamp 1
transform 1 0 98716 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1065
timestamp 1636968456
transform 1 0 99084 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1077
timestamp 1636968456
transform 1 0 100188 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1089
timestamp 1
transform 1 0 101292 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1093
timestamp 1636968456
transform 1 0 101660 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1105
timestamp 1636968456
transform 1 0 102764 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1117
timestamp 1
transform 1 0 103868 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1121
timestamp 1636968456
transform 1 0 104236 0 1 146880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1133
timestamp 1636968456
transform 1 0 105340 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_266_1145
timestamp 1
transform 1 0 106444 0 1 146880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_266_1149
timestamp 1636968456
transform 1 0 106812 0 1 146880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_266_1161
timestamp 1
transform 1 0 107916 0 1 146880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_266_1167
timestamp 1
transform 1 0 108468 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1
transform -1 0 2300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1
transform 1 0 1380 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1
transform 1 0 1380 0 1 80512
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1
transform 1 0 1380 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1
transform 1 0 1380 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1
transform 1 0 1380 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1
transform 1 0 1380 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1
transform 1 0 1380 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1
transform 1 0 1380 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1
transform 1 0 1380 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1
transform 1 0 108284 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1
transform -1 0 108560 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1
transform -1 0 108560 0 1 80512
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1
transform -1 0 108560 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1
transform -1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1
transform 1 0 41952 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1
transform 1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1
transform -1 0 31924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1
transform -1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1
transform -1 0 34500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1
transform 1 0 1380 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1
transform 1 0 1380 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1
transform 1 0 1380 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1
transform 1 0 1380 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1
transform 1 0 1380 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1
transform 1 0 1380 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1
transform 1 0 1380 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1
transform 1 0 1380 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1
transform 1 0 1380 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1
transform 1 0 1380 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1
transform 1 0 1380 0 -1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1
transform 1 0 1380 0 1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1
transform 1 0 1380 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1
transform 1 0 1380 0 -1 88128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1
transform 1 0 1380 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1
transform 1 0 1380 0 -1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1
transform -1 0 108560 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1
transform 1 0 108284 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1
transform 1 0 108284 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1
transform -1 0 108560 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1
transform -1 0 108560 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap76
timestamp 1
transform -1 0 101568 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  max_cap77
timestamp 1
transform 1 0 101292 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap79
timestamp 1
transform -1 0 97336 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap80
timestamp 1
transform -1 0 99360 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap82
timestamp 1
transform 1 0 99544 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap84
timestamp 1
transform -1 0 101200 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap85
timestamp 1
transform -1 0 105064 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap86
timestamp 1
transform 1 0 105984 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i0_114
timestamp 1
transform -1 0 104604 0 1 59840
box -38 -48 314 592
use ram256x16  mem_i0
timestamp 0
transform 1 0 10000 0 1 10000
box 0 0 1 1
use sky130_fd_sc_hd__conb_1  mem_i1_115
timestamp 1
transform -1 0 104604 0 1 129472
box -38 -48 314 592
use ram256x16  mem_i1
timestamp 0
transform 1 0 10000 0 1 80000
box 0 0 1 1
use sky130_fd_sc_hd__buf_2  output60
timestamp 1
transform -1 0 1748 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1
transform 1 0 108192 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1
transform 1 0 108192 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1
transform 1 0 108192 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1
transform 1 0 108192 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1
transform 1 0 108192 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1
transform 1 0 108192 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1
transform -1 0 1748 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1
transform -1 0 1748 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1
transform -1 0 1748 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1
transform -1 0 1748 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1
transform -1 0 1748 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1
transform -1 0 1748 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1
transform 1 0 108192 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1
transform 1 0 108192 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1
transform 1 0 108192 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_267
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 108836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_268
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 108836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_269
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 108836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_270
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 108836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_271
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 108836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_272
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 108836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_273
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 108836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_274
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 108836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_275
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 108836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_276
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 108836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_533
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_747
timestamp 1
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_534
timestamp 1
transform 1 0 104052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_53
timestamp 1
transform -1 0 108836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_277
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_641
timestamp 1
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_535
timestamp 1
transform 1 0 104052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_54
timestamp 1
transform -1 0 108836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_278
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_642
timestamp 1
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_536
timestamp 1
transform 1 0 104052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_55
timestamp 1
transform -1 0 108836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_279
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_643
timestamp 1
transform -1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_537
timestamp 1
transform 1 0 104052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_56
timestamp 1
transform -1 0 108836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_280
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_644
timestamp 1
transform -1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_538
timestamp 1
transform 1 0 104052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_57
timestamp 1
transform -1 0 108836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_281
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_645
timestamp 1
transform -1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_539
timestamp 1
transform 1 0 104052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_58
timestamp 1
transform -1 0 108836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_282
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_646
timestamp 1
transform -1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_540
timestamp 1
transform 1 0 104052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_59
timestamp 1
transform -1 0 108836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_283
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_647
timestamp 1
transform -1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_541
timestamp 1
transform 1 0 104052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_60
timestamp 1
transform -1 0 108836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_284
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_648
timestamp 1
transform -1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_542
timestamp 1
transform 1 0 104052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_61
timestamp 1
transform -1 0 108836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_285
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_649
timestamp 1
transform -1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_543
timestamp 1
transform 1 0 104052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_62
timestamp 1
transform -1 0 108836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_286
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_650
timestamp 1
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_544
timestamp 1
transform 1 0 104052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_63
timestamp 1
transform -1 0 108836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_287
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_651
timestamp 1
transform -1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_545
timestamp 1
transform 1 0 104052 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_64
timestamp 1
transform -1 0 108836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_288
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_652
timestamp 1
transform -1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_546
timestamp 1
transform 1 0 104052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_65
timestamp 1
transform -1 0 108836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_289
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_653
timestamp 1
transform -1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_547
timestamp 1
transform 1 0 104052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_66
timestamp 1
transform -1 0 108836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_290
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_654
timestamp 1
transform -1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_548
timestamp 1
transform 1 0 104052 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_67
timestamp 1
transform -1 0 108836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_291
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_655
timestamp 1
transform -1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_549
timestamp 1
transform 1 0 104052 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_68
timestamp 1
transform -1 0 108836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_292
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_656
timestamp 1
transform -1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_550
timestamp 1
transform 1 0 104052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_69
timestamp 1
transform -1 0 108836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_293
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_657
timestamp 1
transform -1 0 7912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_551
timestamp 1
transform 1 0 104052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_70
timestamp 1
transform -1 0 108836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_294
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_658
timestamp 1
transform -1 0 7912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_552
timestamp 1
transform 1 0 104052 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_71
timestamp 1
transform -1 0 108836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_295
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_659
timestamp 1
transform -1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_553
timestamp 1
transform 1 0 104052 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_72
timestamp 1
transform -1 0 108836 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_296
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_660
timestamp 1
transform -1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_554
timestamp 1
transform 1 0 104052 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_73
timestamp 1
transform -1 0 108836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_297
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_661
timestamp 1
transform -1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_555
timestamp 1
transform 1 0 104052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_74
timestamp 1
transform -1 0 108836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_298
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_662
timestamp 1
transform -1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_556
timestamp 1
transform 1 0 104052 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_75
timestamp 1
transform -1 0 108836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_299
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_663
timestamp 1
transform -1 0 7912 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_557
timestamp 1
transform 1 0 104052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_76
timestamp 1
transform -1 0 108836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_300
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_664
timestamp 1
transform -1 0 7912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_558
timestamp 1
transform 1 0 104052 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_77
timestamp 1
transform -1 0 108836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_301
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_665
timestamp 1
transform -1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_559
timestamp 1
transform 1 0 104052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_78
timestamp 1
transform -1 0 108836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_302
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_666
timestamp 1
transform -1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_560
timestamp 1
transform 1 0 104052 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_79
timestamp 1
transform -1 0 108836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_303
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_667
timestamp 1
transform -1 0 7912 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_561
timestamp 1
transform 1 0 104052 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_80
timestamp 1
transform -1 0 108836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_304
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_668
timestamp 1
transform -1 0 7912 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_562
timestamp 1
transform 1 0 104052 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_81
timestamp 1
transform -1 0 108836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_305
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_669
timestamp 1
transform -1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_563
timestamp 1
transform 1 0 104052 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_82
timestamp 1
transform -1 0 108836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_306
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_670
timestamp 1
transform -1 0 7912 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_564
timestamp 1
transform 1 0 104052 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_83
timestamp 1
transform -1 0 108836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_307
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_671
timestamp 1
transform -1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_565
timestamp 1
transform 1 0 104052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_84
timestamp 1
transform -1 0 108836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_308
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_672
timestamp 1
transform -1 0 7912 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_566
timestamp 1
transform 1 0 104052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_85
timestamp 1
transform -1 0 108836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_309
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_673
timestamp 1
transform -1 0 7912 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_567
timestamp 1
transform 1 0 104052 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_86
timestamp 1
transform -1 0 108836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_310
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_674
timestamp 1
transform -1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_568
timestamp 1
transform 1 0 104052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_87
timestamp 1
transform -1 0 108836 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_311
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_675
timestamp 1
transform -1 0 7912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_569
timestamp 1
transform 1 0 104052 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_88
timestamp 1
transform -1 0 108836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_312
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_676
timestamp 1
transform -1 0 7912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_570
timestamp 1
transform 1 0 104052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_89
timestamp 1
transform -1 0 108836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_313
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_677
timestamp 1
transform -1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_571
timestamp 1
transform 1 0 104052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_90
timestamp 1
transform -1 0 108836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_314
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_678
timestamp 1
transform -1 0 7912 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_572
timestamp 1
transform 1 0 104052 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_91
timestamp 1
transform -1 0 108836 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_315
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_679
timestamp 1
transform -1 0 7912 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_573
timestamp 1
transform 1 0 104052 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_92
timestamp 1
transform -1 0 108836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_316
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_680
timestamp 1
transform -1 0 7912 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_574
timestamp 1
transform 1 0 104052 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_93
timestamp 1
transform -1 0 108836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_317
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_681
timestamp 1
transform -1 0 7912 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_575
timestamp 1
transform 1 0 104052 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_94
timestamp 1
transform -1 0 108836 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_318
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_682
timestamp 1
transform -1 0 7912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_576
timestamp 1
transform 1 0 104052 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_95
timestamp 1
transform -1 0 108836 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_319
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_683
timestamp 1
transform -1 0 7912 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_577
timestamp 1
transform 1 0 104052 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_96
timestamp 1
transform -1 0 108836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_320
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_684
timestamp 1
transform -1 0 7912 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_578
timestamp 1
transform 1 0 104052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_97
timestamp 1
transform -1 0 108836 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_321
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_685
timestamp 1
transform -1 0 7912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_579
timestamp 1
transform 1 0 104052 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_98
timestamp 1
transform -1 0 108836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_322
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_686
timestamp 1
transform -1 0 7912 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_580
timestamp 1
transform 1 0 104052 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_99
timestamp 1
transform -1 0 108836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_323
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_687
timestamp 1
transform -1 0 7912 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_581
timestamp 1
transform 1 0 104052 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_100
timestamp 1
transform -1 0 108836 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_324
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_688
timestamp 1
transform -1 0 7912 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_582
timestamp 1
transform 1 0 104052 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_101
timestamp 1
transform -1 0 108836 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_325
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_689
timestamp 1
transform -1 0 7912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_583
timestamp 1
transform 1 0 104052 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_102
timestamp 1
transform -1 0 108836 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_326
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_690
timestamp 1
transform -1 0 7912 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_584
timestamp 1
transform 1 0 104052 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_103
timestamp 1
transform -1 0 108836 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_327
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_691
timestamp 1
transform -1 0 7912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_585
timestamp 1
transform 1 0 104052 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_104
timestamp 1
transform -1 0 108836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_328
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_692
timestamp 1
transform -1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_586
timestamp 1
transform 1 0 104052 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_105
timestamp 1
transform -1 0 108836 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_329
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_693
timestamp 1
transform -1 0 7912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_587
timestamp 1
transform 1 0 104052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_106
timestamp 1
transform -1 0 108836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_330
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_694
timestamp 1
transform -1 0 7912 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_588
timestamp 1
transform 1 0 104052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_107
timestamp 1
transform -1 0 108836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_331
timestamp 1
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_695
timestamp 1
transform -1 0 7912 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_589
timestamp 1
transform 1 0 104052 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_108
timestamp 1
transform -1 0 108836 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_332
timestamp 1
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_696
timestamp 1
transform -1 0 7912 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_590
timestamp 1
transform 1 0 104052 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_109
timestamp 1
transform -1 0 108836 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_333
timestamp 1
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_697
timestamp 1
transform -1 0 7912 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_591
timestamp 1
transform 1 0 104052 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_110
timestamp 1
transform -1 0 108836 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_334
timestamp 1
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_698
timestamp 1
transform -1 0 7912 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_592
timestamp 1
transform 1 0 104052 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_111
timestamp 1
transform -1 0 108836 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_335
timestamp 1
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_699
timestamp 1
transform -1 0 7912 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_593
timestamp 1
transform 1 0 104052 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_112
timestamp 1
transform -1 0 108836 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_336
timestamp 1
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_700
timestamp 1
transform -1 0 7912 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_594
timestamp 1
transform 1 0 104052 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_113
timestamp 1
transform -1 0 108836 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_337
timestamp 1
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_701
timestamp 1
transform -1 0 7912 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_595
timestamp 1
transform 1 0 104052 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_114
timestamp 1
transform -1 0 108836 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_338
timestamp 1
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_702
timestamp 1
transform -1 0 7912 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_596
timestamp 1
transform 1 0 104052 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_115
timestamp 1
transform -1 0 108836 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_339
timestamp 1
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_703
timestamp 1
transform -1 0 7912 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_597
timestamp 1
transform 1 0 104052 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_116
timestamp 1
transform -1 0 108836 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_340
timestamp 1
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_704
timestamp 1
transform -1 0 7912 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_598
timestamp 1
transform 1 0 104052 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_117
timestamp 1
transform -1 0 108836 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_341
timestamp 1
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_705
timestamp 1
transform -1 0 7912 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_599
timestamp 1
transform 1 0 104052 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_118
timestamp 1
transform -1 0 108836 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_342
timestamp 1
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_706
timestamp 1
transform -1 0 7912 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_600
timestamp 1
transform 1 0 104052 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_119
timestamp 1
transform -1 0 108836 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_343
timestamp 1
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_707
timestamp 1
transform -1 0 7912 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_601
timestamp 1
transform 1 0 104052 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_120
timestamp 1
transform -1 0 108836 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_344
timestamp 1
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_708
timestamp 1
transform -1 0 7912 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_602
timestamp 1
transform 1 0 104052 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_121
timestamp 1
transform -1 0 108836 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_345
timestamp 1
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_709
timestamp 1
transform -1 0 7912 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_603
timestamp 1
transform 1 0 104052 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_122
timestamp 1
transform -1 0 108836 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_346
timestamp 1
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_710
timestamp 1
transform -1 0 7912 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_604
timestamp 1
transform 1 0 104052 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_123
timestamp 1
transform -1 0 108836 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_347
timestamp 1
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_711
timestamp 1
transform -1 0 7912 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_605
timestamp 1
transform 1 0 104052 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_124
timestamp 1
transform -1 0 108836 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_348
timestamp 1
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_712
timestamp 1
transform -1 0 7912 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_606
timestamp 1
transform 1 0 104052 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_125
timestamp 1
transform -1 0 108836 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_349
timestamp 1
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_713
timestamp 1
transform -1 0 7912 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_607
timestamp 1
transform 1 0 104052 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_126
timestamp 1
transform -1 0 108836 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_350
timestamp 1
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_714
timestamp 1
transform -1 0 7912 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_608
timestamp 1
transform 1 0 104052 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_127
timestamp 1
transform -1 0 108836 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_351
timestamp 1
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_715
timestamp 1
transform -1 0 7912 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_609
timestamp 1
transform 1 0 104052 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_128
timestamp 1
transform -1 0 108836 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_352
timestamp 1
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_716
timestamp 1
transform -1 0 7912 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_610
timestamp 1
transform 1 0 104052 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_129
timestamp 1
transform -1 0 108836 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_353
timestamp 1
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_717
timestamp 1
transform -1 0 7912 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_611
timestamp 1
transform 1 0 104052 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_130
timestamp 1
transform -1 0 108836 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_354
timestamp 1
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_718
timestamp 1
transform -1 0 7912 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_612
timestamp 1
transform 1 0 104052 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_131
timestamp 1
transform -1 0 108836 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_355
timestamp 1
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_719
timestamp 1
transform -1 0 7912 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_613
timestamp 1
transform 1 0 104052 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_132
timestamp 1
transform -1 0 108836 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_356
timestamp 1
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_720
timestamp 1
transform -1 0 7912 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_614
timestamp 1
transform 1 0 104052 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_133
timestamp 1
transform -1 0 108836 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_357
timestamp 1
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_721
timestamp 1
transform -1 0 7912 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_615
timestamp 1
transform 1 0 104052 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_134
timestamp 1
transform -1 0 108836 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_358
timestamp 1
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_722
timestamp 1
transform -1 0 7912 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_616
timestamp 1
transform 1 0 104052 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_135
timestamp 1
transform -1 0 108836 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_359
timestamp 1
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_723
timestamp 1
transform -1 0 7912 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_617
timestamp 1
transform 1 0 104052 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_136
timestamp 1
transform -1 0 108836 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_360
timestamp 1
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_724
timestamp 1
transform -1 0 7912 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_618
timestamp 1
transform 1 0 104052 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_137
timestamp 1
transform -1 0 108836 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_361
timestamp 1
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_725
timestamp 1
transform -1 0 7912 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_619
timestamp 1
transform 1 0 104052 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_138
timestamp 1
transform -1 0 108836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_362
timestamp 1
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_726
timestamp 1
transform -1 0 7912 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_620
timestamp 1
transform 1 0 104052 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_139
timestamp 1
transform -1 0 108836 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_363
timestamp 1
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_727
timestamp 1
transform -1 0 7912 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_621
timestamp 1
transform 1 0 104052 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_140
timestamp 1
transform -1 0 108836 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_364
timestamp 1
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_728
timestamp 1
transform -1 0 7912 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_622
timestamp 1
transform 1 0 104052 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_141
timestamp 1
transform -1 0 108836 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_365
timestamp 1
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_729
timestamp 1
transform -1 0 7912 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_623
timestamp 1
transform 1 0 104052 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_142
timestamp 1
transform -1 0 108836 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_366
timestamp 1
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_730
timestamp 1
transform -1 0 7912 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_624
timestamp 1
transform 1 0 104052 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_143
timestamp 1
transform -1 0 108836 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_367
timestamp 1
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_731
timestamp 1
transform -1 0 7912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_625
timestamp 1
transform 1 0 104052 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_144
timestamp 1
transform -1 0 108836 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_368
timestamp 1
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_732
timestamp 1
transform -1 0 7912 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_626
timestamp 1
transform 1 0 104052 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_145
timestamp 1
transform -1 0 108836 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_369
timestamp 1
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_733
timestamp 1
transform -1 0 7912 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_627
timestamp 1
transform 1 0 104052 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_146
timestamp 1
transform -1 0 108836 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_370
timestamp 1
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_734
timestamp 1
transform -1 0 7912 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_628
timestamp 1
transform 1 0 104052 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_147
timestamp 1
transform -1 0 108836 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_371
timestamp 1
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_735
timestamp 1
transform -1 0 7912 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_629
timestamp 1
transform 1 0 104052 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_148
timestamp 1
transform -1 0 108836 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_372
timestamp 1
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_736
timestamp 1
transform -1 0 7912 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_630
timestamp 1
transform 1 0 104052 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_149
timestamp 1
transform -1 0 108836 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_373
timestamp 1
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_737
timestamp 1
transform -1 0 7912 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_631
timestamp 1
transform 1 0 104052 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_150
timestamp 1
transform -1 0 108836 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_374
timestamp 1
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_738
timestamp 1
transform -1 0 7912 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_632
timestamp 1
transform 1 0 104052 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_151
timestamp 1
transform -1 0 108836 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_375
timestamp 1
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_739
timestamp 1
transform -1 0 7912 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_633
timestamp 1
transform 1 0 104052 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_152
timestamp 1
transform -1 0 108836 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_376
timestamp 1
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_740
timestamp 1
transform -1 0 7912 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_634
timestamp 1
transform 1 0 104052 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_153
timestamp 1
transform -1 0 108836 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_377
timestamp 1
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_741
timestamp 1
transform -1 0 7912 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_635
timestamp 1
transform 1 0 104052 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_154
timestamp 1
transform -1 0 108836 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_378
timestamp 1
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_742
timestamp 1
transform -1 0 7912 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_636
timestamp 1
transform 1 0 104052 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_155
timestamp 1
transform -1 0 108836 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_379
timestamp 1
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_743
timestamp 1
transform -1 0 7912 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_637
timestamp 1
transform 1 0 104052 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_156
timestamp 1
transform -1 0 108836 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_380
timestamp 1
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_744
timestamp 1
transform -1 0 7912 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_638
timestamp 1
transform 1 0 104052 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_157
timestamp 1
transform -1 0 108836 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_381
timestamp 1
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_745
timestamp 1
transform -1 0 7912 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_639
timestamp 1
transform 1 0 104052 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_158
timestamp 1
transform -1 0 108836 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_382
timestamp 1
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_746
timestamp 1
transform -1 0 7912 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_640
timestamp 1
transform 1 0 104052 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_159
timestamp 1
transform -1 0 108836 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_384
timestamp 1
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_10
timestamp 1
transform -1 0 108836 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_385
timestamp 1
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_11
timestamp 1
transform -1 0 108836 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_386
timestamp 1
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_12
timestamp 1
transform -1 0 108836 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_387
timestamp 1
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_13
timestamp 1
transform -1 0 108836 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_388
timestamp 1
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_14
timestamp 1
transform -1 0 108836 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_389
timestamp 1
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_15
timestamp 1
transform -1 0 108836 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_390
timestamp 1
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_16
timestamp 1
transform -1 0 108836 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Left_391
timestamp 1
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Right_17
timestamp 1
transform -1 0 108836 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Left_392
timestamp 1
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Right_18
timestamp 1
transform -1 0 108836 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Left_393
timestamp 1
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Right_19
timestamp 1
transform -1 0 108836 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Left_394
timestamp 1
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Right_20
timestamp 1
transform -1 0 108836 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Left_395
timestamp 1
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Right_21
timestamp 1
transform -1 0 108836 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Left_396
timestamp 1
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Right_22
timestamp 1
transform -1 0 108836 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Left_397
timestamp 1
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Right_23
timestamp 1
transform -1 0 108836 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Left_398
timestamp 1
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Right_24
timestamp 1
transform -1 0 108836 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Left_399
timestamp 1
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Right_25
timestamp 1
transform -1 0 108836 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Left_400
timestamp 1
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Right_26
timestamp 1
transform -1 0 108836 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Left_401
timestamp 1
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Right_27
timestamp 1
transform -1 0 108836 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Left_402
timestamp 1
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Right_28
timestamp 1
transform -1 0 108836 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Left_403
timestamp 1
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Right_29
timestamp 1
transform -1 0 108836 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Left_404
timestamp 1
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Right_30
timestamp 1
transform -1 0 108836 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Left_405
timestamp 1
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Right_31
timestamp 1
transform -1 0 108836 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_383
timestamp 1
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_855
timestamp 1
transform -1 0 7912 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Left_748
timestamp 1
transform 1 0 104052 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Right_160
timestamp 1
transform -1 0 108836 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_406
timestamp 1
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_856
timestamp 1
transform -1 0 7912 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Left_749
timestamp 1
transform 1 0 104052 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Right_161
timestamp 1
transform -1 0 108836 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_407
timestamp 1
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_857
timestamp 1
transform -1 0 7912 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Left_750
timestamp 1
transform 1 0 104052 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Right_162
timestamp 1
transform -1 0 108836 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_408
timestamp 1
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_858
timestamp 1
transform -1 0 7912 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Left_751
timestamp 1
transform 1 0 104052 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Right_163
timestamp 1
transform -1 0 108836 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_409
timestamp 1
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_859
timestamp 1
transform -1 0 7912 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Left_752
timestamp 1
transform 1 0 104052 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Right_164
timestamp 1
transform -1 0 108836 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_410
timestamp 1
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_860
timestamp 1
transform -1 0 7912 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Left_753
timestamp 1
transform 1 0 104052 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Right_165
timestamp 1
transform -1 0 108836 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_411
timestamp 1
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_861
timestamp 1
transform -1 0 7912 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Left_754
timestamp 1
transform 1 0 104052 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Right_166
timestamp 1
transform -1 0 108836 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Left_412
timestamp 1
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Right_862
timestamp 1
transform -1 0 7912 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Left_755
timestamp 1
transform 1 0 104052 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Right_167
timestamp 1
transform -1 0 108836 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Left_413
timestamp 1
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Right_863
timestamp 1
transform -1 0 7912 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Left_756
timestamp 1
transform 1 0 104052 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Right_168
timestamp 1
transform -1 0 108836 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Left_414
timestamp 1
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Right_864
timestamp 1
transform -1 0 7912 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Left_757
timestamp 1
transform 1 0 104052 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Right_169
timestamp 1
transform -1 0 108836 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Left_415
timestamp 1
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Right_865
timestamp 1
transform -1 0 7912 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Left_758
timestamp 1
transform 1 0 104052 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Right_170
timestamp 1
transform -1 0 108836 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Left_416
timestamp 1
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_1_Right_866
timestamp 1
transform -1 0 7912 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Left_759
timestamp 1
transform 1 0 104052 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Right_171
timestamp 1
transform -1 0 108836 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Left_417
timestamp 1
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_1_Right_867
timestamp 1
transform -1 0 7912 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Left_760
timestamp 1
transform 1 0 104052 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Right_172
timestamp 1
transform -1 0 108836 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Left_418
timestamp 1
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_1_Right_868
timestamp 1
transform -1 0 7912 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Left_761
timestamp 1
transform 1 0 104052 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Right_173
timestamp 1
transform -1 0 108836 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Left_419
timestamp 1
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_1_Right_869
timestamp 1
transform -1 0 7912 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Left_762
timestamp 1
transform 1 0 104052 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Right_174
timestamp 1
transform -1 0 108836 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Left_420
timestamp 1
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_1_Right_870
timestamp 1
transform -1 0 7912 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Left_763
timestamp 1
transform 1 0 104052 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Right_175
timestamp 1
transform -1 0 108836 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Left_421
timestamp 1
transform 1 0 1104 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_1_Right_871
timestamp 1
transform -1 0 7912 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Left_764
timestamp 1
transform 1 0 104052 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Right_176
timestamp 1
transform -1 0 108836 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Left_422
timestamp 1
transform 1 0 1104 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_1_Right_872
timestamp 1
transform -1 0 7912 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_2_Left_765
timestamp 1
transform 1 0 104052 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_2_Right_177
timestamp 1
transform -1 0 108836 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Left_423
timestamp 1
transform 1 0 1104 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_1_Right_873
timestamp 1
transform -1 0 7912 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_2_Left_766
timestamp 1
transform 1 0 104052 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_2_Right_178
timestamp 1
transform -1 0 108836 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Left_424
timestamp 1
transform 1 0 1104 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_1_Right_874
timestamp 1
transform -1 0 7912 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_2_Left_767
timestamp 1
transform 1 0 104052 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_2_Right_179
timestamp 1
transform -1 0 108836 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Left_425
timestamp 1
transform 1 0 1104 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_1_Right_875
timestamp 1
transform -1 0 7912 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_2_Left_768
timestamp 1
transform 1 0 104052 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_2_Right_180
timestamp 1
transform -1 0 108836 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Left_426
timestamp 1
transform 1 0 1104 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_1_Right_876
timestamp 1
transform -1 0 7912 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_2_Left_769
timestamp 1
transform 1 0 104052 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_2_Right_181
timestamp 1
transform -1 0 108836 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Left_427
timestamp 1
transform 1 0 1104 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_1_Right_877
timestamp 1
transform -1 0 7912 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_2_Left_770
timestamp 1
transform 1 0 104052 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_2_Right_182
timestamp 1
transform -1 0 108836 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Left_428
timestamp 1
transform 1 0 1104 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_1_Right_878
timestamp 1
transform -1 0 7912 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_2_Left_771
timestamp 1
transform 1 0 104052 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_2_Right_183
timestamp 1
transform -1 0 108836 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Left_429
timestamp 1
transform 1 0 1104 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_1_Right_879
timestamp 1
transform -1 0 7912 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_2_Left_772
timestamp 1
transform 1 0 104052 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_2_Right_184
timestamp 1
transform -1 0 108836 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Left_430
timestamp 1
transform 1 0 1104 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_1_Right_880
timestamp 1
transform -1 0 7912 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_2_Left_773
timestamp 1
transform 1 0 104052 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_2_Right_185
timestamp 1
transform -1 0 108836 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_1_Left_431
timestamp 1
transform 1 0 1104 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_1_Right_881
timestamp 1
transform -1 0 7912 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_2_Left_774
timestamp 1
transform 1 0 104052 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_2_Right_186
timestamp 1
transform -1 0 108836 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_1_Left_432
timestamp 1
transform 1 0 1104 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_1_Right_882
timestamp 1
transform -1 0 7912 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_2_Left_775
timestamp 1
transform 1 0 104052 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_2_Right_187
timestamp 1
transform -1 0 108836 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_1_Left_433
timestamp 1
transform 1 0 1104 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_1_Right_883
timestamp 1
transform -1 0 7912 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_2_Left_776
timestamp 1
transform 1 0 104052 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_2_Right_188
timestamp 1
transform -1 0 108836 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_1_Left_434
timestamp 1
transform 1 0 1104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_1_Right_884
timestamp 1
transform -1 0 7912 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_2_Left_777
timestamp 1
transform 1 0 104052 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_2_Right_189
timestamp 1
transform -1 0 108836 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_1_Left_435
timestamp 1
transform 1 0 1104 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_1_Right_885
timestamp 1
transform -1 0 7912 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_2_Left_778
timestamp 1
transform 1 0 104052 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_2_Right_190
timestamp 1
transform -1 0 108836 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_1_Left_436
timestamp 1
transform 1 0 1104 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_1_Right_886
timestamp 1
transform -1 0 7912 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_2_Left_779
timestamp 1
transform 1 0 104052 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_2_Right_191
timestamp 1
transform -1 0 108836 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_1_Left_437
timestamp 1
transform 1 0 1104 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_1_Right_887
timestamp 1
transform -1 0 7912 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_2_Left_780
timestamp 1
transform 1 0 104052 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_2_Right_192
timestamp 1
transform -1 0 108836 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_1_Left_438
timestamp 1
transform 1 0 1104 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_1_Right_888
timestamp 1
transform -1 0 7912 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_2_Left_781
timestamp 1
transform 1 0 104052 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_2_Right_193
timestamp 1
transform -1 0 108836 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_1_Left_439
timestamp 1
transform 1 0 1104 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_1_Right_889
timestamp 1
transform -1 0 7912 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_2_Left_782
timestamp 1
transform 1 0 104052 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_2_Right_194
timestamp 1
transform -1 0 108836 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_1_Left_440
timestamp 1
transform 1 0 1104 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_1_Right_890
timestamp 1
transform -1 0 7912 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_2_Left_783
timestamp 1
transform 1 0 104052 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_2_Right_195
timestamp 1
transform -1 0 108836 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_1_Left_441
timestamp 1
transform 1 0 1104 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_1_Right_891
timestamp 1
transform -1 0 7912 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_2_Left_784
timestamp 1
transform 1 0 104052 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_2_Right_196
timestamp 1
transform -1 0 108836 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_1_Left_442
timestamp 1
transform 1 0 1104 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_1_Right_892
timestamp 1
transform -1 0 7912 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_2_Left_785
timestamp 1
transform 1 0 104052 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_2_Right_197
timestamp 1
transform -1 0 108836 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_1_Left_443
timestamp 1
transform 1 0 1104 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_1_Right_893
timestamp 1
transform -1 0 7912 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_2_Left_786
timestamp 1
transform 1 0 104052 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_2_Right_198
timestamp 1
transform -1 0 108836 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_1_Left_444
timestamp 1
transform 1 0 1104 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_1_Right_894
timestamp 1
transform -1 0 7912 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_2_Left_787
timestamp 1
transform 1 0 104052 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_2_Right_199
timestamp 1
transform -1 0 108836 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_1_Left_445
timestamp 1
transform 1 0 1104 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_1_Right_895
timestamp 1
transform -1 0 7912 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_2_Left_788
timestamp 1
transform 1 0 104052 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_2_Right_200
timestamp 1
transform -1 0 108836 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_1_Left_446
timestamp 1
transform 1 0 1104 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_1_Right_896
timestamp 1
transform -1 0 7912 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_2_Left_789
timestamp 1
transform 1 0 104052 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_2_Right_201
timestamp 1
transform -1 0 108836 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_1_Left_447
timestamp 1
transform 1 0 1104 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_1_Right_897
timestamp 1
transform -1 0 7912 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_2_Left_790
timestamp 1
transform 1 0 104052 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_2_Right_202
timestamp 1
transform -1 0 108836 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_1_Left_448
timestamp 1
transform 1 0 1104 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_1_Right_898
timestamp 1
transform -1 0 7912 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_2_Left_791
timestamp 1
transform 1 0 104052 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_2_Right_203
timestamp 1
transform -1 0 108836 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_1_Left_449
timestamp 1
transform 1 0 1104 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_1_Right_899
timestamp 1
transform -1 0 7912 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_2_Left_792
timestamp 1
transform 1 0 104052 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_183_2_Right_204
timestamp 1
transform -1 0 108836 0 -1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_1_Left_450
timestamp 1
transform 1 0 1104 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_1_Right_900
timestamp 1
transform -1 0 7912 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_2_Left_793
timestamp 1
transform 1 0 104052 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_184_2_Right_205
timestamp 1
transform -1 0 108836 0 1 102272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_1_Left_451
timestamp 1
transform 1 0 1104 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_1_Right_901
timestamp 1
transform -1 0 7912 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_2_Left_794
timestamp 1
transform 1 0 104052 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_185_2_Right_206
timestamp 1
transform -1 0 108836 0 -1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_1_Left_452
timestamp 1
transform 1 0 1104 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_1_Right_902
timestamp 1
transform -1 0 7912 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_2_Left_795
timestamp 1
transform 1 0 104052 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_186_2_Right_207
timestamp 1
transform -1 0 108836 0 1 103360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_1_Left_453
timestamp 1
transform 1 0 1104 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_1_Right_903
timestamp 1
transform -1 0 7912 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_2_Left_796
timestamp 1
transform 1 0 104052 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_187_2_Right_208
timestamp 1
transform -1 0 108836 0 -1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_1_Left_454
timestamp 1
transform 1 0 1104 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_1_Right_904
timestamp 1
transform -1 0 7912 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_2_Left_797
timestamp 1
transform 1 0 104052 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_188_2_Right_209
timestamp 1
transform -1 0 108836 0 1 104448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_1_Left_455
timestamp 1
transform 1 0 1104 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_1_Right_905
timestamp 1
transform -1 0 7912 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_2_Left_798
timestamp 1
transform 1 0 104052 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_189_2_Right_210
timestamp 1
transform -1 0 108836 0 -1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_1_Left_456
timestamp 1
transform 1 0 1104 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_1_Right_906
timestamp 1
transform -1 0 7912 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_2_Left_799
timestamp 1
transform 1 0 104052 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_190_2_Right_211
timestamp 1
transform -1 0 108836 0 1 105536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_1_Left_457
timestamp 1
transform 1 0 1104 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_1_Right_907
timestamp 1
transform -1 0 7912 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_2_Left_800
timestamp 1
transform 1 0 104052 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_191_2_Right_212
timestamp 1
transform -1 0 108836 0 -1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_1_Left_458
timestamp 1
transform 1 0 1104 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_1_Right_908
timestamp 1
transform -1 0 7912 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_2_Left_801
timestamp 1
transform 1 0 104052 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_192_2_Right_213
timestamp 1
transform -1 0 108836 0 1 106624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_1_Left_459
timestamp 1
transform 1 0 1104 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_1_Right_909
timestamp 1
transform -1 0 7912 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_2_Left_802
timestamp 1
transform 1 0 104052 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_193_2_Right_214
timestamp 1
transform -1 0 108836 0 -1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_1_Left_460
timestamp 1
transform 1 0 1104 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_1_Right_910
timestamp 1
transform -1 0 7912 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_2_Left_803
timestamp 1
transform 1 0 104052 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_194_2_Right_215
timestamp 1
transform -1 0 108836 0 1 107712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_1_Left_461
timestamp 1
transform 1 0 1104 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_1_Right_911
timestamp 1
transform -1 0 7912 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_2_Left_804
timestamp 1
transform 1 0 104052 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_195_2_Right_216
timestamp 1
transform -1 0 108836 0 -1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_1_Left_462
timestamp 1
transform 1 0 1104 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_1_Right_912
timestamp 1
transform -1 0 7912 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_2_Left_805
timestamp 1
transform 1 0 104052 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_196_2_Right_217
timestamp 1
transform -1 0 108836 0 1 108800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_1_Left_463
timestamp 1
transform 1 0 1104 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_1_Right_913
timestamp 1
transform -1 0 7912 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_2_Left_806
timestamp 1
transform 1 0 104052 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_197_2_Right_218
timestamp 1
transform -1 0 108836 0 -1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_1_Left_464
timestamp 1
transform 1 0 1104 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_1_Right_914
timestamp 1
transform -1 0 7912 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_2_Left_807
timestamp 1
transform 1 0 104052 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_198_2_Right_219
timestamp 1
transform -1 0 108836 0 1 109888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_1_Left_465
timestamp 1
transform 1 0 1104 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_1_Right_915
timestamp 1
transform -1 0 7912 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_2_Left_808
timestamp 1
transform 1 0 104052 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_199_2_Right_220
timestamp 1
transform -1 0 108836 0 -1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_1_Left_466
timestamp 1
transform 1 0 1104 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_1_Right_916
timestamp 1
transform -1 0 7912 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_2_Left_809
timestamp 1
transform 1 0 104052 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_200_2_Right_221
timestamp 1
transform -1 0 108836 0 1 110976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_1_Left_467
timestamp 1
transform 1 0 1104 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_1_Right_917
timestamp 1
transform -1 0 7912 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_2_Left_810
timestamp 1
transform 1 0 104052 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_201_2_Right_222
timestamp 1
transform -1 0 108836 0 -1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_1_Left_468
timestamp 1
transform 1 0 1104 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_1_Right_918
timestamp 1
transform -1 0 7912 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_2_Left_811
timestamp 1
transform 1 0 104052 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_202_2_Right_223
timestamp 1
transform -1 0 108836 0 1 112064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_1_Left_469
timestamp 1
transform 1 0 1104 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_1_Right_919
timestamp 1
transform -1 0 7912 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_2_Left_812
timestamp 1
transform 1 0 104052 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_203_2_Right_224
timestamp 1
transform -1 0 108836 0 -1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_1_Left_470
timestamp 1
transform 1 0 1104 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_1_Right_920
timestamp 1
transform -1 0 7912 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_2_Left_813
timestamp 1
transform 1 0 104052 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_204_2_Right_225
timestamp 1
transform -1 0 108836 0 1 113152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_1_Left_471
timestamp 1
transform 1 0 1104 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_1_Right_921
timestamp 1
transform -1 0 7912 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_2_Left_814
timestamp 1
transform 1 0 104052 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_205_2_Right_226
timestamp 1
transform -1 0 108836 0 -1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_1_Left_472
timestamp 1
transform 1 0 1104 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_1_Right_922
timestamp 1
transform -1 0 7912 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_2_Left_815
timestamp 1
transform 1 0 104052 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_206_2_Right_227
timestamp 1
transform -1 0 108836 0 1 114240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_1_Left_473
timestamp 1
transform 1 0 1104 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_1_Right_923
timestamp 1
transform -1 0 7912 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_2_Left_816
timestamp 1
transform 1 0 104052 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_207_2_Right_228
timestamp 1
transform -1 0 108836 0 -1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_1_Left_474
timestamp 1
transform 1 0 1104 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_1_Right_924
timestamp 1
transform -1 0 7912 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_2_Left_817
timestamp 1
transform 1 0 104052 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_208_2_Right_229
timestamp 1
transform -1 0 108836 0 1 115328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_1_Left_475
timestamp 1
transform 1 0 1104 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_1_Right_925
timestamp 1
transform -1 0 7912 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_2_Left_818
timestamp 1
transform 1 0 104052 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_209_2_Right_230
timestamp 1
transform -1 0 108836 0 -1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_1_Left_476
timestamp 1
transform 1 0 1104 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_1_Right_926
timestamp 1
transform -1 0 7912 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_2_Left_819
timestamp 1
transform 1 0 104052 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_210_2_Right_231
timestamp 1
transform -1 0 108836 0 1 116416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_1_Left_477
timestamp 1
transform 1 0 1104 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_1_Right_927
timestamp 1
transform -1 0 7912 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_2_Left_820
timestamp 1
transform 1 0 104052 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_211_2_Right_232
timestamp 1
transform -1 0 108836 0 -1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_1_Left_478
timestamp 1
transform 1 0 1104 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_1_Right_928
timestamp 1
transform -1 0 7912 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_2_Left_821
timestamp 1
transform 1 0 104052 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_212_2_Right_233
timestamp 1
transform -1 0 108836 0 1 117504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_1_Left_479
timestamp 1
transform 1 0 1104 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_1_Right_929
timestamp 1
transform -1 0 7912 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_2_Left_822
timestamp 1
transform 1 0 104052 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_213_2_Right_234
timestamp 1
transform -1 0 108836 0 -1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_1_Left_480
timestamp 1
transform 1 0 1104 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_1_Right_930
timestamp 1
transform -1 0 7912 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_2_Left_823
timestamp 1
transform 1 0 104052 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_214_2_Right_235
timestamp 1
transform -1 0 108836 0 1 118592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_1_Left_481
timestamp 1
transform 1 0 1104 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_1_Right_931
timestamp 1
transform -1 0 7912 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_2_Left_824
timestamp 1
transform 1 0 104052 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_215_2_Right_236
timestamp 1
transform -1 0 108836 0 -1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_1_Left_482
timestamp 1
transform 1 0 1104 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_1_Right_932
timestamp 1
transform -1 0 7912 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_2_Left_825
timestamp 1
transform 1 0 104052 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_216_2_Right_237
timestamp 1
transform -1 0 108836 0 1 119680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_1_Left_483
timestamp 1
transform 1 0 1104 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_1_Right_933
timestamp 1
transform -1 0 7912 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_2_Left_826
timestamp 1
transform 1 0 104052 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_217_2_Right_238
timestamp 1
transform -1 0 108836 0 -1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_1_Left_484
timestamp 1
transform 1 0 1104 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_1_Right_934
timestamp 1
transform -1 0 7912 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_2_Left_827
timestamp 1
transform 1 0 104052 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_218_2_Right_239
timestamp 1
transform -1 0 108836 0 1 120768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_1_Left_485
timestamp 1
transform 1 0 1104 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_1_Right_935
timestamp 1
transform -1 0 7912 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_2_Left_828
timestamp 1
transform 1 0 104052 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_219_2_Right_240
timestamp 1
transform -1 0 108836 0 -1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_1_Left_486
timestamp 1
transform 1 0 1104 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_1_Right_936
timestamp 1
transform -1 0 7912 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_2_Left_829
timestamp 1
transform 1 0 104052 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_220_2_Right_241
timestamp 1
transform -1 0 108836 0 1 121856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_1_Left_487
timestamp 1
transform 1 0 1104 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_1_Right_937
timestamp 1
transform -1 0 7912 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_2_Left_830
timestamp 1
transform 1 0 104052 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_221_2_Right_242
timestamp 1
transform -1 0 108836 0 -1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_1_Left_488
timestamp 1
transform 1 0 1104 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_1_Right_938
timestamp 1
transform -1 0 7912 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_2_Left_831
timestamp 1
transform 1 0 104052 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_222_2_Right_243
timestamp 1
transform -1 0 108836 0 1 122944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_1_Left_489
timestamp 1
transform 1 0 1104 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_1_Right_939
timestamp 1
transform -1 0 7912 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_2_Left_832
timestamp 1
transform 1 0 104052 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_223_2_Right_244
timestamp 1
transform -1 0 108836 0 -1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_1_Left_490
timestamp 1
transform 1 0 1104 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_1_Right_940
timestamp 1
transform -1 0 7912 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_2_Left_833
timestamp 1
transform 1 0 104052 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_224_2_Right_245
timestamp 1
transform -1 0 108836 0 1 124032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_1_Left_491
timestamp 1
transform 1 0 1104 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_1_Right_941
timestamp 1
transform -1 0 7912 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_2_Left_834
timestamp 1
transform 1 0 104052 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_225_2_Right_246
timestamp 1
transform -1 0 108836 0 -1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_1_Left_492
timestamp 1
transform 1 0 1104 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_1_Right_942
timestamp 1
transform -1 0 7912 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_2_Left_835
timestamp 1
transform 1 0 104052 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_226_2_Right_247
timestamp 1
transform -1 0 108836 0 1 125120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_1_Left_493
timestamp 1
transform 1 0 1104 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_1_Right_943
timestamp 1
transform -1 0 7912 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_2_Left_836
timestamp 1
transform 1 0 104052 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_227_2_Right_248
timestamp 1
transform -1 0 108836 0 -1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_1_Left_494
timestamp 1
transform 1 0 1104 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_1_Right_944
timestamp 1
transform -1 0 7912 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_2_Left_837
timestamp 1
transform 1 0 104052 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_228_2_Right_249
timestamp 1
transform -1 0 108836 0 1 126208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_1_Left_495
timestamp 1
transform 1 0 1104 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_1_Right_945
timestamp 1
transform -1 0 7912 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_2_Left_838
timestamp 1
transform 1 0 104052 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_229_2_Right_250
timestamp 1
transform -1 0 108836 0 -1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_230_1_Left_496
timestamp 1
transform 1 0 1104 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_230_1_Right_946
timestamp 1
transform -1 0 7912 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_230_2_Left_839
timestamp 1
transform 1 0 104052 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_230_2_Right_251
timestamp 1
transform -1 0 108836 0 1 127296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_231_1_Left_497
timestamp 1
transform 1 0 1104 0 -1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_231_1_Right_947
timestamp 1
transform -1 0 7912 0 -1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_231_2_Left_840
timestamp 1
transform 1 0 104052 0 -1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_231_2_Right_252
timestamp 1
transform -1 0 108836 0 -1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_232_1_Left_498
timestamp 1
transform 1 0 1104 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_232_1_Right_948
timestamp 1
transform -1 0 7912 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_232_2_Left_841
timestamp 1
transform 1 0 104052 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_232_2_Right_253
timestamp 1
transform -1 0 108836 0 1 128384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_233_1_Left_499
timestamp 1
transform 1 0 1104 0 -1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_233_1_Right_949
timestamp 1
transform -1 0 7912 0 -1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_233_2_Left_842
timestamp 1
transform 1 0 104052 0 -1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_233_2_Right_254
timestamp 1
transform -1 0 108836 0 -1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_234_1_Left_500
timestamp 1
transform 1 0 1104 0 1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_234_1_Right_950
timestamp 1
transform -1 0 7912 0 1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_234_2_Left_843
timestamp 1
transform 1 0 104052 0 1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_234_2_Right_255
timestamp 1
transform -1 0 108836 0 1 129472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_235_1_Left_501
timestamp 1
transform 1 0 1104 0 -1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_235_1_Right_951
timestamp 1
transform -1 0 7912 0 -1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_235_2_Left_844
timestamp 1
transform 1 0 104052 0 -1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_235_2_Right_256
timestamp 1
transform -1 0 108836 0 -1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_236_1_Left_502
timestamp 1
transform 1 0 1104 0 1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_236_1_Right_952
timestamp 1
transform -1 0 7912 0 1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_236_2_Left_845
timestamp 1
transform 1 0 104052 0 1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_236_2_Right_257
timestamp 1
transform -1 0 108836 0 1 130560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_237_1_Left_503
timestamp 1
transform 1 0 1104 0 -1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_237_1_Right_953
timestamp 1
transform -1 0 7912 0 -1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_237_2_Left_846
timestamp 1
transform 1 0 104052 0 -1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_237_2_Right_258
timestamp 1
transform -1 0 108836 0 -1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_238_1_Left_504
timestamp 1
transform 1 0 1104 0 1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_238_1_Right_954
timestamp 1
transform -1 0 7912 0 1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_238_2_Left_847
timestamp 1
transform 1 0 104052 0 1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_238_2_Right_259
timestamp 1
transform -1 0 108836 0 1 131648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_239_1_Left_505
timestamp 1
transform 1 0 1104 0 -1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_239_1_Right_955
timestamp 1
transform -1 0 7912 0 -1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_239_2_Left_848
timestamp 1
transform 1 0 104052 0 -1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_239_2_Right_260
timestamp 1
transform -1 0 108836 0 -1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_240_1_Left_506
timestamp 1
transform 1 0 1104 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_240_1_Right_956
timestamp 1
transform -1 0 7912 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_240_2_Left_849
timestamp 1
transform 1 0 104052 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_240_2_Right_261
timestamp 1
transform -1 0 108836 0 1 132736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_241_1_Left_507
timestamp 1
transform 1 0 1104 0 -1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_241_1_Right_957
timestamp 1
transform -1 0 7912 0 -1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_241_2_Left_850
timestamp 1
transform 1 0 104052 0 -1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_241_2_Right_262
timestamp 1
transform -1 0 108836 0 -1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_242_1_Left_508
timestamp 1
transform 1 0 1104 0 1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_242_1_Right_958
timestamp 1
transform -1 0 7912 0 1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_242_2_Left_851
timestamp 1
transform 1 0 104052 0 1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_242_2_Right_263
timestamp 1
transform -1 0 108836 0 1 133824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_243_1_Left_509
timestamp 1
transform 1 0 1104 0 -1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_243_1_Right_959
timestamp 1
transform -1 0 7912 0 -1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_243_2_Left_852
timestamp 1
transform 1 0 104052 0 -1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_243_2_Right_264
timestamp 1
transform -1 0 108836 0 -1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_244_1_Left_510
timestamp 1
transform 1 0 1104 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_244_1_Right_960
timestamp 1
transform -1 0 7912 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_244_2_Left_853
timestamp 1
transform 1 0 104052 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_244_2_Right_265
timestamp 1
transform -1 0 108836 0 1 134912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_245_1_Left_511
timestamp 1
transform 1 0 1104 0 -1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_245_1_Right_961
timestamp 1
transform -1 0 7912 0 -1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_245_2_Left_854
timestamp 1
transform 1 0 104052 0 -1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_245_2_Right_266
timestamp 1
transform -1 0 108836 0 -1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_246_Left_512
timestamp 1
transform 1 0 1104 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_246_Right_32
timestamp 1
transform -1 0 108836 0 1 136000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_247_Left_513
timestamp 1
transform 1 0 1104 0 -1 137088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_247_Right_33
timestamp 1
transform -1 0 108836 0 -1 137088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_248_Left_514
timestamp 1
transform 1 0 1104 0 1 137088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_248_Right_34
timestamp 1
transform -1 0 108836 0 1 137088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_249_Left_515
timestamp 1
transform 1 0 1104 0 -1 138176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_249_Right_35
timestamp 1
transform -1 0 108836 0 -1 138176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_250_Left_516
timestamp 1
transform 1 0 1104 0 1 138176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_250_Right_36
timestamp 1
transform -1 0 108836 0 1 138176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_251_Left_517
timestamp 1
transform 1 0 1104 0 -1 139264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_251_Right_37
timestamp 1
transform -1 0 108836 0 -1 139264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_252_Left_518
timestamp 1
transform 1 0 1104 0 1 139264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_252_Right_38
timestamp 1
transform -1 0 108836 0 1 139264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_253_Left_519
timestamp 1
transform 1 0 1104 0 -1 140352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_253_Right_39
timestamp 1
transform -1 0 108836 0 -1 140352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_254_Left_520
timestamp 1
transform 1 0 1104 0 1 140352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_254_Right_40
timestamp 1
transform -1 0 108836 0 1 140352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_255_Left_521
timestamp 1
transform 1 0 1104 0 -1 141440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_255_Right_41
timestamp 1
transform -1 0 108836 0 -1 141440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_256_Left_522
timestamp 1
transform 1 0 1104 0 1 141440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_256_Right_42
timestamp 1
transform -1 0 108836 0 1 141440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_257_Left_523
timestamp 1
transform 1 0 1104 0 -1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_257_Right_43
timestamp 1
transform -1 0 108836 0 -1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_258_Left_524
timestamp 1
transform 1 0 1104 0 1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_258_Right_44
timestamp 1
transform -1 0 108836 0 1 142528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_259_Left_525
timestamp 1
transform 1 0 1104 0 -1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_259_Right_45
timestamp 1
transform -1 0 108836 0 -1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_260_Left_526
timestamp 1
transform 1 0 1104 0 1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_260_Right_46
timestamp 1
transform -1 0 108836 0 1 143616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_261_Left_527
timestamp 1
transform 1 0 1104 0 -1 144704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_261_Right_47
timestamp 1
transform -1 0 108836 0 -1 144704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_262_Left_528
timestamp 1
transform 1 0 1104 0 1 144704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_262_Right_48
timestamp 1
transform -1 0 108836 0 1 144704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_263_Left_529
timestamp 1
transform 1 0 1104 0 -1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_263_Right_49
timestamp 1
transform -1 0 108836 0 -1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_264_Left_530
timestamp 1
transform 1 0 1104 0 1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_264_Right_50
timestamp 1
transform -1 0 108836 0 1 145792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_265_Left_531
timestamp 1
transform 1 0 1104 0 -1 146880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_265_Right_51
timestamp 1
transform -1 0 108836 0 -1 146880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_266_Left_532
timestamp 1
transform 1 0 1104 0 1 146880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_266_Right_52
timestamp 1
transform -1 0 108836 0 1 146880
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1
timestamp 1
transform -1 0 89516 0 -1 75072
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 1
transform 1 0 89976 0 1 77248
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp 1
transform 1 0 90620 0 1 77248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_962
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_963
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_964
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_965
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_966
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_967
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_968
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_969
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_970
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_971
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_972
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_973
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_974
timestamp 1
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_975
timestamp 1
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_976
timestamp 1
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_977
timestamp 1
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_978
timestamp 1
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_979
timestamp 1
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_980
timestamp 1
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_981
timestamp 1
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_982
timestamp 1
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_983
timestamp 1
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_984
timestamp 1
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_985
timestamp 1
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_986
timestamp 1
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_987
timestamp 1
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_988
timestamp 1
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_989
timestamp 1
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_990
timestamp 1
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_991
timestamp 1
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_992
timestamp 1
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_993
timestamp 1
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_994
timestamp 1
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_995
timestamp 1
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_996
timestamp 1
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_997
timestamp 1
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_998
timestamp 1
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_999
timestamp 1
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_1000
timestamp 1
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_1001
timestamp 1
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_1002
timestamp 1
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1003
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1004
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1005
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1006
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1007
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1008
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1009
timestamp 1
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1010
timestamp 1
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1011
timestamp 1
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1012
timestamp 1
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1013
timestamp 1
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1014
timestamp 1
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1015
timestamp 1
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1016
timestamp 1
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1017
timestamp 1
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1018
timestamp 1
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1019
timestamp 1
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1020
timestamp 1
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1021
timestamp 1
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_1022
timestamp 1
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1023
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1024
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1025
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1026
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1027
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1028
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1029
timestamp 1
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1030
timestamp 1
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1031
timestamp 1
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1032
timestamp 1
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1033
timestamp 1
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1034
timestamp 1
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1035
timestamp 1
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1036
timestamp 1
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1037
timestamp 1
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1038
timestamp 1
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1039
timestamp 1
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1040
timestamp 1
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1041
timestamp 1
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1042
timestamp 1
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_1043
timestamp 1
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1044
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1045
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1046
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1047
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1048
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1049
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1050
timestamp 1
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1051
timestamp 1
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1052
timestamp 1
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1053
timestamp 1
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1054
timestamp 1
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1055
timestamp 1
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1056
timestamp 1
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1057
timestamp 1
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1058
timestamp 1
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1059
timestamp 1
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1060
timestamp 1
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1061
timestamp 1
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1062
timestamp 1
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_1063
timestamp 1
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1064
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1065
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1066
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1067
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1068
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1069
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1070
timestamp 1
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1071
timestamp 1
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1072
timestamp 1
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1073
timestamp 1
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1074
timestamp 1
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1075
timestamp 1
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1076
timestamp 1
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1077
timestamp 1
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1078
timestamp 1
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1079
timestamp 1
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1080
timestamp 1
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1081
timestamp 1
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1082
timestamp 1
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1083
timestamp 1
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_1084
timestamp 1
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1085
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1086
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1087
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1088
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1089
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1090
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1091
timestamp 1
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1092
timestamp 1
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1093
timestamp 1
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1094
timestamp 1
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1095
timestamp 1
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1096
timestamp 1
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1097
timestamp 1
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1098
timestamp 1
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1099
timestamp 1
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1100
timestamp 1
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1101
timestamp 1
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1102
timestamp 1
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1103
timestamp 1
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1104
timestamp 1
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1105
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1106
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1107
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1108
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1109
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1110
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1111
timestamp 1
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1112
timestamp 1
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1113
timestamp 1
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1114
timestamp 1
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1115
timestamp 1
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1116
timestamp 1
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1117
timestamp 1
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1118
timestamp 1
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1119
timestamp 1
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1120
timestamp 1
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1121
timestamp 1
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1122
timestamp 1
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1123
timestamp 1
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1124
timestamp 1
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1125
timestamp 1
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1126
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1127
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1128
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1129
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1130
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1131
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1132
timestamp 1
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1133
timestamp 1
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1134
timestamp 1
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1135
timestamp 1
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1136
timestamp 1
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1137
timestamp 1
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1138
timestamp 1
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1139
timestamp 1
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1140
timestamp 1
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1141
timestamp 1
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1142
timestamp 1
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1143
timestamp 1
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1144
timestamp 1
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1145
timestamp 1
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1146
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1147
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1148
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1149
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1150
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1151
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1152
timestamp 1
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1153
timestamp 1
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1154
timestamp 1
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1155
timestamp 1
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1156
timestamp 1
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1157
timestamp 1
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1158
timestamp 1
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1159
timestamp 1
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1160
timestamp 1
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1161
timestamp 1
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1162
timestamp 1
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1163
timestamp 1
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1164
timestamp 1
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1165
timestamp 1
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1166
timestamp 1
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1167
timestamp 1
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1168
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1169
timestamp 1
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1170
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1171
timestamp 1
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1172
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1173
timestamp 1
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1174
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1175
timestamp 1
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1176
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1177
timestamp 1
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1178
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1179
timestamp 1
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1180
timestamp 1
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1181
timestamp 1
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1182
timestamp 1
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1183
timestamp 1
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1184
timestamp 1
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1185
timestamp 1
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1186
timestamp 1
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1187
timestamp 1
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1188
timestamp 1
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1189
timestamp 1
transform 1 0 60352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1190
timestamp 1
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1191
timestamp 1
transform 1 0 65504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1192
timestamp 1
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1193
timestamp 1
transform 1 0 70656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1194
timestamp 1
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1195
timestamp 1
transform 1 0 75808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1196
timestamp 1
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1197
timestamp 1
transform 1 0 80960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1198
timestamp 1
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1199
timestamp 1
transform 1 0 86112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1200
timestamp 1
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1201
timestamp 1
transform 1 0 91264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1202
timestamp 1
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1203
timestamp 1
transform 1 0 96416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1204
timestamp 1
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1205
timestamp 1
transform 1 0 101568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1206
timestamp 1
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1207
timestamp 1
transform 1 0 106720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_2384
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_2385
timestamp 1
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_1_1208
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_1209
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_2386
timestamp 1
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_1_1210
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_1211
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_2387
timestamp 1
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_1_1212
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_1213
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_2388
timestamp 1
transform 1 0 106628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_1_1214
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_1215
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_2389
timestamp 1
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_1_1216
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_1217
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_2390
timestamp 1
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_1_1218
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_1219
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_2391
timestamp 1
transform 1 0 106628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_1_1220
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_1221
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_2392
timestamp 1
transform 1 0 106628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_1_1222
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_1223
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_2393
timestamp 1
transform 1 0 106628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_1_1224
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_1225
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_2394
timestamp 1
transform 1 0 106628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_1_1226
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_1227
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_2395
timestamp 1
transform 1 0 106628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_1_1228
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_1229
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_2396
timestamp 1
transform 1 0 106628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_1_1230
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_1231
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_2397
timestamp 1
transform 1 0 106628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_1_1232
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_1233
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_2398
timestamp 1
transform 1 0 106628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_1_1234
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_1235
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_2399
timestamp 1
transform 1 0 106628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_1_1236
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_1237
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_2400
timestamp 1
transform 1 0 106628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_1_1238
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_1239
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_2401
timestamp 1
transform 1 0 106628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_1_1240
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_1241
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_2402
timestamp 1
transform 1 0 106628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_1_1242
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_1243
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_2403
timestamp 1
transform 1 0 106628 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_1_1244
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_1245
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_2404
timestamp 1
transform 1 0 106628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1_1246
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_1247
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_2405
timestamp 1
transform 1 0 106628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1_1248
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_1249
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_2406
timestamp 1
transform 1 0 106628 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1_1250
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_1251
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_2407
timestamp 1
transform 1 0 106628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1_1252
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_1253
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_2408
timestamp 1
transform 1 0 106628 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1_1254
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_1255
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_2409
timestamp 1
transform 1 0 106628 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1_1256
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_1257
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_2410
timestamp 1
transform 1 0 106628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1_1258
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_1259
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_2411
timestamp 1
transform 1 0 106628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1_1260
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_1261
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_2412
timestamp 1
transform 1 0 106628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1_1262
timestamp 1
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_1263
timestamp 1
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_2413
timestamp 1
transform 1 0 106628 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1_1264
timestamp 1
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_1265
timestamp 1
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_2414
timestamp 1
transform 1 0 106628 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1_1266
timestamp 1
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_1267
timestamp 1
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_2415
timestamp 1
transform 1 0 106628 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1_1268
timestamp 1
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_1269
timestamp 1
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_2416
timestamp 1
transform 1 0 106628 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1_1270
timestamp 1
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_1271
timestamp 1
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_2417
timestamp 1
transform 1 0 106628 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1_1272
timestamp 1
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_1273
timestamp 1
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_2418
timestamp 1
transform 1 0 106628 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1_1274
timestamp 1
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_1275
timestamp 1
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_2419
timestamp 1
transform 1 0 106628 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1_1276
timestamp 1
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_1277
timestamp 1
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_2420
timestamp 1
transform 1 0 106628 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1_1278
timestamp 1
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_1279
timestamp 1
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_2421
timestamp 1
transform 1 0 106628 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1_1280
timestamp 1
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_1281
timestamp 1
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_2422
timestamp 1
transform 1 0 106628 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1_1282
timestamp 1
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_1283
timestamp 1
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_2423
timestamp 1
transform 1 0 106628 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1_1284
timestamp 1
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_1285
timestamp 1
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_2424
timestamp 1
transform 1 0 106628 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1_1286
timestamp 1
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_1287
timestamp 1
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_2425
timestamp 1
transform 1 0 106628 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1_1288
timestamp 1
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_1289
timestamp 1
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_2426
timestamp 1
transform 1 0 106628 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1_1290
timestamp 1
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_1291
timestamp 1
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_2427
timestamp 1
transform 1 0 106628 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1_1292
timestamp 1
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_1293
timestamp 1
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_2428
timestamp 1
transform 1 0 106628 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1_1294
timestamp 1
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_1295
timestamp 1
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_2429
timestamp 1
transform 1 0 106628 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1_1296
timestamp 1
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_1297
timestamp 1
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_2430
timestamp 1
transform 1 0 106628 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1_1298
timestamp 1
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_1299
timestamp 1
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_2431
timestamp 1
transform 1 0 106628 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1_1300
timestamp 1
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_1301
timestamp 1
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_2432
timestamp 1
transform 1 0 106628 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1_1302
timestamp 1
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_1303
timestamp 1
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_2433
timestamp 1
transform 1 0 106628 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1_1304
timestamp 1
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_1305
timestamp 1
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_2434
timestamp 1
transform 1 0 106628 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1_1306
timestamp 1
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_1307
timestamp 1
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_2435
timestamp 1
transform 1 0 106628 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1_1308
timestamp 1
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_1309
timestamp 1
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_2436
timestamp 1
transform 1 0 106628 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1_1310
timestamp 1
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_1311
timestamp 1
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_2437
timestamp 1
transform 1 0 106628 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1_1312
timestamp 1
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_1313
timestamp 1
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_2438
timestamp 1
transform 1 0 106628 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1315
timestamp 1
transform 1 0 3680 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1316
timestamp 1
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1317
timestamp 1
transform 1 0 8832 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1318
timestamp 1
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1319
timestamp 1
transform 1 0 13984 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1320
timestamp 1
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1321
timestamp 1
transform 1 0 19136 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1322
timestamp 1
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1323
timestamp 1
transform 1 0 24288 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1324
timestamp 1
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1325
timestamp 1
transform 1 0 29440 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1326
timestamp 1
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1327
timestamp 1
transform 1 0 34592 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1328
timestamp 1
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1329
timestamp 1
transform 1 0 39744 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1330
timestamp 1
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1331
timestamp 1
transform 1 0 44896 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1332
timestamp 1
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1333
timestamp 1
transform 1 0 50048 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1334
timestamp 1
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1335
timestamp 1
transform 1 0 55200 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1336
timestamp 1
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1337
timestamp 1
transform 1 0 60352 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1338
timestamp 1
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1339
timestamp 1
transform 1 0 65504 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1340
timestamp 1
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1341
timestamp 1
transform 1 0 70656 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1342
timestamp 1
transform 1 0 73232 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1343
timestamp 1
transform 1 0 75808 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1344
timestamp 1
transform 1 0 78384 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1345
timestamp 1
transform 1 0 80960 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1346
timestamp 1
transform 1 0 83536 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1347
timestamp 1
transform 1 0 86112 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1348
timestamp 1
transform 1 0 88688 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1349
timestamp 1
transform 1 0 91264 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1350
timestamp 1
transform 1 0 93840 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1351
timestamp 1
transform 1 0 96416 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1352
timestamp 1
transform 1 0 98992 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1353
timestamp 1
transform 1 0 101568 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1354
timestamp 1
transform 1 0 104144 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1355
timestamp 1
transform 1 0 106720 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1356
timestamp 1
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1357
timestamp 1
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1358
timestamp 1
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1359
timestamp 1
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1360
timestamp 1
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1361
timestamp 1
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1362
timestamp 1
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1363
timestamp 1
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1364
timestamp 1
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1365
timestamp 1
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1366
timestamp 1
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1367
timestamp 1
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1368
timestamp 1
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1369
timestamp 1
transform 1 0 70656 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1370
timestamp 1
transform 1 0 75808 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1371
timestamp 1
transform 1 0 80960 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1372
timestamp 1
transform 1 0 86112 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1373
timestamp 1
transform 1 0 91264 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1374
timestamp 1
transform 1 0 96416 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1375
timestamp 1
transform 1 0 101568 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1376
timestamp 1
transform 1 0 106720 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1377
timestamp 1
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1378
timestamp 1
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1379
timestamp 1
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1380
timestamp 1
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1381
timestamp 1
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1382
timestamp 1
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1383
timestamp 1
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1384
timestamp 1
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1385
timestamp 1
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1386
timestamp 1
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1387
timestamp 1
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1388
timestamp 1
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1389
timestamp 1
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1390
timestamp 1
transform 1 0 73232 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1391
timestamp 1
transform 1 0 78384 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1392
timestamp 1
transform 1 0 83536 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1393
timestamp 1
transform 1 0 88688 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1394
timestamp 1
transform 1 0 93840 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1395
timestamp 1
transform 1 0 98992 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_1396
timestamp 1
transform 1 0 104144 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1397
timestamp 1
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1398
timestamp 1
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1399
timestamp 1
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1400
timestamp 1
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1401
timestamp 1
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1402
timestamp 1
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1403
timestamp 1
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1404
timestamp 1
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1405
timestamp 1
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1406
timestamp 1
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1407
timestamp 1
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1408
timestamp 1
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1409
timestamp 1
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1410
timestamp 1
transform 1 0 70656 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1411
timestamp 1
transform 1 0 75808 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1412
timestamp 1
transform 1 0 80960 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1413
timestamp 1
transform 1 0 86112 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1414
timestamp 1
transform 1 0 91264 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1415
timestamp 1
transform 1 0 96416 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1416
timestamp 1
transform 1 0 101568 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1417
timestamp 1
transform 1 0 106720 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1418
timestamp 1
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1419
timestamp 1
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1420
timestamp 1
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1421
timestamp 1
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1422
timestamp 1
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1423
timestamp 1
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1424
timestamp 1
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1425
timestamp 1
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1426
timestamp 1
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1427
timestamp 1
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1428
timestamp 1
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1429
timestamp 1
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1430
timestamp 1
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1431
timestamp 1
transform 1 0 73232 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1432
timestamp 1
transform 1 0 78384 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1433
timestamp 1
transform 1 0 83536 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1434
timestamp 1
transform 1 0 88688 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1435
timestamp 1
transform 1 0 93840 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1436
timestamp 1
transform 1 0 98992 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_1437
timestamp 1
transform 1 0 104144 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1438
timestamp 1
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1439
timestamp 1
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1440
timestamp 1
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1441
timestamp 1
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1442
timestamp 1
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1443
timestamp 1
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1444
timestamp 1
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1445
timestamp 1
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1446
timestamp 1
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1447
timestamp 1
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1448
timestamp 1
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1449
timestamp 1
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1450
timestamp 1
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1451
timestamp 1
transform 1 0 70656 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1452
timestamp 1
transform 1 0 75808 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1453
timestamp 1
transform 1 0 80960 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1454
timestamp 1
transform 1 0 86112 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1455
timestamp 1
transform 1 0 91264 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1456
timestamp 1
transform 1 0 96416 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1457
timestamp 1
transform 1 0 101568 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1458
timestamp 1
transform 1 0 106720 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1459
timestamp 1
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1460
timestamp 1
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1461
timestamp 1
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1462
timestamp 1
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1463
timestamp 1
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1464
timestamp 1
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1465
timestamp 1
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1466
timestamp 1
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1467
timestamp 1
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1468
timestamp 1
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1469
timestamp 1
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1470
timestamp 1
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1471
timestamp 1
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1472
timestamp 1
transform 1 0 73232 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1473
timestamp 1
transform 1 0 78384 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1474
timestamp 1
transform 1 0 83536 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1475
timestamp 1
transform 1 0 88688 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1476
timestamp 1
transform 1 0 93840 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1477
timestamp 1
transform 1 0 98992 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_1478
timestamp 1
transform 1 0 104144 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1479
timestamp 1
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1480
timestamp 1
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1481
timestamp 1
transform 1 0 13984 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1482
timestamp 1
transform 1 0 19136 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1483
timestamp 1
transform 1 0 24288 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1484
timestamp 1
transform 1 0 29440 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1485
timestamp 1
transform 1 0 34592 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1486
timestamp 1
transform 1 0 39744 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1487
timestamp 1
transform 1 0 44896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1488
timestamp 1
transform 1 0 50048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1489
timestamp 1
transform 1 0 55200 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1490
timestamp 1
transform 1 0 60352 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1491
timestamp 1
transform 1 0 65504 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1492
timestamp 1
transform 1 0 70656 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1493
timestamp 1
transform 1 0 75808 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1494
timestamp 1
transform 1 0 80960 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1495
timestamp 1
transform 1 0 86112 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1496
timestamp 1
transform 1 0 91264 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1497
timestamp 1
transform 1 0 96416 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1498
timestamp 1
transform 1 0 101568 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1499
timestamp 1
transform 1 0 106720 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1500
timestamp 1
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1501
timestamp 1
transform 1 0 11408 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1502
timestamp 1
transform 1 0 16560 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1503
timestamp 1
transform 1 0 21712 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1504
timestamp 1
transform 1 0 26864 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1505
timestamp 1
transform 1 0 32016 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1506
timestamp 1
transform 1 0 37168 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1507
timestamp 1
transform 1 0 42320 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1508
timestamp 1
transform 1 0 47472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1509
timestamp 1
transform 1 0 52624 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1510
timestamp 1
transform 1 0 57776 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1511
timestamp 1
transform 1 0 62928 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1512
timestamp 1
transform 1 0 68080 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1513
timestamp 1
transform 1 0 73232 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1514
timestamp 1
transform 1 0 78384 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1515
timestamp 1
transform 1 0 83536 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1516
timestamp 1
transform 1 0 88688 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1517
timestamp 1
transform 1 0 93840 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1518
timestamp 1
transform 1 0 98992 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1519
timestamp 1
transform 1 0 104144 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1520
timestamp 1
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1521
timestamp 1
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1522
timestamp 1
transform 1 0 13984 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1523
timestamp 1
transform 1 0 19136 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1524
timestamp 1
transform 1 0 24288 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1525
timestamp 1
transform 1 0 29440 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1526
timestamp 1
transform 1 0 34592 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1527
timestamp 1
transform 1 0 39744 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1528
timestamp 1
transform 1 0 44896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1529
timestamp 1
transform 1 0 50048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1530
timestamp 1
transform 1 0 55200 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1531
timestamp 1
transform 1 0 60352 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1532
timestamp 1
transform 1 0 65504 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1533
timestamp 1
transform 1 0 70656 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1534
timestamp 1
transform 1 0 75808 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1535
timestamp 1
transform 1 0 80960 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1536
timestamp 1
transform 1 0 86112 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1537
timestamp 1
transform 1 0 91264 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1538
timestamp 1
transform 1 0 96416 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1539
timestamp 1
transform 1 0 101568 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1540
timestamp 1
transform 1 0 106720 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1541
timestamp 1
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1542
timestamp 1
transform 1 0 11408 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1543
timestamp 1
transform 1 0 16560 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1544
timestamp 1
transform 1 0 21712 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1545
timestamp 1
transform 1 0 26864 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1546
timestamp 1
transform 1 0 32016 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1547
timestamp 1
transform 1 0 37168 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1548
timestamp 1
transform 1 0 42320 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1549
timestamp 1
transform 1 0 47472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1550
timestamp 1
transform 1 0 52624 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1551
timestamp 1
transform 1 0 57776 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1552
timestamp 1
transform 1 0 62928 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1553
timestamp 1
transform 1 0 68080 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1554
timestamp 1
transform 1 0 73232 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1555
timestamp 1
transform 1 0 78384 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1556
timestamp 1
transform 1 0 83536 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1557
timestamp 1
transform 1 0 88688 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1558
timestamp 1
transform 1 0 93840 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1559
timestamp 1
transform 1 0 98992 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1560
timestamp 1
transform 1 0 104144 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1561
timestamp 1
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1562
timestamp 1
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1563
timestamp 1
transform 1 0 13984 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1564
timestamp 1
transform 1 0 19136 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1565
timestamp 1
transform 1 0 24288 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1566
timestamp 1
transform 1 0 29440 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1567
timestamp 1
transform 1 0 34592 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1568
timestamp 1
transform 1 0 39744 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1569
timestamp 1
transform 1 0 44896 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1570
timestamp 1
transform 1 0 50048 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1571
timestamp 1
transform 1 0 55200 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1572
timestamp 1
transform 1 0 60352 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1573
timestamp 1
transform 1 0 65504 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1574
timestamp 1
transform 1 0 70656 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1575
timestamp 1
transform 1 0 75808 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1576
timestamp 1
transform 1 0 80960 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1577
timestamp 1
transform 1 0 86112 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1578
timestamp 1
transform 1 0 91264 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1579
timestamp 1
transform 1 0 96416 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1580
timestamp 1
transform 1 0 101568 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1581
timestamp 1
transform 1 0 106720 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1582
timestamp 1
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1583
timestamp 1
transform 1 0 11408 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1584
timestamp 1
transform 1 0 16560 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1585
timestamp 1
transform 1 0 21712 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1586
timestamp 1
transform 1 0 26864 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1587
timestamp 1
transform 1 0 32016 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1588
timestamp 1
transform 1 0 37168 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1589
timestamp 1
transform 1 0 42320 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1590
timestamp 1
transform 1 0 47472 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1591
timestamp 1
transform 1 0 52624 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1592
timestamp 1
transform 1 0 57776 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1593
timestamp 1
transform 1 0 62928 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1594
timestamp 1
transform 1 0 68080 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1595
timestamp 1
transform 1 0 73232 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1596
timestamp 1
transform 1 0 78384 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1597
timestamp 1
transform 1 0 83536 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1598
timestamp 1
transform 1 0 88688 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1599
timestamp 1
transform 1 0 93840 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1600
timestamp 1
transform 1 0 98992 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1601
timestamp 1
transform 1 0 104144 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1602
timestamp 1
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1603
timestamp 1
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1604
timestamp 1
transform 1 0 13984 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1605
timestamp 1
transform 1 0 19136 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1606
timestamp 1
transform 1 0 24288 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1607
timestamp 1
transform 1 0 29440 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1608
timestamp 1
transform 1 0 34592 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1609
timestamp 1
transform 1 0 39744 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1610
timestamp 1
transform 1 0 44896 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1611
timestamp 1
transform 1 0 50048 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1612
timestamp 1
transform 1 0 55200 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1613
timestamp 1
transform 1 0 60352 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1614
timestamp 1
transform 1 0 65504 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1615
timestamp 1
transform 1 0 70656 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1616
timestamp 1
transform 1 0 75808 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1617
timestamp 1
transform 1 0 80960 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1618
timestamp 1
transform 1 0 86112 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1619
timestamp 1
transform 1 0 91264 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1620
timestamp 1
transform 1 0 96416 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1621
timestamp 1
transform 1 0 101568 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1622
timestamp 1
transform 1 0 106720 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1623
timestamp 1
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1624
timestamp 1
transform 1 0 11408 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1625
timestamp 1
transform 1 0 16560 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1626
timestamp 1
transform 1 0 21712 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1627
timestamp 1
transform 1 0 26864 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1628
timestamp 1
transform 1 0 32016 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1629
timestamp 1
transform 1 0 37168 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1630
timestamp 1
transform 1 0 42320 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1631
timestamp 1
transform 1 0 47472 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1632
timestamp 1
transform 1 0 52624 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1633
timestamp 1
transform 1 0 57776 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1634
timestamp 1
transform 1 0 62928 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1635
timestamp 1
transform 1 0 68080 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1636
timestamp 1
transform 1 0 73232 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1637
timestamp 1
transform 1 0 78384 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1638
timestamp 1
transform 1 0 83536 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1639
timestamp 1
transform 1 0 88688 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1640
timestamp 1
transform 1 0 93840 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1641
timestamp 1
transform 1 0 98992 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1642
timestamp 1
transform 1 0 104144 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1643
timestamp 1
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1644
timestamp 1
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1645
timestamp 1
transform 1 0 13984 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1646
timestamp 1
transform 1 0 19136 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1647
timestamp 1
transform 1 0 24288 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1648
timestamp 1
transform 1 0 29440 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1649
timestamp 1
transform 1 0 34592 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1650
timestamp 1
transform 1 0 39744 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1651
timestamp 1
transform 1 0 44896 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1652
timestamp 1
transform 1 0 50048 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1653
timestamp 1
transform 1 0 55200 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1654
timestamp 1
transform 1 0 60352 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1655
timestamp 1
transform 1 0 65504 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1656
timestamp 1
transform 1 0 70656 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1657
timestamp 1
transform 1 0 75808 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1658
timestamp 1
transform 1 0 80960 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1659
timestamp 1
transform 1 0 86112 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1660
timestamp 1
transform 1 0 91264 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1661
timestamp 1
transform 1 0 96416 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1662
timestamp 1
transform 1 0 101568 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1663
timestamp 1
transform 1 0 106720 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1664
timestamp 1
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1665
timestamp 1
transform 1 0 11408 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1666
timestamp 1
transform 1 0 16560 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1667
timestamp 1
transform 1 0 21712 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1668
timestamp 1
transform 1 0 26864 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1669
timestamp 1
transform 1 0 32016 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1670
timestamp 1
transform 1 0 37168 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1671
timestamp 1
transform 1 0 42320 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1672
timestamp 1
transform 1 0 47472 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1673
timestamp 1
transform 1 0 52624 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1674
timestamp 1
transform 1 0 57776 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1675
timestamp 1
transform 1 0 62928 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1676
timestamp 1
transform 1 0 68080 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1677
timestamp 1
transform 1 0 73232 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1678
timestamp 1
transform 1 0 78384 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1679
timestamp 1
transform 1 0 83536 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1680
timestamp 1
transform 1 0 88688 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1681
timestamp 1
transform 1 0 93840 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1682
timestamp 1
transform 1 0 98992 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1683
timestamp 1
transform 1 0 104144 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1684
timestamp 1
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1685
timestamp 1
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1686
timestamp 1
transform 1 0 13984 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1687
timestamp 1
transform 1 0 19136 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1688
timestamp 1
transform 1 0 24288 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1689
timestamp 1
transform 1 0 29440 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1690
timestamp 1
transform 1 0 34592 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1691
timestamp 1
transform 1 0 39744 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1692
timestamp 1
transform 1 0 44896 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1693
timestamp 1
transform 1 0 50048 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1694
timestamp 1
transform 1 0 55200 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1695
timestamp 1
transform 1 0 60352 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1696
timestamp 1
transform 1 0 65504 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1697
timestamp 1
transform 1 0 70656 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1698
timestamp 1
transform 1 0 75808 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1699
timestamp 1
transform 1 0 80960 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1700
timestamp 1
transform 1 0 86112 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1701
timestamp 1
transform 1 0 91264 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1702
timestamp 1
transform 1 0 96416 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1703
timestamp 1
transform 1 0 101568 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1704
timestamp 1
transform 1 0 106720 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1705
timestamp 1
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1706
timestamp 1
transform 1 0 11408 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1707
timestamp 1
transform 1 0 16560 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1708
timestamp 1
transform 1 0 21712 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1709
timestamp 1
transform 1 0 26864 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1710
timestamp 1
transform 1 0 32016 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1711
timestamp 1
transform 1 0 37168 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1712
timestamp 1
transform 1 0 42320 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1713
timestamp 1
transform 1 0 47472 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1714
timestamp 1
transform 1 0 52624 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1715
timestamp 1
transform 1 0 57776 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1716
timestamp 1
transform 1 0 62928 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1717
timestamp 1
transform 1 0 68080 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1718
timestamp 1
transform 1 0 73232 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1719
timestamp 1
transform 1 0 78384 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1720
timestamp 1
transform 1 0 83536 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1721
timestamp 1
transform 1 0 88688 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1722
timestamp 1
transform 1 0 93840 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1723
timestamp 1
transform 1 0 98992 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1724
timestamp 1
transform 1 0 104144 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1725
timestamp 1
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1726
timestamp 1
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1727
timestamp 1
transform 1 0 13984 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1728
timestamp 1
transform 1 0 19136 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1729
timestamp 1
transform 1 0 24288 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1730
timestamp 1
transform 1 0 29440 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1731
timestamp 1
transform 1 0 34592 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1732
timestamp 1
transform 1 0 39744 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1733
timestamp 1
transform 1 0 44896 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1734
timestamp 1
transform 1 0 50048 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1735
timestamp 1
transform 1 0 55200 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1736
timestamp 1
transform 1 0 60352 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1737
timestamp 1
transform 1 0 65504 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1738
timestamp 1
transform 1 0 70656 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1739
timestamp 1
transform 1 0 75808 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1740
timestamp 1
transform 1 0 80960 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1741
timestamp 1
transform 1 0 86112 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1742
timestamp 1
transform 1 0 91264 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1743
timestamp 1
transform 1 0 96416 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1744
timestamp 1
transform 1 0 101568 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1745
timestamp 1
transform 1 0 106720 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1746
timestamp 1
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1747
timestamp 1
transform 1 0 11408 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1748
timestamp 1
transform 1 0 16560 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1749
timestamp 1
transform 1 0 21712 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1750
timestamp 1
transform 1 0 26864 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1751
timestamp 1
transform 1 0 32016 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1752
timestamp 1
transform 1 0 37168 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1753
timestamp 1
transform 1 0 42320 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1754
timestamp 1
transform 1 0 47472 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1755
timestamp 1
transform 1 0 52624 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1756
timestamp 1
transform 1 0 57776 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1757
timestamp 1
transform 1 0 62928 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1758
timestamp 1
transform 1 0 68080 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1759
timestamp 1
transform 1 0 73232 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1760
timestamp 1
transform 1 0 78384 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1761
timestamp 1
transform 1 0 83536 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1762
timestamp 1
transform 1 0 88688 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1763
timestamp 1
transform 1 0 93840 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1764
timestamp 1
transform 1 0 98992 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1765
timestamp 1
transform 1 0 104144 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1766
timestamp 1
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1767
timestamp 1
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1768
timestamp 1
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1769
timestamp 1
transform 1 0 11408 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1770
timestamp 1
transform 1 0 13984 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1771
timestamp 1
transform 1 0 16560 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1772
timestamp 1
transform 1 0 19136 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1773
timestamp 1
transform 1 0 21712 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1774
timestamp 1
transform 1 0 24288 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1775
timestamp 1
transform 1 0 26864 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1776
timestamp 1
transform 1 0 29440 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1777
timestamp 1
transform 1 0 32016 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1778
timestamp 1
transform 1 0 34592 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1779
timestamp 1
transform 1 0 37168 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1780
timestamp 1
transform 1 0 39744 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1781
timestamp 1
transform 1 0 42320 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1782
timestamp 1
transform 1 0 44896 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1783
timestamp 1
transform 1 0 47472 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1784
timestamp 1
transform 1 0 50048 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1785
timestamp 1
transform 1 0 52624 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1786
timestamp 1
transform 1 0 55200 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1787
timestamp 1
transform 1 0 57776 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1788
timestamp 1
transform 1 0 60352 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1789
timestamp 1
transform 1 0 62928 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1790
timestamp 1
transform 1 0 65504 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1791
timestamp 1
transform 1 0 68080 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1792
timestamp 1
transform 1 0 70656 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1793
timestamp 1
transform 1 0 73232 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1794
timestamp 1
transform 1 0 75808 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1795
timestamp 1
transform 1 0 78384 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1796
timestamp 1
transform 1 0 80960 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1797
timestamp 1
transform 1 0 83536 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1798
timestamp 1
transform 1 0 86112 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1799
timestamp 1
transform 1 0 88688 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1800
timestamp 1
transform 1 0 91264 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1801
timestamp 1
transform 1 0 93840 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1802
timestamp 1
transform 1 0 96416 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1803
timestamp 1
transform 1 0 98992 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1804
timestamp 1
transform 1 0 101568 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1805
timestamp 1
transform 1 0 104144 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1806
timestamp 1
transform 1 0 106720 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1_1314
timestamp 1
transform 1 0 6256 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_1807
timestamp 1
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_2439
timestamp 1
transform 1 0 106628 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1_1808
timestamp 1
transform 1 0 6256 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_1809
timestamp 1
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_2440
timestamp 1
transform 1 0 106628 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1_1810
timestamp 1
transform 1 0 6256 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_1811
timestamp 1
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_2441
timestamp 1
transform 1 0 106628 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1_1812
timestamp 1
transform 1 0 6256 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1_1813
timestamp 1
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_2442
timestamp 1
transform 1 0 106628 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1_1814
timestamp 1
transform 1 0 6256 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1_1815
timestamp 1
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_2443
timestamp 1
transform 1 0 106628 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1_1816
timestamp 1
transform 1 0 6256 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1_1817
timestamp 1
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_2444
timestamp 1
transform 1 0 106628 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1_1818
timestamp 1
transform 1 0 6256 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1_1819
timestamp 1
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_2445
timestamp 1
transform 1 0 106628 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1_1820
timestamp 1
transform 1 0 6256 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1_1821
timestamp 1
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_2446
timestamp 1
transform 1 0 106628 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1_1822
timestamp 1
transform 1 0 6256 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1_1823
timestamp 1
transform 1 0 3680 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_2_2447
timestamp 1
transform 1 0 106628 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1_1824
timestamp 1
transform 1 0 6256 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1_1825
timestamp 1
transform 1 0 3680 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_2_2448
timestamp 1
transform 1 0 106628 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1_1826
timestamp 1
transform 1 0 6256 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1_1827
timestamp 1
transform 1 0 3680 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_2_2449
timestamp 1
transform 1 0 106628 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1_1828
timestamp 1
transform 1 0 6256 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1_1829
timestamp 1
transform 1 0 3680 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_2_2450
timestamp 1
transform 1 0 106628 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1_1830
timestamp 1
transform 1 0 6256 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1_1831
timestamp 1
transform 1 0 3680 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_2_2451
timestamp 1
transform 1 0 106628 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1_1832
timestamp 1
transform 1 0 6256 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1_1833
timestamp 1
transform 1 0 3680 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_2_2452
timestamp 1
transform 1 0 106628 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1_1834
timestamp 1
transform 1 0 6256 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1_1835
timestamp 1
transform 1 0 3680 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_2_2453
timestamp 1
transform 1 0 106628 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1_1836
timestamp 1
transform 1 0 6256 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1_1837
timestamp 1
transform 1 0 3680 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_2_2454
timestamp 1
transform 1 0 106628 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1_1838
timestamp 1
transform 1 0 6256 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1_1839
timestamp 1
transform 1 0 3680 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_2_2455
timestamp 1
transform 1 0 106628 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1_1840
timestamp 1
transform 1 0 6256 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1_1841
timestamp 1
transform 1 0 3680 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_2_2456
timestamp 1
transform 1 0 106628 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1_1842
timestamp 1
transform 1 0 6256 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1_1843
timestamp 1
transform 1 0 3680 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_2_2457
timestamp 1
transform 1 0 106628 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1_1844
timestamp 1
transform 1 0 6256 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1_1845
timestamp 1
transform 1 0 3680 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_2_2458
timestamp 1
transform 1 0 106628 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1_1846
timestamp 1
transform 1 0 6256 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_1_1847
timestamp 1
transform 1 0 3680 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2_2459
timestamp 1
transform 1 0 106628 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_1_1848
timestamp 1
transform 1 0 6256 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_1_1849
timestamp 1
transform 1 0 3680 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2_2460
timestamp 1
transform 1 0 106628 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_183_1_1850
timestamp 1
transform 1 0 6256 0 -1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_184_1_1851
timestamp 1
transform 1 0 3680 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_184_2_2461
timestamp 1
transform 1 0 106628 0 1 102272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_185_1_1852
timestamp 1
transform 1 0 6256 0 -1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_186_1_1853
timestamp 1
transform 1 0 3680 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_186_2_2462
timestamp 1
transform 1 0 106628 0 1 103360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_187_1_1854
timestamp 1
transform 1 0 6256 0 -1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_188_1_1855
timestamp 1
transform 1 0 3680 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_188_2_2463
timestamp 1
transform 1 0 106628 0 1 104448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_189_1_1856
timestamp 1
transform 1 0 6256 0 -1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_190_1_1857
timestamp 1
transform 1 0 3680 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_190_2_2464
timestamp 1
transform 1 0 106628 0 1 105536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_191_1_1858
timestamp 1
transform 1 0 6256 0 -1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_192_1_1859
timestamp 1
transform 1 0 3680 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_192_2_2465
timestamp 1
transform 1 0 106628 0 1 106624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_193_1_1860
timestamp 1
transform 1 0 6256 0 -1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_194_1_1861
timestamp 1
transform 1 0 3680 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_194_2_2466
timestamp 1
transform 1 0 106628 0 1 107712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_195_1_1862
timestamp 1
transform 1 0 6256 0 -1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_196_1_1863
timestamp 1
transform 1 0 3680 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_196_2_2467
timestamp 1
transform 1 0 106628 0 1 108800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_197_1_1864
timestamp 1
transform 1 0 6256 0 -1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_198_1_1865
timestamp 1
transform 1 0 3680 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_198_2_2468
timestamp 1
transform 1 0 106628 0 1 109888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_199_1_1866
timestamp 1
transform 1 0 6256 0 -1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_200_1_1867
timestamp 1
transform 1 0 3680 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_200_2_2469
timestamp 1
transform 1 0 106628 0 1 110976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_201_1_1868
timestamp 1
transform 1 0 6256 0 -1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_202_1_1869
timestamp 1
transform 1 0 3680 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_202_2_2470
timestamp 1
transform 1 0 106628 0 1 112064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_203_1_1870
timestamp 1
transform 1 0 6256 0 -1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_204_1_1871
timestamp 1
transform 1 0 3680 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_204_2_2471
timestamp 1
transform 1 0 106628 0 1 113152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_205_1_1872
timestamp 1
transform 1 0 6256 0 -1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_206_1_1873
timestamp 1
transform 1 0 3680 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_206_2_2472
timestamp 1
transform 1 0 106628 0 1 114240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_207_1_1874
timestamp 1
transform 1 0 6256 0 -1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_208_1_1875
timestamp 1
transform 1 0 3680 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_208_2_2473
timestamp 1
transform 1 0 106628 0 1 115328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_209_1_1876
timestamp 1
transform 1 0 6256 0 -1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_210_1_1877
timestamp 1
transform 1 0 3680 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_210_2_2474
timestamp 1
transform 1 0 106628 0 1 116416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_211_1_1878
timestamp 1
transform 1 0 6256 0 -1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_212_1_1879
timestamp 1
transform 1 0 3680 0 1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_212_2_2475
timestamp 1
transform 1 0 106628 0 1 117504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_213_1_1880
timestamp 1
transform 1 0 6256 0 -1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_214_1_1881
timestamp 1
transform 1 0 3680 0 1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_214_2_2476
timestamp 1
transform 1 0 106628 0 1 118592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_215_1_1882
timestamp 1
transform 1 0 6256 0 -1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_216_1_1883
timestamp 1
transform 1 0 3680 0 1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_216_2_2477
timestamp 1
transform 1 0 106628 0 1 119680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_217_1_1884
timestamp 1
transform 1 0 6256 0 -1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_218_1_1885
timestamp 1
transform 1 0 3680 0 1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_218_2_2478
timestamp 1
transform 1 0 106628 0 1 120768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_219_1_1886
timestamp 1
transform 1 0 6256 0 -1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_220_1_1887
timestamp 1
transform 1 0 3680 0 1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_220_2_2479
timestamp 1
transform 1 0 106628 0 1 121856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_221_1_1888
timestamp 1
transform 1 0 6256 0 -1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_222_1_1889
timestamp 1
transform 1 0 3680 0 1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_222_2_2480
timestamp 1
transform 1 0 106628 0 1 122944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_223_1_1890
timestamp 1
transform 1 0 6256 0 -1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_224_1_1891
timestamp 1
transform 1 0 3680 0 1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_224_2_2481
timestamp 1
transform 1 0 106628 0 1 124032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_225_1_1892
timestamp 1
transform 1 0 6256 0 -1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_226_1_1893
timestamp 1
transform 1 0 3680 0 1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_226_2_2482
timestamp 1
transform 1 0 106628 0 1 125120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_227_1_1894
timestamp 1
transform 1 0 6256 0 -1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_1_1895
timestamp 1
transform 1 0 3680 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_228_2_2483
timestamp 1
transform 1 0 106628 0 1 126208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_229_1_1896
timestamp 1
transform 1 0 6256 0 -1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_230_1_1897
timestamp 1
transform 1 0 3680 0 1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_230_2_2484
timestamp 1
transform 1 0 106628 0 1 127296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_231_1_1898
timestamp 1
transform 1 0 6256 0 -1 128384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_232_1_1899
timestamp 1
transform 1 0 3680 0 1 128384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_232_2_2485
timestamp 1
transform 1 0 106628 0 1 128384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_233_1_1900
timestamp 1
transform 1 0 6256 0 -1 129472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_234_1_1901
timestamp 1
transform 1 0 3680 0 1 129472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_234_2_2486
timestamp 1
transform 1 0 106628 0 1 129472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_235_1_1902
timestamp 1
transform 1 0 6256 0 -1 130560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_236_1_1903
timestamp 1
transform 1 0 3680 0 1 130560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_236_2_2487
timestamp 1
transform 1 0 106628 0 1 130560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_237_1_1904
timestamp 1
transform 1 0 6256 0 -1 131648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_238_1_1905
timestamp 1
transform 1 0 3680 0 1 131648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_238_2_2488
timestamp 1
transform 1 0 106628 0 1 131648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_239_1_1906
timestamp 1
transform 1 0 6256 0 -1 132736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_240_1_1907
timestamp 1
transform 1 0 3680 0 1 132736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_240_2_2489
timestamp 1
transform 1 0 106628 0 1 132736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_241_1_1908
timestamp 1
transform 1 0 6256 0 -1 133824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_242_1_1909
timestamp 1
transform 1 0 3680 0 1 133824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_242_2_2490
timestamp 1
transform 1 0 106628 0 1 133824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_243_1_1910
timestamp 1
transform 1 0 6256 0 -1 134912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_244_1_1911
timestamp 1
transform 1 0 3680 0 1 134912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_244_2_2491
timestamp 1
transform 1 0 106628 0 1 134912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_245_1_1912
timestamp 1
transform 1 0 6256 0 -1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1913
timestamp 1
transform 1 0 3680 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1914
timestamp 1
transform 1 0 6256 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1915
timestamp 1
transform 1 0 8832 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1916
timestamp 1
transform 1 0 11408 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1917
timestamp 1
transform 1 0 13984 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1918
timestamp 1
transform 1 0 16560 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1919
timestamp 1
transform 1 0 19136 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1920
timestamp 1
transform 1 0 21712 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1921
timestamp 1
transform 1 0 24288 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1922
timestamp 1
transform 1 0 26864 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1923
timestamp 1
transform 1 0 29440 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1924
timestamp 1
transform 1 0 32016 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1925
timestamp 1
transform 1 0 34592 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1926
timestamp 1
transform 1 0 37168 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1927
timestamp 1
transform 1 0 39744 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1928
timestamp 1
transform 1 0 42320 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1929
timestamp 1
transform 1 0 44896 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1930
timestamp 1
transform 1 0 47472 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1931
timestamp 1
transform 1 0 50048 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1932
timestamp 1
transform 1 0 52624 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1933
timestamp 1
transform 1 0 55200 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1934
timestamp 1
transform 1 0 57776 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1935
timestamp 1
transform 1 0 60352 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1936
timestamp 1
transform 1 0 62928 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1937
timestamp 1
transform 1 0 65504 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1938
timestamp 1
transform 1 0 68080 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1939
timestamp 1
transform 1 0 70656 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1940
timestamp 1
transform 1 0 73232 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1941
timestamp 1
transform 1 0 75808 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1942
timestamp 1
transform 1 0 78384 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1943
timestamp 1
transform 1 0 80960 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1944
timestamp 1
transform 1 0 83536 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1945
timestamp 1
transform 1 0 86112 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1946
timestamp 1
transform 1 0 88688 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1947
timestamp 1
transform 1 0 91264 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1948
timestamp 1
transform 1 0 93840 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1949
timestamp 1
transform 1 0 96416 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1950
timestamp 1
transform 1 0 98992 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1951
timestamp 1
transform 1 0 101568 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1952
timestamp 1
transform 1 0 104144 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_246_1953
timestamp 1
transform 1 0 106720 0 1 136000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1954
timestamp 1
transform 1 0 6256 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1955
timestamp 1
transform 1 0 11408 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1956
timestamp 1
transform 1 0 16560 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1957
timestamp 1
transform 1 0 21712 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1958
timestamp 1
transform 1 0 26864 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1959
timestamp 1
transform 1 0 32016 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1960
timestamp 1
transform 1 0 37168 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1961
timestamp 1
transform 1 0 42320 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1962
timestamp 1
transform 1 0 47472 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1963
timestamp 1
transform 1 0 52624 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1964
timestamp 1
transform 1 0 57776 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1965
timestamp 1
transform 1 0 62928 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1966
timestamp 1
transform 1 0 68080 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1967
timestamp 1
transform 1 0 73232 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1968
timestamp 1
transform 1 0 78384 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1969
timestamp 1
transform 1 0 83536 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1970
timestamp 1
transform 1 0 88688 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1971
timestamp 1
transform 1 0 93840 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1972
timestamp 1
transform 1 0 98992 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_247_1973
timestamp 1
transform 1 0 104144 0 -1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1974
timestamp 1
transform 1 0 3680 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1975
timestamp 1
transform 1 0 8832 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1976
timestamp 1
transform 1 0 13984 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1977
timestamp 1
transform 1 0 19136 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1978
timestamp 1
transform 1 0 24288 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1979
timestamp 1
transform 1 0 29440 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1980
timestamp 1
transform 1 0 34592 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1981
timestamp 1
transform 1 0 39744 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1982
timestamp 1
transform 1 0 44896 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1983
timestamp 1
transform 1 0 50048 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1984
timestamp 1
transform 1 0 55200 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1985
timestamp 1
transform 1 0 60352 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1986
timestamp 1
transform 1 0 65504 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1987
timestamp 1
transform 1 0 70656 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1988
timestamp 1
transform 1 0 75808 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1989
timestamp 1
transform 1 0 80960 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1990
timestamp 1
transform 1 0 86112 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1991
timestamp 1
transform 1 0 91264 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1992
timestamp 1
transform 1 0 96416 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1993
timestamp 1
transform 1 0 101568 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_248_1994
timestamp 1
transform 1 0 106720 0 1 137088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1995
timestamp 1
transform 1 0 6256 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1996
timestamp 1
transform 1 0 11408 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1997
timestamp 1
transform 1 0 16560 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1998
timestamp 1
transform 1 0 21712 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_1999
timestamp 1
transform 1 0 26864 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2000
timestamp 1
transform 1 0 32016 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2001
timestamp 1
transform 1 0 37168 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2002
timestamp 1
transform 1 0 42320 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2003
timestamp 1
transform 1 0 47472 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2004
timestamp 1
transform 1 0 52624 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2005
timestamp 1
transform 1 0 57776 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2006
timestamp 1
transform 1 0 62928 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2007
timestamp 1
transform 1 0 68080 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2008
timestamp 1
transform 1 0 73232 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2009
timestamp 1
transform 1 0 78384 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2010
timestamp 1
transform 1 0 83536 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2011
timestamp 1
transform 1 0 88688 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2012
timestamp 1
transform 1 0 93840 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2013
timestamp 1
transform 1 0 98992 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_249_2014
timestamp 1
transform 1 0 104144 0 -1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2015
timestamp 1
transform 1 0 3680 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2016
timestamp 1
transform 1 0 8832 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2017
timestamp 1
transform 1 0 13984 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2018
timestamp 1
transform 1 0 19136 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2019
timestamp 1
transform 1 0 24288 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2020
timestamp 1
transform 1 0 29440 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2021
timestamp 1
transform 1 0 34592 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2022
timestamp 1
transform 1 0 39744 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2023
timestamp 1
transform 1 0 44896 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2024
timestamp 1
transform 1 0 50048 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2025
timestamp 1
transform 1 0 55200 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2026
timestamp 1
transform 1 0 60352 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2027
timestamp 1
transform 1 0 65504 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2028
timestamp 1
transform 1 0 70656 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2029
timestamp 1
transform 1 0 75808 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2030
timestamp 1
transform 1 0 80960 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2031
timestamp 1
transform 1 0 86112 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2032
timestamp 1
transform 1 0 91264 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2033
timestamp 1
transform 1 0 96416 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2034
timestamp 1
transform 1 0 101568 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_250_2035
timestamp 1
transform 1 0 106720 0 1 138176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2036
timestamp 1
transform 1 0 6256 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2037
timestamp 1
transform 1 0 11408 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2038
timestamp 1
transform 1 0 16560 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2039
timestamp 1
transform 1 0 21712 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2040
timestamp 1
transform 1 0 26864 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2041
timestamp 1
transform 1 0 32016 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2042
timestamp 1
transform 1 0 37168 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2043
timestamp 1
transform 1 0 42320 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2044
timestamp 1
transform 1 0 47472 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2045
timestamp 1
transform 1 0 52624 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2046
timestamp 1
transform 1 0 57776 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2047
timestamp 1
transform 1 0 62928 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2048
timestamp 1
transform 1 0 68080 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2049
timestamp 1
transform 1 0 73232 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2050
timestamp 1
transform 1 0 78384 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2051
timestamp 1
transform 1 0 83536 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2052
timestamp 1
transform 1 0 88688 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2053
timestamp 1
transform 1 0 93840 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2054
timestamp 1
transform 1 0 98992 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_251_2055
timestamp 1
transform 1 0 104144 0 -1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2056
timestamp 1
transform 1 0 3680 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2057
timestamp 1
transform 1 0 8832 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2058
timestamp 1
transform 1 0 13984 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2059
timestamp 1
transform 1 0 19136 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2060
timestamp 1
transform 1 0 24288 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2061
timestamp 1
transform 1 0 29440 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2062
timestamp 1
transform 1 0 34592 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2063
timestamp 1
transform 1 0 39744 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2064
timestamp 1
transform 1 0 44896 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2065
timestamp 1
transform 1 0 50048 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2066
timestamp 1
transform 1 0 55200 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2067
timestamp 1
transform 1 0 60352 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2068
timestamp 1
transform 1 0 65504 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2069
timestamp 1
transform 1 0 70656 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2070
timestamp 1
transform 1 0 75808 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2071
timestamp 1
transform 1 0 80960 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2072
timestamp 1
transform 1 0 86112 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2073
timestamp 1
transform 1 0 91264 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2074
timestamp 1
transform 1 0 96416 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2075
timestamp 1
transform 1 0 101568 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_252_2076
timestamp 1
transform 1 0 106720 0 1 139264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2077
timestamp 1
transform 1 0 6256 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2078
timestamp 1
transform 1 0 11408 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2079
timestamp 1
transform 1 0 16560 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2080
timestamp 1
transform 1 0 21712 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2081
timestamp 1
transform 1 0 26864 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2082
timestamp 1
transform 1 0 32016 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2083
timestamp 1
transform 1 0 37168 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2084
timestamp 1
transform 1 0 42320 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2085
timestamp 1
transform 1 0 47472 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2086
timestamp 1
transform 1 0 52624 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2087
timestamp 1
transform 1 0 57776 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2088
timestamp 1
transform 1 0 62928 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2089
timestamp 1
transform 1 0 68080 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2090
timestamp 1
transform 1 0 73232 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2091
timestamp 1
transform 1 0 78384 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2092
timestamp 1
transform 1 0 83536 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2093
timestamp 1
transform 1 0 88688 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2094
timestamp 1
transform 1 0 93840 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2095
timestamp 1
transform 1 0 98992 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_253_2096
timestamp 1
transform 1 0 104144 0 -1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2097
timestamp 1
transform 1 0 3680 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2098
timestamp 1
transform 1 0 8832 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2099
timestamp 1
transform 1 0 13984 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2100
timestamp 1
transform 1 0 19136 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2101
timestamp 1
transform 1 0 24288 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2102
timestamp 1
transform 1 0 29440 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2103
timestamp 1
transform 1 0 34592 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2104
timestamp 1
transform 1 0 39744 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2105
timestamp 1
transform 1 0 44896 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2106
timestamp 1
transform 1 0 50048 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2107
timestamp 1
transform 1 0 55200 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2108
timestamp 1
transform 1 0 60352 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2109
timestamp 1
transform 1 0 65504 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2110
timestamp 1
transform 1 0 70656 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2111
timestamp 1
transform 1 0 75808 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2112
timestamp 1
transform 1 0 80960 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2113
timestamp 1
transform 1 0 86112 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2114
timestamp 1
transform 1 0 91264 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2115
timestamp 1
transform 1 0 96416 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2116
timestamp 1
transform 1 0 101568 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_254_2117
timestamp 1
transform 1 0 106720 0 1 140352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2118
timestamp 1
transform 1 0 6256 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2119
timestamp 1
transform 1 0 11408 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2120
timestamp 1
transform 1 0 16560 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2121
timestamp 1
transform 1 0 21712 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2122
timestamp 1
transform 1 0 26864 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2123
timestamp 1
transform 1 0 32016 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2124
timestamp 1
transform 1 0 37168 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2125
timestamp 1
transform 1 0 42320 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2126
timestamp 1
transform 1 0 47472 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2127
timestamp 1
transform 1 0 52624 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2128
timestamp 1
transform 1 0 57776 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2129
timestamp 1
transform 1 0 62928 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2130
timestamp 1
transform 1 0 68080 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2131
timestamp 1
transform 1 0 73232 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2132
timestamp 1
transform 1 0 78384 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2133
timestamp 1
transform 1 0 83536 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2134
timestamp 1
transform 1 0 88688 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2135
timestamp 1
transform 1 0 93840 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2136
timestamp 1
transform 1 0 98992 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_255_2137
timestamp 1
transform 1 0 104144 0 -1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2138
timestamp 1
transform 1 0 3680 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2139
timestamp 1
transform 1 0 8832 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2140
timestamp 1
transform 1 0 13984 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2141
timestamp 1
transform 1 0 19136 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2142
timestamp 1
transform 1 0 24288 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2143
timestamp 1
transform 1 0 29440 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2144
timestamp 1
transform 1 0 34592 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2145
timestamp 1
transform 1 0 39744 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2146
timestamp 1
transform 1 0 44896 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2147
timestamp 1
transform 1 0 50048 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2148
timestamp 1
transform 1 0 55200 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2149
timestamp 1
transform 1 0 60352 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2150
timestamp 1
transform 1 0 65504 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2151
timestamp 1
transform 1 0 70656 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2152
timestamp 1
transform 1 0 75808 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2153
timestamp 1
transform 1 0 80960 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2154
timestamp 1
transform 1 0 86112 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2155
timestamp 1
transform 1 0 91264 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2156
timestamp 1
transform 1 0 96416 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2157
timestamp 1
transform 1 0 101568 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_256_2158
timestamp 1
transform 1 0 106720 0 1 141440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2159
timestamp 1
transform 1 0 6256 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2160
timestamp 1
transform 1 0 11408 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2161
timestamp 1
transform 1 0 16560 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2162
timestamp 1
transform 1 0 21712 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2163
timestamp 1
transform 1 0 26864 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2164
timestamp 1
transform 1 0 32016 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2165
timestamp 1
transform 1 0 37168 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2166
timestamp 1
transform 1 0 42320 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2167
timestamp 1
transform 1 0 47472 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2168
timestamp 1
transform 1 0 52624 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2169
timestamp 1
transform 1 0 57776 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2170
timestamp 1
transform 1 0 62928 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2171
timestamp 1
transform 1 0 68080 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2172
timestamp 1
transform 1 0 73232 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2173
timestamp 1
transform 1 0 78384 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2174
timestamp 1
transform 1 0 83536 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2175
timestamp 1
transform 1 0 88688 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2176
timestamp 1
transform 1 0 93840 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2177
timestamp 1
transform 1 0 98992 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_257_2178
timestamp 1
transform 1 0 104144 0 -1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2179
timestamp 1
transform 1 0 3680 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2180
timestamp 1
transform 1 0 8832 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2181
timestamp 1
transform 1 0 13984 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2182
timestamp 1
transform 1 0 19136 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2183
timestamp 1
transform 1 0 24288 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2184
timestamp 1
transform 1 0 29440 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2185
timestamp 1
transform 1 0 34592 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2186
timestamp 1
transform 1 0 39744 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2187
timestamp 1
transform 1 0 44896 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2188
timestamp 1
transform 1 0 50048 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2189
timestamp 1
transform 1 0 55200 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2190
timestamp 1
transform 1 0 60352 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2191
timestamp 1
transform 1 0 65504 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2192
timestamp 1
transform 1 0 70656 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2193
timestamp 1
transform 1 0 75808 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2194
timestamp 1
transform 1 0 80960 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2195
timestamp 1
transform 1 0 86112 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2196
timestamp 1
transform 1 0 91264 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2197
timestamp 1
transform 1 0 96416 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2198
timestamp 1
transform 1 0 101568 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_258_2199
timestamp 1
transform 1 0 106720 0 1 142528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2200
timestamp 1
transform 1 0 6256 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2201
timestamp 1
transform 1 0 11408 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2202
timestamp 1
transform 1 0 16560 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2203
timestamp 1
transform 1 0 21712 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2204
timestamp 1
transform 1 0 26864 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2205
timestamp 1
transform 1 0 32016 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2206
timestamp 1
transform 1 0 37168 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2207
timestamp 1
transform 1 0 42320 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2208
timestamp 1
transform 1 0 47472 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2209
timestamp 1
transform 1 0 52624 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2210
timestamp 1
transform 1 0 57776 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2211
timestamp 1
transform 1 0 62928 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2212
timestamp 1
transform 1 0 68080 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2213
timestamp 1
transform 1 0 73232 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2214
timestamp 1
transform 1 0 78384 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2215
timestamp 1
transform 1 0 83536 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2216
timestamp 1
transform 1 0 88688 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2217
timestamp 1
transform 1 0 93840 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2218
timestamp 1
transform 1 0 98992 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_259_2219
timestamp 1
transform 1 0 104144 0 -1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2220
timestamp 1
transform 1 0 3680 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2221
timestamp 1
transform 1 0 8832 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2222
timestamp 1
transform 1 0 13984 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2223
timestamp 1
transform 1 0 19136 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2224
timestamp 1
transform 1 0 24288 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2225
timestamp 1
transform 1 0 29440 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2226
timestamp 1
transform 1 0 34592 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2227
timestamp 1
transform 1 0 39744 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2228
timestamp 1
transform 1 0 44896 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2229
timestamp 1
transform 1 0 50048 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2230
timestamp 1
transform 1 0 55200 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2231
timestamp 1
transform 1 0 60352 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2232
timestamp 1
transform 1 0 65504 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2233
timestamp 1
transform 1 0 70656 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2234
timestamp 1
transform 1 0 75808 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2235
timestamp 1
transform 1 0 80960 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2236
timestamp 1
transform 1 0 86112 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2237
timestamp 1
transform 1 0 91264 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2238
timestamp 1
transform 1 0 96416 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2239
timestamp 1
transform 1 0 101568 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_260_2240
timestamp 1
transform 1 0 106720 0 1 143616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2241
timestamp 1
transform 1 0 6256 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2242
timestamp 1
transform 1 0 11408 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2243
timestamp 1
transform 1 0 16560 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2244
timestamp 1
transform 1 0 21712 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2245
timestamp 1
transform 1 0 26864 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2246
timestamp 1
transform 1 0 32016 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2247
timestamp 1
transform 1 0 37168 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2248
timestamp 1
transform 1 0 42320 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2249
timestamp 1
transform 1 0 47472 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2250
timestamp 1
transform 1 0 52624 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2251
timestamp 1
transform 1 0 57776 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2252
timestamp 1
transform 1 0 62928 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2253
timestamp 1
transform 1 0 68080 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2254
timestamp 1
transform 1 0 73232 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2255
timestamp 1
transform 1 0 78384 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2256
timestamp 1
transform 1 0 83536 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2257
timestamp 1
transform 1 0 88688 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2258
timestamp 1
transform 1 0 93840 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2259
timestamp 1
transform 1 0 98992 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_261_2260
timestamp 1
transform 1 0 104144 0 -1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2261
timestamp 1
transform 1 0 3680 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2262
timestamp 1
transform 1 0 8832 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2263
timestamp 1
transform 1 0 13984 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2264
timestamp 1
transform 1 0 19136 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2265
timestamp 1
transform 1 0 24288 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2266
timestamp 1
transform 1 0 29440 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2267
timestamp 1
transform 1 0 34592 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2268
timestamp 1
transform 1 0 39744 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2269
timestamp 1
transform 1 0 44896 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2270
timestamp 1
transform 1 0 50048 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2271
timestamp 1
transform 1 0 55200 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2272
timestamp 1
transform 1 0 60352 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2273
timestamp 1
transform 1 0 65504 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2274
timestamp 1
transform 1 0 70656 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2275
timestamp 1
transform 1 0 75808 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2276
timestamp 1
transform 1 0 80960 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2277
timestamp 1
transform 1 0 86112 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2278
timestamp 1
transform 1 0 91264 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2279
timestamp 1
transform 1 0 96416 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2280
timestamp 1
transform 1 0 101568 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_262_2281
timestamp 1
transform 1 0 106720 0 1 144704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2282
timestamp 1
transform 1 0 6256 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2283
timestamp 1
transform 1 0 11408 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2284
timestamp 1
transform 1 0 16560 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2285
timestamp 1
transform 1 0 21712 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2286
timestamp 1
transform 1 0 26864 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2287
timestamp 1
transform 1 0 32016 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2288
timestamp 1
transform 1 0 37168 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2289
timestamp 1
transform 1 0 42320 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2290
timestamp 1
transform 1 0 47472 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2291
timestamp 1
transform 1 0 52624 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2292
timestamp 1
transform 1 0 57776 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2293
timestamp 1
transform 1 0 62928 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2294
timestamp 1
transform 1 0 68080 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2295
timestamp 1
transform 1 0 73232 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2296
timestamp 1
transform 1 0 78384 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2297
timestamp 1
transform 1 0 83536 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2298
timestamp 1
transform 1 0 88688 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2299
timestamp 1
transform 1 0 93840 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2300
timestamp 1
transform 1 0 98992 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_263_2301
timestamp 1
transform 1 0 104144 0 -1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2302
timestamp 1
transform 1 0 3680 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2303
timestamp 1
transform 1 0 8832 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2304
timestamp 1
transform 1 0 13984 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2305
timestamp 1
transform 1 0 19136 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2306
timestamp 1
transform 1 0 24288 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2307
timestamp 1
transform 1 0 29440 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2308
timestamp 1
transform 1 0 34592 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2309
timestamp 1
transform 1 0 39744 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2310
timestamp 1
transform 1 0 44896 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2311
timestamp 1
transform 1 0 50048 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2312
timestamp 1
transform 1 0 55200 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2313
timestamp 1
transform 1 0 60352 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2314
timestamp 1
transform 1 0 65504 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2315
timestamp 1
transform 1 0 70656 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2316
timestamp 1
transform 1 0 75808 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2317
timestamp 1
transform 1 0 80960 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2318
timestamp 1
transform 1 0 86112 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2319
timestamp 1
transform 1 0 91264 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2320
timestamp 1
transform 1 0 96416 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2321
timestamp 1
transform 1 0 101568 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_264_2322
timestamp 1
transform 1 0 106720 0 1 145792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2323
timestamp 1
transform 1 0 6256 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2324
timestamp 1
transform 1 0 11408 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2325
timestamp 1
transform 1 0 16560 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2326
timestamp 1
transform 1 0 21712 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2327
timestamp 1
transform 1 0 26864 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2328
timestamp 1
transform 1 0 32016 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2329
timestamp 1
transform 1 0 37168 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2330
timestamp 1
transform 1 0 42320 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2331
timestamp 1
transform 1 0 47472 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2332
timestamp 1
transform 1 0 52624 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2333
timestamp 1
transform 1 0 57776 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2334
timestamp 1
transform 1 0 62928 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2335
timestamp 1
transform 1 0 68080 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2336
timestamp 1
transform 1 0 73232 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2337
timestamp 1
transform 1 0 78384 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2338
timestamp 1
transform 1 0 83536 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2339
timestamp 1
transform 1 0 88688 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2340
timestamp 1
transform 1 0 93840 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2341
timestamp 1
transform 1 0 98992 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_265_2342
timestamp 1
transform 1 0 104144 0 -1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2343
timestamp 1
transform 1 0 3680 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2344
timestamp 1
transform 1 0 6256 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2345
timestamp 1
transform 1 0 8832 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2346
timestamp 1
transform 1 0 11408 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2347
timestamp 1
transform 1 0 13984 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2348
timestamp 1
transform 1 0 16560 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2349
timestamp 1
transform 1 0 19136 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2350
timestamp 1
transform 1 0 21712 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2351
timestamp 1
transform 1 0 24288 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2352
timestamp 1
transform 1 0 26864 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2353
timestamp 1
transform 1 0 29440 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2354
timestamp 1
transform 1 0 32016 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2355
timestamp 1
transform 1 0 34592 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2356
timestamp 1
transform 1 0 37168 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2357
timestamp 1
transform 1 0 39744 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2358
timestamp 1
transform 1 0 42320 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2359
timestamp 1
transform 1 0 44896 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2360
timestamp 1
transform 1 0 47472 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2361
timestamp 1
transform 1 0 50048 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2362
timestamp 1
transform 1 0 52624 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2363
timestamp 1
transform 1 0 55200 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2364
timestamp 1
transform 1 0 57776 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2365
timestamp 1
transform 1 0 60352 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2366
timestamp 1
transform 1 0 62928 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2367
timestamp 1
transform 1 0 65504 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2368
timestamp 1
transform 1 0 68080 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2369
timestamp 1
transform 1 0 70656 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2370
timestamp 1
transform 1 0 73232 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2371
timestamp 1
transform 1 0 75808 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2372
timestamp 1
transform 1 0 78384 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2373
timestamp 1
transform 1 0 80960 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2374
timestamp 1
transform 1 0 83536 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2375
timestamp 1
transform 1 0 86112 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2376
timestamp 1
transform 1 0 88688 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2377
timestamp 1
transform 1 0 91264 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2378
timestamp 1
transform 1 0 93840 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2379
timestamp 1
transform 1 0 96416 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2380
timestamp 1
transform 1 0 98992 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2381
timestamp 1
transform 1 0 101568 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2382
timestamp 1
transform 1 0 104144 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_266_2383
timestamp 1
transform 1 0 106720 0 1 146880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire81
timestamp 1
transform 1 0 99728 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire83
timestamp 1
transform 1 0 100004 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  wire87
timestamp 1
transform 1 0 60444 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire88
timestamp 1
transform 1 0 57868 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire89
timestamp 1
transform 1 0 55292 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire90
timestamp 1
transform -1 0 50508 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire91
timestamp 1
transform -1 0 47932 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire92
timestamp 1
transform -1 0 43332 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire93
timestamp 1
transform -1 0 36340 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire94
timestamp 1
transform -1 0 35328 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire95
timestamp 1
transform 1 0 77280 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire96
timestamp 1
transform 1 0 73324 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire97
timestamp 1
transform 1 0 72404 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire98
timestamp 1
transform 1 0 63020 0 1 136000
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire99
timestamp 1
transform -1 0 34500 0 1 136000
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 addr00[0]
port 0 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 addr00[1]
port 1 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 addr00[2]
port 2 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 addr00[3]
port 3 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 addr00[4]
port 4 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 addr00[5]
port 5 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 addr00[6]
port 6 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 addr00[7]
port 7 nsew signal input
flabel metal3 s 0 71408 800 71528 0 FreeSans 480 0 0 0 addr01[0]
port 8 nsew signal input
flabel metal3 s 0 80248 800 80368 0 FreeSans 480 0 0 0 addr01[1]
port 9 nsew signal input
flabel metal3 s 0 104048 800 104168 0 FreeSans 480 0 0 0 addr01[2]
port 10 nsew signal input
flabel metal3 s 0 105408 800 105528 0 FreeSans 480 0 0 0 addr01[3]
port 11 nsew signal input
flabel metal3 s 0 106768 800 106888 0 FreeSans 480 0 0 0 addr01[4]
port 12 nsew signal input
flabel metal3 s 0 108128 800 108248 0 FreeSans 480 0 0 0 addr01[5]
port 13 nsew signal input
flabel metal3 s 0 109488 800 109608 0 FreeSans 480 0 0 0 addr01[6]
port 14 nsew signal input
flabel metal3 s 0 110848 800 110968 0 FreeSans 480 0 0 0 addr01[7]
port 15 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 csb00
port 17 nsew signal input
flabel metal3 s 0 85688 800 85808 0 FreeSans 480 0 0 0 csb01
port 18 nsew signal input
flabel metal3 s 109200 72088 110000 72208 0 FreeSans 480 0 0 0 denum[0]
port 19 nsew signal input
flabel metal3 s 109200 73448 110000 73568 0 FreeSans 480 0 0 0 denum[1]
port 20 nsew signal input
flabel metal3 s 109200 80248 110000 80368 0 FreeSans 480 0 0 0 denum[2]
port 21 nsew signal input
flabel metal3 s 109200 72768 110000 72888 0 FreeSans 480 0 0 0 denum[3]
port 22 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 din00[0]
port 23 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 din00[10]
port 24 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 din00[11]
port 25 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 din00[12]
port 26 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 din00[13]
port 27 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 din00[14]
port 28 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 din00[15]
port 29 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 din00[1]
port 30 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 din00[2]
port 31 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 din00[3]
port 32 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 din00[4]
port 33 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 din00[5]
port 34 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 din00[6]
port 35 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 din00[7]
port 36 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 din00[8]
port 37 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 din00[9]
port 38 nsew signal input
flabel metal3 s 0 77528 800 77648 0 FreeSans 480 0 0 0 din01[0]
port 39 nsew signal input
flabel metal3 s 0 79568 800 79688 0 FreeSans 480 0 0 0 din01[10]
port 40 nsew signal input
flabel metal3 s 0 81608 800 81728 0 FreeSans 480 0 0 0 din01[11]
port 41 nsew signal input
flabel metal3 s 0 82288 800 82408 0 FreeSans 480 0 0 0 din01[12]
port 42 nsew signal input
flabel metal3 s 0 82968 800 83088 0 FreeSans 480 0 0 0 din01[13]
port 43 nsew signal input
flabel metal3 s 0 78888 800 79008 0 FreeSans 480 0 0 0 din01[14]
port 44 nsew signal input
flabel metal3 s 0 83648 800 83768 0 FreeSans 480 0 0 0 din01[15]
port 45 nsew signal input
flabel metal3 s 0 84328 800 84448 0 FreeSans 480 0 0 0 din01[1]
port 46 nsew signal input
flabel metal3 s 0 85008 800 85128 0 FreeSans 480 0 0 0 din01[2]
port 47 nsew signal input
flabel metal3 s 0 78208 800 78328 0 FreeSans 480 0 0 0 din01[3]
port 48 nsew signal input
flabel metal3 s 0 86368 800 86488 0 FreeSans 480 0 0 0 din01[4]
port 49 nsew signal input
flabel metal3 s 0 87048 800 87168 0 FreeSans 480 0 0 0 din01[5]
port 50 nsew signal input
flabel metal3 s 0 80928 800 81048 0 FreeSans 480 0 0 0 din01[6]
port 51 nsew signal input
flabel metal3 s 0 87728 800 87848 0 FreeSans 480 0 0 0 din01[7]
port 52 nsew signal input
flabel metal3 s 0 76848 800 76968 0 FreeSans 480 0 0 0 din01[8]
port 53 nsew signal input
flabel metal3 s 0 88408 800 88528 0 FreeSans 480 0 0 0 din01[9]
port 54 nsew signal input
flabel metal3 s 109200 69368 110000 69488 0 FreeSans 480 0 0 0 num[0]
port 55 nsew signal input
flabel metal3 s 109200 70048 110000 70168 0 FreeSans 480 0 0 0 num[1]
port 56 nsew signal input
flabel metal3 s 109200 70728 110000 70848 0 FreeSans 480 0 0 0 num[2]
port 57 nsew signal input
flabel metal3 s 109200 71408 110000 71528 0 FreeSans 480 0 0 0 num[3]
port 58 nsew signal input
flabel metal3 s 109200 67328 110000 67448 0 FreeSans 480 0 0 0 rst
port 59 nsew signal input
flabel metal3 s 0 72088 800 72208 0 FreeSans 480 0 0 0 sine_out[0]
port 60 nsew signal output
flabel metal3 s 109200 76168 110000 76288 0 FreeSans 480 0 0 0 sine_out[10]
port 61 nsew signal output
flabel metal3 s 109200 79568 110000 79688 0 FreeSans 480 0 0 0 sine_out[11]
port 62 nsew signal output
flabel metal3 s 109200 78888 110000 79008 0 FreeSans 480 0 0 0 sine_out[12]
port 63 nsew signal output
flabel metal3 s 109200 77528 110000 77648 0 FreeSans 480 0 0 0 sine_out[13]
port 64 nsew signal output
flabel metal3 s 109200 76848 110000 76968 0 FreeSans 480 0 0 0 sine_out[14]
port 65 nsew signal output
flabel metal3 s 109200 78208 110000 78328 0 FreeSans 480 0 0 0 sine_out[15]
port 66 nsew signal output
flabel metal3 s 0 76168 800 76288 0 FreeSans 480 0 0 0 sine_out[1]
port 67 nsew signal output
flabel metal3 s 0 74808 800 74928 0 FreeSans 480 0 0 0 sine_out[2]
port 68 nsew signal output
flabel metal3 s 0 73448 800 73568 0 FreeSans 480 0 0 0 sine_out[3]
port 69 nsew signal output
flabel metal3 s 0 75488 800 75608 0 FreeSans 480 0 0 0 sine_out[4]
port 70 nsew signal output
flabel metal3 s 0 74128 800 74248 0 FreeSans 480 0 0 0 sine_out[5]
port 71 nsew signal output
flabel metal3 s 0 72768 800 72888 0 FreeSans 480 0 0 0 sine_out[6]
port 72 nsew signal output
flabel metal3 s 109200 74128 110000 74248 0 FreeSans 480 0 0 0 sine_out[7]
port 73 nsew signal output
flabel metal3 s 109200 74808 110000 74928 0 FreeSans 480 0 0 0 sine_out[8]
port 74 nsew signal output
flabel metal3 s 109200 75488 110000 75608 0 FreeSans 480 0 0 0 sine_out[9]
port 75 nsew signal output
flabel metal4 s 4208 2128 4528 147472 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 34928 2128 35248 7880 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 34928 65650 35248 77880 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 34928 135650 35248 147472 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 65648 2128 65968 8064 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 65648 65776 65968 78064 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 65648 135834 65968 147472 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 96368 2128 96688 8064 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 96368 65650 96688 78064 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 96368 135650 96688 147472 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 1056 5346 108884 5666 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 1056 35982 108884 36302 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 1056 66618 108884 66938 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 1056 97254 108884 97574 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 1056 127890 108884 128210 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 105916 7024 106236 66416 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 105916 77200 106236 136592 0 FreeSans 1920 90 0 0 vccd1
port 76 nsew power bidirectional
flabel metal5 s 4208 140940 108884 141260 0 FreeSans 2560 0 0 0 vccd1
port 76 nsew power bidirectional
flabel metal4 s 4868 2128 5188 147472 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 8064 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 35588 65650 35908 78064 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 35588 135650 35908 147472 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 66308 2128 66628 8064 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 66308 65650 66628 78064 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 66308 135650 66628 147472 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 97028 2128 97348 8064 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 97028 65650 97348 78064 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 97028 135650 97348 147472 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 1056 6006 108884 6326 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 1056 36642 108884 36962 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 1056 67278 108884 67598 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 1056 97914 108884 98234 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 1056 128550 108884 128870 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 106652 7024 106972 66416 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal4 s 106652 77200 106972 136592 0 FreeSans 1920 90 0 0 vssd1
port 77 nsew ground bidirectional
flabel metal5 s 4208 141620 108884 141940 0 FreeSans 2560 0 0 0 vssd1
port 77 nsew ground bidirectional
rlabel via4 101806 128050 101806 128050 0 vccd1
rlabel via4 101110 128710 101110 128710 0 vssd1
rlabel metal2 24702 73729 24702 73729 0 _000_
rlabel metal1 74934 73678 74934 73678 0 _001_
rlabel metal2 85882 76908 85882 76908 0 _002_
rlabel metal1 90666 75956 90666 75956 0 _003_
rlabel metal1 93518 77146 93518 77146 0 _004_
rlabel metal1 89930 77452 89930 77452 0 _005_
rlabel metal1 92874 77010 92874 77010 0 _006_
rlabel metal2 19366 76160 19366 76160 0 _007_
rlabel metal2 28566 75514 28566 75514 0 _008_
rlabel metal2 29394 73372 29394 73372 0 _009_
rlabel metal2 16238 77724 16238 77724 0 _010_
rlabel metal1 36432 72998 36432 72998 0 _011_
rlabel metal1 39882 73066 39882 73066 0 _012_
rlabel via1 74750 73797 74750 73797 0 _013_
rlabel metal2 78614 73508 78614 73508 0 _014_
rlabel metal2 73094 72896 73094 72896 0 _015_
rlabel metal2 87814 75038 87814 75038 0 _016_
rlabel metal2 89930 75446 89930 75446 0 _017_
rlabel metal1 90206 73576 90206 73576 0 _018_
rlabel metal1 91724 68850 91724 68850 0 _019_
rlabel metal2 91586 68952 91586 68952 0 _020_
rlabel metal1 89332 66538 89332 66538 0 _021_
rlabel metal1 89148 67762 89148 67762 0 _022_
rlabel metal1 88550 66198 88550 66198 0 _023_
rlabel metal1 87906 70618 87906 70618 0 _024_
rlabel metal2 23414 73984 23414 73984 0 _025_
rlabel metal2 22310 75786 22310 75786 0 _026_
rlabel metal2 19182 75072 19182 75072 0 _027_
rlabel metal1 22685 73066 22685 73066 0 _028_
rlabel metal1 15969 77418 15969 77418 0 _029_
rlabel metal1 22218 74263 22218 74263 0 _030_
rlabel metal1 27009 73814 27009 73814 0 _031_
rlabel metal1 85468 73882 85468 73882 0 _032_
rlabel metal2 85514 72488 85514 72488 0 _033_
rlabel metal1 88734 73134 88734 73134 0 _034_
rlabel metal1 87492 74154 87492 74154 0 _035_
rlabel metal1 92184 76058 92184 76058 0 _036_
rlabel metal1 92322 74426 92322 74426 0 _037_
rlabel metal1 96462 77690 96462 77690 0 _038_
rlabel metal1 94983 75990 94983 75990 0 _039_
rlabel metal2 96554 77350 96554 77350 0 _040_
rlabel metal2 85698 74664 85698 74664 0 _041_
rlabel metal2 89654 75106 89654 75106 0 _042_
rlabel metal2 90114 71808 90114 71808 0 _043_
rlabel metal1 90574 68646 90574 68646 0 _044_
rlabel metal1 89969 69462 89969 69462 0 _045_
rlabel metal2 86802 66810 86802 66810 0 _046_
rlabel metal2 86802 68204 86802 68204 0 _047_
rlabel metal1 85974 66538 85974 66538 0 _048_
rlabel metal1 86059 70890 86059 70890 0 _049_
rlabel metal1 103546 74868 103546 74868 0 _050_
rlabel metal1 103868 74834 103868 74834 0 _051_
rlabel metal2 106306 70924 106306 70924 0 _052_
rlabel metal2 100234 75344 100234 75344 0 _053_
rlabel metal2 101430 71842 101430 71842 0 _054_
rlabel metal2 104190 75412 104190 75412 0 _055_
rlabel metal1 101200 67218 101200 67218 0 _056_
rlabel metal1 104282 73712 104282 73712 0 _057_
rlabel metal1 103914 73100 103914 73100 0 _058_
rlabel metal1 103408 75242 103408 75242 0 _059_
rlabel metal1 103086 75514 103086 75514 0 _060_
rlabel metal1 103070 75242 103070 75242 0 _061_
rlabel metal1 102948 74290 102948 74290 0 _062_
rlabel metal2 103454 74086 103454 74086 0 _063_
rlabel metal1 104006 72590 104006 72590 0 _064_
rlabel metal1 103040 74222 103040 74222 0 _065_
rlabel metal2 103546 72794 103546 72794 0 _066_
rlabel metal1 104512 70414 104512 70414 0 _067_
rlabel metal1 104780 75174 104780 75174 0 _068_
rlabel metal2 105294 74698 105294 74698 0 _069_
rlabel metal2 104466 75038 104466 75038 0 _070_
rlabel metal1 104558 74698 104558 74698 0 _071_
rlabel metal1 105064 74834 105064 74834 0 _072_
rlabel metal1 104834 74222 104834 74222 0 _073_
rlabel metal1 104466 72658 104466 72658 0 _074_
rlabel metal2 103178 72250 103178 72250 0 _075_
rlabel metal2 103086 72250 103086 72250 0 _076_
rlabel metal2 102810 71740 102810 71740 0 _077_
rlabel metal1 103546 71536 103546 71536 0 _078_
rlabel metal1 105018 72794 105018 72794 0 _079_
rlabel metal2 105386 73270 105386 73270 0 _080_
rlabel metal1 105386 73882 105386 73882 0 _081_
rlabel metal2 105386 74460 105386 74460 0 _082_
rlabel metal1 104282 71536 104282 71536 0 _083_
rlabel metal1 103454 71604 103454 71604 0 _084_
rlabel metal1 103730 71502 103730 71502 0 _085_
rlabel metal1 105800 72046 105800 72046 0 _086_
rlabel metal1 106030 71978 106030 71978 0 _087_
rlabel metal1 105064 71366 105064 71366 0 _088_
rlabel metal2 105570 71468 105570 71468 0 _089_
rlabel metal2 105846 71536 105846 71536 0 _090_
rlabel metal1 105202 71026 105202 71026 0 _091_
rlabel metal1 105754 70550 105754 70550 0 _092_
rlabel metal1 104052 71026 104052 71026 0 _093_
rlabel metal1 103868 70482 103868 70482 0 _094_
rlabel metal1 102258 70924 102258 70924 0 _095_
rlabel metal1 95082 71434 95082 71434 0 _096_
rlabel metal1 103822 70822 103822 70822 0 _097_
rlabel metal2 103178 69836 103178 69836 0 _098_
rlabel metal1 102948 69394 102948 69394 0 _099_
rlabel metal2 106030 70822 106030 70822 0 _100_
rlabel metal1 105110 69802 105110 69802 0 _101_
rlabel metal1 103270 66640 103270 66640 0 _102_
rlabel metal2 103638 68986 103638 68986 0 _103_
rlabel metal2 103454 68986 103454 68986 0 _104_
rlabel metal1 104512 68442 104512 68442 0 _105_
rlabel metal1 105094 68714 105094 68714 0 _106_
rlabel metal1 103730 67286 103730 67286 0 _107_
rlabel metal1 104604 68782 104604 68782 0 _108_
rlabel metal1 105064 68986 105064 68986 0 _109_
rlabel metal2 104558 68714 104558 68714 0 _110_
rlabel metal1 104374 66130 104374 66130 0 _111_
rlabel metal1 102718 68442 102718 68442 0 _112_
rlabel metal1 103270 68646 103270 68646 0 _113_
rlabel metal1 101936 70958 101936 70958 0 _114_
rlabel metal1 102856 70890 102856 70890 0 _115_
rlabel metal1 98210 67354 98210 67354 0 _116_
rlabel metal1 96922 66164 96922 66164 0 _117_
rlabel metal1 103132 68986 103132 68986 0 _118_
rlabel metal1 101890 69428 101890 69428 0 _119_
rlabel metal1 103822 66130 103822 66130 0 _120_
rlabel metal1 104144 66266 104144 66266 0 _121_
rlabel metal1 104604 66606 104604 66606 0 _122_
rlabel metal2 103178 67184 103178 67184 0 _123_
rlabel metal2 103730 67456 103730 67456 0 _124_
rlabel metal2 102074 67830 102074 67830 0 _125_
rlabel metal2 102166 67745 102166 67745 0 _126_
rlabel metal1 101016 69734 101016 69734 0 _127_
rlabel metal1 102948 67354 102948 67354 0 _128_
rlabel metal2 102534 67932 102534 67932 0 _129_
rlabel metal1 101706 67252 101706 67252 0 _130_
rlabel metal1 101568 66130 101568 66130 0 _131_
rlabel metal2 101338 66334 101338 66334 0 _132_
rlabel metal1 102212 66674 102212 66674 0 _133_
rlabel metal1 101936 68442 101936 68442 0 _134_
rlabel metal1 100648 66130 100648 66130 0 _135_
rlabel metal1 100602 68170 100602 68170 0 _136_
rlabel metal1 102074 68170 102074 68170 0 _137_
rlabel metal1 101430 69802 101430 69802 0 _138_
rlabel metal1 101108 68782 101108 68782 0 _139_
rlabel metal2 98302 69190 98302 69190 0 _140_
rlabel metal1 100648 65926 100648 65926 0 _141_
rlabel metal2 99682 67388 99682 67388 0 _142_
rlabel metal1 100142 67320 100142 67320 0 _143_
rlabel metal1 100280 70074 100280 70074 0 _144_
rlabel metal2 101430 68612 101430 68612 0 _145_
rlabel metal1 101384 68442 101384 68442 0 _146_
rlabel metal1 98210 67728 98210 67728 0 _147_
rlabel metal1 99130 67898 99130 67898 0 _148_
rlabel metal1 97796 66606 97796 66606 0 _149_
rlabel metal2 98578 68034 98578 68034 0 _150_
rlabel metal2 99682 66368 99682 66368 0 _151_
rlabel metal1 99866 66810 99866 66810 0 _152_
rlabel metal1 100832 67014 100832 67014 0 _153_
rlabel metal2 102258 69292 102258 69292 0 _154_
rlabel metal1 101982 68850 101982 68850 0 _155_
rlabel metal1 100418 68272 100418 68272 0 _156_
rlabel metal1 99912 67286 99912 67286 0 _157_
rlabel metal1 98854 70958 98854 70958 0 _158_
rlabel metal2 99958 66266 99958 66266 0 _159_
rlabel metal1 99728 65994 99728 65994 0 _160_
rlabel metal1 100188 67898 100188 67898 0 _161_
rlabel metal1 100188 68442 100188 68442 0 _162_
rlabel metal1 100234 69904 100234 69904 0 _163_
rlabel metal1 98762 71604 98762 71604 0 _164_
rlabel metal1 97336 66266 97336 66266 0 _165_
rlabel metal2 97658 67524 97658 67524 0 _166_
rlabel metal1 98486 70992 98486 70992 0 _167_
rlabel metal1 97428 71570 97428 71570 0 _168_
rlabel metal1 97888 71638 97888 71638 0 _169_
rlabel metal1 99130 69836 99130 69836 0 _170_
rlabel metal1 98854 69360 98854 69360 0 _171_
rlabel metal1 98532 69326 98532 69326 0 _172_
rlabel metal1 97796 70482 97796 70482 0 _173_
rlabel metal1 97198 71094 97198 71094 0 _174_
rlabel metal1 98210 70414 98210 70414 0 _175_
rlabel metal1 99314 70448 99314 70448 0 _176_
rlabel metal1 96646 71162 96646 71162 0 _177_
rlabel metal1 98440 71570 98440 71570 0 _178_
rlabel metal1 97612 70414 97612 70414 0 _179_
rlabel metal1 97382 70448 97382 70448 0 _180_
rlabel metal1 97842 71536 97842 71536 0 _181_
rlabel metal1 99038 73338 99038 73338 0 _182_
rlabel metal1 98164 71706 98164 71706 0 _183_
rlabel metal1 97842 72624 97842 72624 0 _184_
rlabel metal2 99406 71264 99406 71264 0 _185_
rlabel metal1 99360 70074 99360 70074 0 _186_
rlabel metal2 99498 70788 99498 70788 0 _187_
rlabel metal2 100050 72318 100050 72318 0 _188_
rlabel metal1 98854 72726 98854 72726 0 _189_
rlabel metal1 101062 72794 101062 72794 0 _190_
rlabel metal2 98762 72386 98762 72386 0 _191_
rlabel metal1 98302 72794 98302 72794 0 _192_
rlabel metal1 96876 71706 96876 71706 0 _193_
rlabel metal1 97336 72046 97336 72046 0 _194_
rlabel metal1 98302 72012 98302 72012 0 _195_
rlabel metal1 98348 72658 98348 72658 0 _196_
rlabel metal2 100326 71332 100326 71332 0 _197_
rlabel metal1 100464 71706 100464 71706 0 _198_
rlabel metal1 100096 74834 100096 74834 0 _199_
rlabel metal2 100786 76534 100786 76534 0 _200_
rlabel metal2 100510 75004 100510 75004 0 _201_
rlabel metal1 101522 72250 101522 72250 0 _202_
rlabel metal1 101062 73168 101062 73168 0 _203_
rlabel metal1 101752 73066 101752 73066 0 _204_
rlabel metal1 102166 74902 102166 74902 0 _205_
rlabel metal1 101798 74800 101798 74800 0 _206_
rlabel metal2 101982 74630 101982 74630 0 _207_
rlabel metal2 101338 73372 101338 73372 0 _208_
rlabel metal2 101154 75616 101154 75616 0 _209_
rlabel metal1 100096 74970 100096 74970 0 _210_
rlabel metal2 101062 76636 101062 76636 0 _211_
rlabel metal1 97845 72794 97845 72794 0 _212_
rlabel via2 98578 73355 98578 73355 0 _213_
rlabel metal1 99222 73644 99222 73644 0 _214_
rlabel metal2 100326 74732 100326 74732 0 _215_
rlabel metal1 101154 75378 101154 75378 0 _216_
rlabel metal1 101430 75242 101430 75242 0 _217_
rlabel metal1 98578 75480 98578 75480 0 _218_
rlabel metal2 98486 76602 98486 76602 0 _219_
rlabel metal1 100142 74256 100142 74256 0 _220_
rlabel metal1 100510 73338 100510 73338 0 _221_
rlabel metal1 97106 75174 97106 75174 0 _222_
rlabel metal2 98670 76160 98670 76160 0 _223_
rlabel metal1 98026 74868 98026 74868 0 _224_
rlabel metal2 98578 75412 98578 75412 0 _225_
rlabel metal1 100556 76330 100556 76330 0 _226_
rlabel metal1 98762 76330 98762 76330 0 _227_
rlabel metal2 98762 76500 98762 76500 0 _228_
rlabel metal2 98302 75888 98302 75888 0 _229_
rlabel metal1 97060 75378 97060 75378 0 _230_
rlabel metal1 99774 74902 99774 74902 0 _231_
rlabel metal2 99222 73576 99222 73576 0 _232_
rlabel metal2 100418 74409 100418 74409 0 _233_
rlabel via1 97931 74222 97931 74222 0 _234_
rlabel metal2 96738 74596 96738 74596 0 _235_
rlabel metal1 97244 74970 97244 74970 0 _236_
rlabel metal1 97934 75174 97934 75174 0 _237_
rlabel metal2 98670 73916 98670 73916 0 _238_
rlabel metal2 97750 73610 97750 73610 0 _239_
rlabel metal2 97566 75276 97566 75276 0 _240_
rlabel metal2 98394 75514 98394 75514 0 _241_
rlabel metal2 97750 75140 97750 75140 0 _242_
rlabel metal1 96968 73134 96968 73134 0 _243_
rlabel metal1 94024 73746 94024 73746 0 _244_
rlabel metal2 96186 72318 96186 72318 0 _245_
rlabel metal2 95910 67932 95910 67932 0 _246_
rlabel metal1 96876 67014 96876 67014 0 _247_
rlabel metal2 95818 67218 95818 67218 0 _248_
rlabel metal1 95726 66062 95726 66062 0 _249_
rlabel metal2 94990 66844 94990 66844 0 _250_
rlabel metal2 96738 67150 96738 67150 0 _251_
rlabel metal2 95634 66436 95634 66436 0 _252_
rlabel metal1 94254 66130 94254 66130 0 _253_
rlabel metal2 94438 66878 94438 66878 0 _254_
rlabel metal2 96002 66368 96002 66368 0 _255_
rlabel metal2 95542 68000 95542 68000 0 _256_
rlabel metal1 95358 67354 95358 67354 0 _257_
rlabel metal1 95082 68850 95082 68850 0 _258_
rlabel metal2 95174 68374 95174 68374 0 _259_
rlabel metal1 96692 71434 96692 71434 0 _260_
rlabel metal1 95404 69938 95404 69938 0 _261_
rlabel metal2 94438 74188 94438 74188 0 _262_
rlabel via1 93592 72046 93592 72046 0 _263_
rlabel metal1 93426 72080 93426 72080 0 _264_
rlabel metal1 94576 71910 94576 71910 0 _265_
rlabel metal1 94898 68374 94898 68374 0 _266_
rlabel metal2 95358 67898 95358 67898 0 _267_
rlabel via1 96822 67354 96822 67354 0 _268_
rlabel metal2 96186 66844 96186 66844 0 _269_
rlabel metal1 96692 66606 96692 66606 0 _270_
rlabel metal1 95772 66810 95772 66810 0 _271_
rlabel metal1 89470 67660 89470 67660 0 _272_
rlabel metal2 90114 76534 90114 76534 0 _273_
rlabel metal1 90290 76058 90290 76058 0 _274_
rlabel metal1 90850 73576 90850 73576 0 _275_
rlabel metal1 90888 73814 90888 73814 0 _276_
rlabel metal1 93334 70822 93334 70822 0 _277_
rlabel metal1 92322 69190 92322 69190 0 _278_
rlabel metal1 92544 69530 92544 69530 0 _279_
rlabel metal2 93426 67728 93426 67728 0 _280_
rlabel metal2 92966 67898 92966 67898 0 _281_
rlabel metal2 91218 67014 91218 67014 0 _282_
rlabel metal2 89838 66912 89838 66912 0 _283_
rlabel metal1 91678 66232 91678 66232 0 _284_
rlabel metal1 90482 67286 90482 67286 0 _285_
rlabel metal2 90850 66980 90850 66980 0 _286_
rlabel metal1 90022 66198 90022 66198 0 _287_
rlabel metal1 89194 67898 89194 67898 0 _288_
rlabel metal1 89470 67354 89470 67354 0 _289_
rlabel metal1 88504 70482 88504 70482 0 _290_
rlabel metal1 1426 5202 1426 5202 0 addr00[0]
rlabel metal2 1978 8143 1978 8143 0 addr00[1]
rlabel metal1 1426 10642 1426 10642 0 addr00[2]
rlabel metal1 1380 11730 1380 11730 0 addr00[3]
rlabel metal2 1518 12563 1518 12563 0 addr00[4]
rlabel metal1 1426 13226 1426 13226 0 addr00[5]
rlabel metal2 1518 10999 1518 10999 0 addr00[6]
rlabel metal2 1518 13787 1518 13787 0 addr00[7]
rlabel metal1 1380 71570 1380 71570 0 addr01[0]
rlabel metal1 1380 80342 1380 80342 0 addr01[1]
rlabel metal1 1380 104210 1380 104210 0 addr01[2]
rlabel metal1 1380 105774 1380 105774 0 addr01[3]
rlabel metal1 1334 106862 1334 106862 0 addr01[4]
rlabel metal1 1380 108562 1380 108562 0 addr01[5]
rlabel metal1 1380 109650 1380 109650 0 addr01[6]
rlabel metal1 1380 111214 1380 111214 0 addr01[7]
rlabel metal1 55292 73746 55292 73746 0 clk
rlabel metal1 5244 82382 5244 82382 0 clknet_0_clk
rlabel metal1 82938 67626 82938 67626 0 clknet_2_0_0_clk
rlabel metal1 105248 91562 105248 91562 0 clknet_2_1_0_clk
rlabel metal1 5796 82246 5796 82246 0 clknet_2_2_0_clk
rlabel metal1 55246 77418 55246 77418 0 clknet_2_3_0_clk
rlabel metal1 63618 76398 63618 76398 0 clknet_3_0__leaf_clk
rlabel metal2 79534 70448 79534 70448 0 clknet_3_1__leaf_clk
rlabel metal1 91632 73542 91632 73542 0 clknet_3_2__leaf_clk
rlabel metal2 96002 136374 96002 136374 0 clknet_3_3__leaf_clk
rlabel metal4 16090 9798 16090 9798 0 clknet_3_4__leaf_clk
rlabel metal1 6624 94418 6624 94418 0 clknet_3_5__leaf_clk
rlabel metal1 37122 70006 37122 70006 0 clknet_3_6__leaf_clk
rlabel metal1 44482 76398 44482 76398 0 clknet_3_7__leaf_clk
rlabel metal2 1426 5593 1426 5593 0 csb00
rlabel metal1 1380 86190 1380 86190 0 csb01
rlabel metal2 108514 72403 108514 72403 0 denum[0]
rlabel metal2 108514 73627 108514 73627 0 denum[1]
rlabel via2 108514 80325 108514 80325 0 denum[2]
rlabel metal2 108514 72981 108514 72981 0 denum[3]
rlabel metal1 1380 6290 1380 6290 0 din00[0]
rlabel metal2 37398 1520 37398 1520 0 din00[10]
rlabel metal2 38686 1520 38686 1520 0 din00[11]
rlabel metal2 39974 1520 39974 1520 0 din00[12]
rlabel metal2 41262 1520 41262 1520 0 din00[13]
rlabel metal2 41906 1520 41906 1520 0 din00[14]
rlabel metal2 43194 1520 43194 1520 0 din00[15]
rlabel metal1 1380 8874 1380 8874 0 din00[1]
rlabel metal3 1004 6868 1004 6868 0 din00[2]
rlabel metal2 1518 9775 1518 9775 0 din00[3]
rlabel metal1 1426 7786 1426 7786 0 din00[4]
rlabel metal2 31602 1520 31602 1520 0 din00[5]
rlabel metal2 32890 1520 32890 1520 0 din00[6]
rlabel metal2 34178 1520 34178 1520 0 din00[7]
rlabel metal2 35466 1520 35466 1520 0 din00[8]
rlabel metal2 36110 1520 36110 1520 0 din00[9]
rlabel metal1 1426 78098 1426 78098 0 din01[0]
rlabel metal1 1380 79594 1380 79594 0 din01[10]
rlabel metal1 1380 81770 1380 81770 0 din01[11]
rlabel metal1 1380 82450 1380 82450 0 din01[12]
rlabel metal1 1426 83538 1426 83538 0 din01[13]
rlabel metal1 1426 79186 1426 79186 0 din01[14]
rlabel metal1 1380 84014 1380 84014 0 din01[15]
rlabel metal1 1426 84626 1426 84626 0 din01[1]
rlabel metal1 1380 85034 1380 85034 0 din01[2]
rlabel metal1 1426 78506 1426 78506 0 din01[3]
rlabel metal1 1426 86802 1426 86802 0 din01[4]
rlabel metal1 1380 87210 1380 87210 0 din01[5]
rlabel metal1 1426 81362 1426 81362 0 din01[6]
rlabel metal1 1380 87890 1380 87890 0 din01[7]
rlabel metal1 1380 77010 1380 77010 0 din01[8]
rlabel metal1 1426 88978 1426 88978 0 din01[9]
rlabel metal1 1794 5066 1794 5066 0 net1
rlabel metal1 4002 80614 4002 80614 0 net10
rlabel metal2 68310 73440 68310 73440 0 net100
rlabel metal1 74934 74426 74934 74426 0 net101
rlabel metal4 87342 63983 87342 63983 0 net102
rlabel metal1 86940 67354 86940 67354 0 net103
rlabel metal1 85100 66606 85100 66606 0 net104
rlabel metal2 36202 72726 36202 72726 0 net105
rlabel metal1 97980 71570 97980 71570 0 net106
rlabel metal1 101062 67286 101062 67286 0 net107
rlabel metal1 103132 73134 103132 73134 0 net108
rlabel metal1 98762 74868 98762 74868 0 net109
rlabel metal2 9522 104003 9522 104003 0 net11
rlabel metal1 99038 67762 99038 67762 0 net110
rlabel metal1 105386 72998 105386 72998 0 net111
rlabel metal2 105662 73066 105662 73066 0 net112
rlabel metal2 101154 68476 101154 68476 0 net113
rlabel metal3 102279 59738 102279 59738 0 net114
rlabel metal3 102279 129738 102279 129738 0 net115
rlabel metal4 86174 63983 86174 63983 0 net116
rlabel metal1 90666 77588 90666 77588 0 net117
rlabel metal2 86342 135762 86342 135762 0 net118
rlabel metal2 9522 105761 9522 105761 0 net12
rlabel metal2 9522 106847 9522 106847 0 net13
rlabel via2 9522 108411 9522 108411 0 net14
rlabel via2 9522 109519 9522 109519 0 net15
rlabel metal2 9522 111287 9522 111287 0 net16
rlabel metal1 1702 5882 1702 5882 0 net17
rlabel metal2 5566 85765 5566 85765 0 net18
rlabel metal1 108054 71570 108054 71570 0 net19
rlabel metal1 1978 8364 1978 8364 0 net2
rlabel metal1 105662 73848 105662 73848 0 net20
rlabel metal1 108008 80750 108008 80750 0 net21
rlabel metal1 106306 73100 106306 73100 0 net22
rlabel metal1 1794 6154 1794 6154 0 net23
rlabel metal4 37486 9934 37486 9934 0 net24
rlabel metal4 38654 9934 38654 9934 0 net25
rlabel metal1 40020 2618 40020 2618 0 net26
rlabel metal4 40990 9934 40990 9934 0 net27
rlabel metal4 42158 9934 42158 9934 0 net28
rlabel metal3 43401 8228 43401 8228 0 net29
rlabel metal1 1702 10778 1702 10778 0 net3
rlabel metal1 1794 8874 1794 8874 0 net30
rlabel metal1 1794 7242 1794 7242 0 net31
rlabel metal1 1794 9962 1794 9962 0 net32
rlabel metal1 1794 7786 1794 7786 0 net33
rlabel via3 31717 8228 31717 8228 0 net34
rlabel metal4 32814 9866 32814 9866 0 net35
rlabel metal4 33982 9866 33982 9866 0 net36
rlabel metal1 35512 2618 35512 2618 0 net37
rlabel metal4 36318 9934 36318 9934 0 net38
rlabel metal1 1794 77962 1794 77962 0 net39
rlabel metal1 1702 11866 1702 11866 0 net4
rlabel metal1 1794 79594 1794 79594 0 net40
rlabel metal2 1886 81260 1886 81260 0 net41
rlabel metal1 2300 82246 2300 82246 0 net42
rlabel metal1 1978 83334 1978 83334 0 net43
rlabel metal1 1794 79050 1794 79050 0 net44
rlabel metal1 2208 83878 2208 83878 0 net45
rlabel metal1 1748 84490 1748 84490 0 net46
rlabel metal1 1978 84966 1978 84966 0 net47
rlabel metal1 1794 78506 1794 78506 0 net48
rlabel metal1 1794 86666 1794 86666 0 net49
rlabel metal1 1748 12954 1748 12954 0 net5
rlabel metal2 1886 86360 1886 86360 0 net50
rlabel metal1 1794 81226 1794 81226 0 net51
rlabel metal1 1794 87754 1794 87754 0 net52
rlabel metal1 1978 77146 1978 77146 0 net53
rlabel metal1 1794 88842 1794 88842 0 net54
rlabel metal1 105708 71570 105708 71570 0 net55
rlabel metal1 108238 70618 108238 70618 0 net56
rlabel metal1 107824 71162 107824 71162 0 net57
rlabel metal2 104558 71876 104558 71876 0 net58
rlabel metal1 91356 70482 91356 70482 0 net59
rlabel metal1 1978 13498 1978 13498 0 net6
rlabel metal1 1794 72658 1794 72658 0 net60
rlabel metal1 94484 74358 94484 74358 0 net61
rlabel metal1 96278 76602 96278 76602 0 net62
rlabel metal1 95864 75514 95864 75514 0 net63
rlabel metal2 108238 77860 108238 77860 0 net64
rlabel metal2 100602 76500 100602 76500 0 net65
rlabel metal2 107686 77724 107686 77724 0 net66
rlabel metal1 14720 75854 14720 75854 0 net67
rlabel metal2 18170 75038 18170 75038 0 net68
rlabel metal2 1886 73440 1886 73440 0 net69
rlabel metal1 1748 11322 1748 11322 0 net7
rlabel metal2 11086 76772 11086 76772 0 net70
rlabel metal1 1794 74222 1794 74222 0 net71
rlabel metal1 1794 73134 1794 73134 0 net72
rlabel metal1 90022 74120 90022 74120 0 net73
rlabel metal2 94530 72488 94530 72488 0 net74
rlabel metal1 92460 73814 92460 73814 0 net75
rlabel metal1 99590 74732 99590 74732 0 net76
rlabel metal2 102074 74596 102074 74596 0 net77
rlabel metal1 96140 69734 96140 69734 0 net78
rlabel metal2 97106 70550 97106 70550 0 net79
rlabel metal1 2668 14042 2668 14042 0 net8
rlabel metal1 96922 70958 96922 70958 0 net80
rlabel metal1 99636 68646 99636 68646 0 net81
rlabel metal2 99682 69564 99682 69564 0 net82
rlabel metal2 99774 70074 99774 70074 0 net83
rlabel metal1 97934 68782 97934 68782 0 net84
rlabel metal1 105248 71978 105248 71978 0 net85
rlabel metal1 105800 71502 105800 71502 0 net86
rlabel metal2 60950 135932 60950 135932 0 net87
rlabel via1 63153 76330 63153 76330 0 net88
rlabel via1 61037 76330 61037 76330 0 net89
rlabel metal1 1794 71434 1794 71434 0 net9
rlabel metal2 46966 76874 46966 76874 0 net90
rlabel metal1 44210 76330 44210 76330 0 net91
rlabel metal2 43102 135966 43102 135966 0 net92
rlabel metal1 36248 136102 36248 136102 0 net93
rlabel metal1 8326 101082 8326 101082 0 net94
rlabel metal2 77786 135796 77786 135796 0 net95
rlabel metal2 73830 135830 73830 135830 0 net96
rlabel metal2 72910 135864 72910 135864 0 net97
rlabel metal2 63526 135898 63526 135898 0 net98
rlabel metal2 34178 135388 34178 135388 0 net99
rlabel metal2 108514 69649 108514 69649 0 num[0]
rlabel metal1 108376 70482 108376 70482 0 num[1]
rlabel metal2 108514 70873 108514 70873 0 num[2]
rlabel metal2 108514 71519 108514 71519 0 num[3]
rlabel metal2 108514 67541 108514 67541 0 rst
rlabel metal3 751 72148 751 72148 0 sine_out[0]
rlabel via2 108422 76245 108422 76245 0 sine_out[10]
rlabel metal2 108422 79577 108422 79577 0 sine_out[11]
rlabel via2 108422 78965 108422 78965 0 sine_out[12]
rlabel metal2 108422 77741 108422 77741 0 sine_out[13]
rlabel via2 108422 76891 108422 76891 0 sine_out[14]
rlabel metal2 108422 78353 108422 78353 0 sine_out[15]
rlabel metal3 751 76228 751 76228 0 sine_out[1]
rlabel metal3 751 74868 751 74868 0 sine_out[2]
rlabel metal3 751 73508 751 73508 0 sine_out[3]
rlabel metal3 1096 75548 1096 75548 0 sine_out[4]
rlabel metal3 751 74188 751 74188 0 sine_out[5]
rlabel metal3 751 72828 751 72828 0 sine_out[6]
rlabel metal2 108422 74137 108422 74137 0 sine_out[7]
rlabel metal2 108422 75021 108422 75021 0 sine_out[8]
rlabel metal2 108422 75803 108422 75803 0 sine_out[9]
rlabel metal1 31947 70618 31947 70618 0 sine_out_reg0\[0\]
rlabel metal2 74566 71468 74566 71468 0 sine_out_reg0\[10\]
rlabel metal2 84042 74256 84042 74256 0 sine_out_reg0\[11\]
rlabel metal1 77832 70074 77832 70074 0 sine_out_reg0\[12\]
rlabel metal1 90666 76976 90666 76976 0 sine_out_reg0\[13\]
rlabel metal1 79718 69836 79718 69836 0 sine_out_reg0\[14\]
rlabel metal1 84640 70006 84640 70006 0 sine_out_reg0\[15\]
rlabel metal2 30590 73338 30590 73338 0 sine_out_reg0\[1\]
rlabel metal2 34546 70720 34546 70720 0 sine_out_reg0\[2\]
rlabel metal1 37168 73746 37168 73746 0 sine_out_reg0\[3\]
rlabel metal1 34362 70006 34362 70006 0 sine_out_reg0\[4\]
rlabel metal2 42458 71128 42458 71128 0 sine_out_reg0\[5\]
rlabel metal1 43884 68918 43884 68918 0 sine_out_reg0\[6\]
rlabel metal1 62583 68986 62583 68986 0 sine_out_reg0\[7\]
rlabel metal1 67298 69462 67298 69462 0 sine_out_reg0\[8\]
rlabel metal1 68724 68918 68724 68918 0 sine_out_reg0\[9\]
rlabel metal1 7360 93670 7360 93670 0 sine_out_reg1\[0\]
rlabel metal2 74566 75072 74566 75072 0 sine_out_reg1\[10\]
rlabel metal1 98003 136850 98003 136850 0 sine_out_reg1\[11\]
rlabel metal1 83398 76330 83398 76330 0 sine_out_reg1\[12\]
rlabel metal1 105800 113254 105800 113254 0 sine_out_reg1\[13\]
rlabel metal1 103914 80070 103914 80070 0 sine_out_reg1\[14\]
rlabel metal2 105754 96254 105754 96254 0 sine_out_reg1\[15\]
rlabel metal1 7452 100198 7452 100198 0 sine_out_reg1\[1\]
rlabel metal1 28290 76466 28290 76466 0 sine_out_reg1\[2\]
rlabel metal1 37720 73882 37720 73882 0 sine_out_reg1\[3\]
rlabel metal1 8234 102170 8234 102170 0 sine_out_reg1\[4\]
rlabel metal2 42918 74528 42918 74528 0 sine_out_reg1\[5\]
rlabel metal2 45494 74698 45494 74698 0 sine_out_reg1\[6\]
rlabel metal2 62146 76160 62146 76160 0 sine_out_reg1\[7\]
rlabel metal2 64262 76126 64262 76126 0 sine_out_reg1\[8\]
rlabel metal1 67988 76602 67988 76602 0 sine_out_reg1\[9\]
rlabel metal4 36107 63983 36107 63983 0 sine_out_temp0\[0\]
rlabel metal4 61134 64260 61134 64260 0 sine_out_temp0\[10\]
rlabel metal4 63572 66771 63572 66771 0 sine_out_temp0\[11\]
rlabel metal4 66059 63847 66059 63847 0 sine_out_temp0\[12\]
rlabel metal1 79472 70890 79472 70890 0 sine_out_temp0\[13\]
rlabel via1 77873 69802 77873 69802 0 sine_out_temp0\[14\]
rlabel via2 79350 69853 79350 69853 0 sine_out_temp0\[15\]
rlabel metal4 38575 64260 38575 64260 0 sine_out_temp0\[1\]
rlabel metal4 41099 63983 41099 63983 0 sine_out_temp0\[2\]
rlabel metal4 43595 63915 43595 63915 0 sine_out_temp0\[3\]
rlabel metal2 45126 67711 45126 67711 0 sine_out_temp0\[4\]
rlabel metal1 43664 69394 43664 69394 0 sine_out_temp0\[5\]
rlabel metal3 48794 64124 48794 64124 0 sine_out_temp0\[6\]
rlabel via2 58742 68731 58742 68731 0 sine_out_temp0\[7\]
rlabel metal4 56075 63983 56075 63983 0 sine_out_temp0\[8\]
rlabel metal4 58571 63915 58571 63915 0 sine_out_temp0\[9\]
rlabel metal2 36018 135065 36018 135065 0 sine_out_temp1\[0\]
rlabel metal4 61088 134003 61088 134003 0 sine_out_temp1\[10\]
rlabel metal2 63618 135609 63618 135609 0 sine_out_temp1\[11\]
rlabel metal4 66059 133935 66059 133935 0 sine_out_temp1\[12\]
rlabel metal4 68555 133799 68555 133799 0 sine_out_temp1\[13\]
rlabel metal4 71051 134003 71051 134003 0 sine_out_temp1\[14\]
rlabel metal2 77418 135303 77418 135303 0 sine_out_temp1\[15\]
rlabel metal1 36110 136204 36110 136204 0 sine_out_temp1\[1\]
rlabel metal4 41099 133935 41099 133935 0 sine_out_temp1\[2\]
rlabel metal4 43595 133935 43595 133935 0 sine_out_temp1\[3\]
rlabel metal1 7452 118490 7452 118490 0 sine_out_temp1\[4\]
rlabel metal4 48576 133799 48576 133799 0 sine_out_temp1\[5\]
rlabel metal4 51083 133799 51083 133799 0 sine_out_temp1\[6\]
rlabel metal2 55430 135167 55430 135167 0 sine_out_temp1\[7\]
rlabel metal4 56075 133935 56075 133935 0 sine_out_temp1\[8\]
rlabel metal4 58571 134003 58571 134003 0 sine_out_temp1\[9\]
rlabel metal4 87342 133799 87342 133799 0 tcout\[0\]
rlabel metal1 93242 70924 93242 70924 0 tcout\[1\]
rlabel via2 102279 25060 102279 25060 0 tcout\[2\]
rlabel metal3 102095 23360 102095 23360 0 tcout\[3\]
rlabel metal3 102072 22232 102072 22232 0 tcout\[4\]
rlabel metal2 90574 7939 90574 7939 0 tcout\[5\]
rlabel metal1 90712 7514 90712 7514 0 tcout\[6\]
rlabel metal1 90896 7514 90896 7514 0 tcout\[7\]
rlabel metal1 87768 69394 87768 69394 0 tcout\[8\]
rlabel metal1 76866 74222 76866 74222 0 tcout_delay\[0\]
rlabel metal2 82018 72658 82018 72658 0 tcout_delay\[1\]
<< properties >>
string FIXED_BBOX 0 0 110000 150000
<< end >>
