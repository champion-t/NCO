magic
tech sky130A
magscale 1 2
timestamp 1741069072
<< viali >>
rect 44649 71689 44683 71723
rect 47225 71689 47259 71723
rect 49893 71689 49927 71723
rect 51825 71689 51859 71723
rect 53757 71689 53791 71723
rect 55689 71689 55723 71723
rect 57621 71689 57655 71723
rect 59461 71689 59495 71723
rect 61393 71689 61427 71723
rect 63417 71689 63451 71723
rect 65993 71689 66027 71723
rect 67925 71689 67959 71723
rect 69765 71689 69799 71723
rect 71697 71689 71731 71723
rect 74365 71689 74399 71723
rect 77585 71689 77619 71723
rect 44833 71553 44867 71587
rect 47409 71553 47443 71587
rect 49709 71553 49743 71587
rect 51641 71553 51675 71587
rect 53573 71553 53607 71587
rect 55505 71553 55539 71587
rect 57437 71553 57471 71587
rect 59645 71553 59679 71587
rect 61577 71553 61611 71587
rect 63233 71553 63267 71587
rect 65809 71553 65843 71587
rect 67741 71553 67775 71587
rect 69949 71553 69983 71587
rect 71881 71553 71915 71587
rect 74181 71553 74215 71587
rect 77401 71553 77435 71587
rect 45201 67337 45235 67371
rect 49525 67337 49559 67371
rect 51457 67337 51491 67371
rect 55321 67337 55355 67371
rect 57161 67337 57195 67371
rect 59645 67337 59679 67371
rect 61485 67337 61519 67371
rect 65441 67337 65475 67371
rect 67373 67337 67407 67371
rect 69949 67337 69983 67371
rect 71789 67337 71823 67371
rect 76113 67337 76147 67371
rect 70317 67269 70351 67303
rect 74641 67269 74675 67303
rect 45569 67201 45603 67235
rect 47777 67201 47811 67235
rect 65625 67201 65659 67235
rect 43361 67133 43395 67167
rect 43637 67133 43671 67167
rect 45109 67133 45143 67167
rect 45845 67133 45879 67167
rect 47317 67133 47351 67167
rect 48053 67133 48087 67167
rect 49709 67133 49743 67167
rect 49985 67133 50019 67167
rect 51549 67133 51583 67167
rect 53573 67133 53607 67167
rect 53849 67133 53883 67167
rect 55413 67133 55447 67167
rect 55689 67133 55723 67167
rect 57345 67133 57379 67167
rect 57713 67133 57747 67167
rect 57897 67133 57931 67167
rect 58173 67133 58207 67167
rect 59737 67133 59771 67167
rect 60013 67133 60047 67167
rect 63693 67133 63727 67167
rect 63969 67133 64003 67167
rect 65901 67133 65935 67167
rect 68201 67133 68235 67167
rect 68477 67133 68511 67167
rect 70041 67133 70075 67167
rect 74365 67133 74399 67167
rect 43177 66997 43211 67031
rect 45385 66997 45419 67031
rect 47593 66997 47627 67031
rect 51733 66997 51767 67031
rect 63601 66997 63635 67031
rect 68017 66997 68051 67031
rect 76297 66997 76331 67031
rect 47685 66793 47719 66827
rect 49709 66793 49743 66827
rect 53389 66793 53423 66827
rect 59645 66793 59679 66827
rect 61301 66793 61335 66827
rect 65717 66793 65751 66827
rect 69949 66793 69983 66827
rect 73721 66793 73755 66827
rect 63141 66725 63175 66759
rect 51641 66657 51675 66691
rect 53481 66657 53515 66691
rect 61393 66657 61427 66691
rect 71789 66657 71823 66691
rect 51917 66521 51951 66555
rect 61669 66521 61703 66555
rect 72065 66521 72099 66555
rect 55505 66453 55539 66487
rect 73537 66453 73571 66487
rect 56425 66249 56459 66283
rect 75561 66249 75595 66283
rect 48697 66181 48731 66215
rect 50537 66181 50571 66215
rect 52469 66181 52503 66215
rect 54033 66181 54067 66215
rect 55689 66181 55723 66215
rect 58449 66181 58483 66215
rect 60841 66181 60875 66215
rect 64889 66181 64923 66215
rect 66269 66181 66303 66215
rect 67925 66181 67959 66215
rect 69581 66181 69615 66215
rect 71421 66181 71455 66215
rect 73445 66181 73479 66215
rect 76021 66181 76055 66215
rect 95893 66181 95927 66215
rect 48789 66113 48823 66147
rect 50629 66113 50663 66147
rect 52561 66113 52595 66147
rect 54125 66113 54159 66147
rect 55781 66113 55815 66147
rect 57713 66113 57747 66147
rect 57989 66113 58023 66147
rect 58081 66113 58115 66147
rect 59093 66113 59127 66147
rect 60933 66113 60967 66147
rect 62865 66113 62899 66147
rect 63233 66113 63267 66147
rect 64429 66113 64463 66147
rect 64705 66113 64739 66147
rect 64797 66113 64831 66147
rect 66361 66113 66395 66147
rect 68017 66113 68051 66147
rect 69673 66113 69707 66147
rect 71513 66113 71547 66147
rect 73537 66113 73571 66147
rect 75745 66113 75779 66147
rect 75929 66113 75963 66147
rect 91937 66113 91971 66147
rect 92397 66113 92431 66147
rect 58265 65977 58299 66011
rect 61577 65977 61611 66011
rect 63601 65977 63635 66011
rect 59001 65909 59035 65943
rect 63141 65909 63175 65943
rect 63417 65909 63451 65943
rect 65165 65909 65199 65943
rect 76205 65909 76239 65943
rect 86325 65909 86359 65943
rect 87337 65909 87371 65943
rect 92029 65909 92063 65943
rect 92305 65909 92339 65943
rect 104357 60061 104391 60095
rect 104357 57749 104391 57783
rect 104357 57409 104391 57443
rect 104633 57341 104667 57375
rect 106381 57341 106415 57375
rect 106473 57341 106507 57375
rect 106657 57205 106691 57239
rect 105001 56865 105035 56899
rect 105185 56865 105219 56899
rect 104449 56661 104483 56695
rect 104449 55913 104483 55947
rect 104541 55709 104575 55743
rect 104357 54689 104391 54723
rect 106749 54689 106783 54723
rect 104633 54553 104667 54587
rect 106381 54553 106415 54587
rect 106473 54553 106507 54587
rect 104449 54281 104483 54315
rect 104357 54145 104391 54179
rect 104633 53941 104667 53975
rect 104357 53737 104391 53771
rect 105001 53737 105035 53771
rect 104633 53601 104667 53635
rect 105185 53601 105219 53635
rect 104725 53533 104759 53567
rect 104817 46121 104851 46155
rect 104357 46053 104391 46087
rect 104541 45917 104575 45951
rect 104633 45917 104667 45951
rect 104357 45849 104391 45883
rect 104909 45781 104943 45815
rect 105185 45781 105219 45815
rect 104541 45033 104575 45067
rect 105277 45033 105311 45067
rect 105093 44965 105127 44999
rect 104357 44761 104391 44795
rect 104541 44693 104575 44727
rect 104725 44693 104759 44727
rect 104909 44693 104943 44727
rect 105461 44693 105495 44727
rect 104633 43945 104667 43979
rect 104357 43741 104391 43775
rect 104449 43673 104483 43707
rect 104357 42721 104391 42755
rect 104633 42585 104667 42619
rect 106105 42517 106139 42551
rect 106197 42517 106231 42551
rect 106381 42517 106415 42551
rect 104541 42177 104575 42211
rect 106565 41973 106599 42007
rect 104357 41565 104391 41599
rect 106105 41497 106139 41531
rect 106197 41497 106231 41531
rect 7573 41429 7607 41463
rect 104449 41225 104483 41259
rect 104909 41225 104943 41259
rect 104357 41089 104391 41123
rect 104541 41089 104575 41123
rect 104725 40885 104759 40919
rect 7573 39797 7607 39831
rect 7573 38709 7607 38743
rect 104633 36873 104667 36907
rect 7573 36737 7607 36771
rect 104357 36737 104391 36771
rect 104449 36533 104483 36567
rect 104357 35649 104391 35683
rect 7573 35513 7607 35547
rect 104449 35445 104483 35479
rect 104725 35445 104759 35479
rect 7573 34017 7607 34051
rect 106105 33949 106139 33983
rect 105829 33881 105863 33915
rect 104357 33813 104391 33847
rect 106197 33813 106231 33847
rect 104817 33405 104851 33439
rect 105369 33269 105403 33303
rect 105829 32929 105863 32963
rect 106105 32861 106139 32895
rect 104357 32725 104391 32759
rect 106289 32725 106323 32759
rect 105277 32385 105311 32419
rect 104541 32317 104575 32351
rect 105369 32317 105403 32351
rect 106013 31977 106047 32011
rect 110337 31977 110371 32011
rect 104449 31909 104483 31943
rect 106105 31909 106139 31943
rect 105737 31841 105771 31875
rect 104357 31773 104391 31807
rect 104725 31773 104759 31807
rect 105369 31773 105403 31807
rect 105645 31773 105679 31807
rect 110245 31773 110279 31807
rect 110521 31773 110555 31807
rect 104633 31093 104667 31127
rect 105829 30277 105863 30311
rect 105001 30209 105035 30243
rect 105461 30209 105495 30243
rect 105645 30209 105679 30243
rect 105093 30141 105127 30175
rect 105553 30141 105587 30175
rect 105369 30073 105403 30107
rect 104357 29597 104391 29631
rect 104449 29461 104483 29495
rect 104725 29461 104759 29495
rect 104357 28577 104391 28611
rect 104633 28441 104667 28475
rect 106105 28373 106139 28407
rect 106289 28373 106323 28407
rect 106473 28373 106507 28407
rect 104725 28169 104759 28203
rect 104817 28101 104851 28135
rect 105033 28101 105067 28135
rect 105001 27829 105035 27863
rect 105185 27829 105219 27863
rect 104449 27081 104483 27115
rect 104633 27081 104667 27115
rect 105185 27081 105219 27115
rect 105461 27081 105495 27115
rect 104630 26945 104664 26979
rect 105001 26945 105035 26979
rect 105093 26945 105127 26979
rect 104357 25857 104391 25891
rect 104633 25789 104667 25823
rect 106105 25653 106139 25687
rect 106197 25653 106231 25687
rect 106381 25653 106415 25687
rect 104541 25449 104575 25483
rect 104725 25449 104759 25483
rect 104817 25245 104851 25279
rect 105093 25245 105127 25279
rect 104357 25177 104391 25211
rect 105277 25177 105311 25211
rect 104557 25109 104591 25143
rect 104909 25109 104943 25143
rect 104357 24769 104391 24803
rect 104817 24361 104851 24395
rect 104541 24157 104575 24191
rect 104633 24157 104667 24191
rect 104357 24089 104391 24123
rect 104909 24089 104943 24123
rect 104455 24021 104489 24055
rect 104567 23817 104601 23851
rect 105093 23817 105127 23851
rect 105277 23817 105311 23851
rect 104357 23749 104391 23783
rect 104817 23681 104851 23715
rect 105001 23681 105035 23715
rect 104817 23545 104851 23579
rect 104541 23477 104575 23511
rect 104725 23477 104759 23511
rect 104357 20961 104391 20995
rect 106381 20961 106415 20995
rect 104633 20825 104667 20859
rect 106105 20757 106139 20791
rect 106197 20757 106231 20791
rect 105001 20349 105035 20383
rect 104449 20213 104483 20247
rect 104357 19669 104391 19703
rect 104725 19329 104759 19363
rect 104357 19261 104391 19295
rect 104633 19261 104667 19295
rect 7573 15521 7607 15555
rect 16129 7497 16163 7531
rect 23489 7497 23523 7531
rect 24685 7497 24719 7531
rect 25881 7497 25915 7531
rect 26985 7497 27019 7531
rect 28273 7497 28307 7531
rect 29561 7497 29595 7531
rect 30481 7497 30515 7531
rect 31769 7497 31803 7531
rect 32873 7497 32907 7531
rect 33977 7497 34011 7531
rect 35265 7497 35299 7531
rect 36369 7497 36403 7531
rect 37473 7497 37507 7531
rect 38669 7497 38703 7531
rect 39865 7497 39899 7531
rect 41061 7497 41095 7531
rect 42165 7497 42199 7531
rect 43361 7497 43395 7531
rect 90557 7497 90591 7531
rect 90741 7497 90775 7531
rect 91017 7497 91051 7531
<< metal1 >>
rect 1104 71834 110860 71856
rect 1104 71782 4874 71834
rect 4926 71782 4938 71834
rect 4990 71782 5002 71834
rect 5054 71782 5066 71834
rect 5118 71782 5130 71834
rect 5182 71782 35594 71834
rect 35646 71782 35658 71834
rect 35710 71782 35722 71834
rect 35774 71782 35786 71834
rect 35838 71782 35850 71834
rect 35902 71782 66314 71834
rect 66366 71782 66378 71834
rect 66430 71782 66442 71834
rect 66494 71782 66506 71834
rect 66558 71782 66570 71834
rect 66622 71782 97034 71834
rect 97086 71782 97098 71834
rect 97150 71782 97162 71834
rect 97214 71782 97226 71834
rect 97278 71782 97290 71834
rect 97342 71782 110860 71834
rect 1104 71760 110860 71782
rect 44450 71680 44456 71732
rect 44508 71720 44514 71732
rect 44637 71723 44695 71729
rect 44637 71720 44649 71723
rect 44508 71692 44649 71720
rect 44508 71680 44514 71692
rect 44637 71689 44649 71692
rect 44683 71689 44695 71723
rect 44637 71683 44695 71689
rect 47026 71680 47032 71732
rect 47084 71720 47090 71732
rect 47213 71723 47271 71729
rect 47213 71720 47225 71723
rect 47084 71692 47225 71720
rect 47084 71680 47090 71692
rect 47213 71689 47225 71692
rect 47259 71689 47271 71723
rect 47213 71683 47271 71689
rect 49602 71680 49608 71732
rect 49660 71720 49666 71732
rect 49881 71723 49939 71729
rect 49881 71720 49893 71723
rect 49660 71692 49893 71720
rect 49660 71680 49666 71692
rect 49881 71689 49893 71692
rect 49927 71689 49939 71723
rect 49881 71683 49939 71689
rect 51534 71680 51540 71732
rect 51592 71720 51598 71732
rect 51813 71723 51871 71729
rect 51813 71720 51825 71723
rect 51592 71692 51825 71720
rect 51592 71680 51598 71692
rect 51813 71689 51825 71692
rect 51859 71689 51871 71723
rect 51813 71683 51871 71689
rect 53466 71680 53472 71732
rect 53524 71720 53530 71732
rect 53745 71723 53803 71729
rect 53745 71720 53757 71723
rect 53524 71692 53757 71720
rect 53524 71680 53530 71692
rect 53745 71689 53757 71692
rect 53791 71689 53803 71723
rect 53745 71683 53803 71689
rect 55398 71680 55404 71732
rect 55456 71720 55462 71732
rect 55677 71723 55735 71729
rect 55677 71720 55689 71723
rect 55456 71692 55689 71720
rect 55456 71680 55462 71692
rect 55677 71689 55689 71692
rect 55723 71689 55735 71723
rect 55677 71683 55735 71689
rect 57330 71680 57336 71732
rect 57388 71720 57394 71732
rect 57609 71723 57667 71729
rect 57609 71720 57621 71723
rect 57388 71692 57621 71720
rect 57388 71680 57394 71692
rect 57609 71689 57621 71692
rect 57655 71689 57667 71723
rect 57609 71683 57667 71689
rect 59262 71680 59268 71732
rect 59320 71720 59326 71732
rect 59449 71723 59507 71729
rect 59449 71720 59461 71723
rect 59320 71692 59461 71720
rect 59320 71680 59326 71692
rect 59449 71689 59461 71692
rect 59495 71689 59507 71723
rect 59449 71683 59507 71689
rect 61194 71680 61200 71732
rect 61252 71720 61258 71732
rect 61381 71723 61439 71729
rect 61381 71720 61393 71723
rect 61252 71692 61393 71720
rect 61252 71680 61258 71692
rect 61381 71689 61393 71692
rect 61427 71689 61439 71723
rect 61381 71683 61439 71689
rect 63126 71680 63132 71732
rect 63184 71720 63190 71732
rect 63405 71723 63463 71729
rect 63405 71720 63417 71723
rect 63184 71692 63417 71720
rect 63184 71680 63190 71692
rect 63405 71689 63417 71692
rect 63451 71689 63463 71723
rect 63405 71683 63463 71689
rect 65702 71680 65708 71732
rect 65760 71720 65766 71732
rect 65981 71723 66039 71729
rect 65981 71720 65993 71723
rect 65760 71692 65993 71720
rect 65760 71680 65766 71692
rect 65981 71689 65993 71692
rect 66027 71689 66039 71723
rect 65981 71683 66039 71689
rect 67634 71680 67640 71732
rect 67692 71720 67698 71732
rect 67913 71723 67971 71729
rect 67913 71720 67925 71723
rect 67692 71692 67925 71720
rect 67692 71680 67698 71692
rect 67913 71689 67925 71692
rect 67959 71689 67971 71723
rect 67913 71683 67971 71689
rect 69566 71680 69572 71732
rect 69624 71720 69630 71732
rect 69753 71723 69811 71729
rect 69753 71720 69765 71723
rect 69624 71692 69765 71720
rect 69624 71680 69630 71692
rect 69753 71689 69765 71692
rect 69799 71689 69811 71723
rect 69753 71683 69811 71689
rect 71498 71680 71504 71732
rect 71556 71720 71562 71732
rect 71685 71723 71743 71729
rect 71685 71720 71697 71723
rect 71556 71692 71697 71720
rect 71556 71680 71562 71692
rect 71685 71689 71697 71692
rect 71731 71689 71743 71723
rect 71685 71683 71743 71689
rect 74074 71680 74080 71732
rect 74132 71720 74138 71732
rect 74353 71723 74411 71729
rect 74353 71720 74365 71723
rect 74132 71692 74365 71720
rect 74132 71680 74138 71692
rect 74353 71689 74365 71692
rect 74399 71689 74411 71723
rect 74353 71683 74411 71689
rect 77294 71680 77300 71732
rect 77352 71720 77358 71732
rect 77573 71723 77631 71729
rect 77573 71720 77585 71723
rect 77352 71692 77585 71720
rect 77352 71680 77358 71692
rect 77573 71689 77585 71692
rect 77619 71689 77631 71723
rect 77573 71683 77631 71689
rect 44821 71587 44879 71593
rect 44821 71553 44833 71587
rect 44867 71584 44879 71587
rect 45094 71584 45100 71596
rect 44867 71556 45100 71584
rect 44867 71553 44879 71556
rect 44821 71547 44879 71553
rect 45094 71544 45100 71556
rect 45152 71544 45158 71596
rect 47302 71544 47308 71596
rect 47360 71584 47366 71596
rect 47397 71587 47455 71593
rect 47397 71584 47409 71587
rect 47360 71556 47409 71584
rect 47360 71544 47366 71556
rect 47397 71553 47409 71556
rect 47443 71553 47455 71587
rect 47397 71547 47455 71553
rect 49510 71544 49516 71596
rect 49568 71584 49574 71596
rect 49697 71587 49755 71593
rect 49697 71584 49709 71587
rect 49568 71556 49709 71584
rect 49568 71544 49574 71556
rect 49697 71553 49709 71556
rect 49743 71553 49755 71587
rect 49697 71547 49755 71553
rect 51626 71544 51632 71596
rect 51684 71544 51690 71596
rect 53558 71544 53564 71596
rect 53616 71544 53622 71596
rect 55490 71544 55496 71596
rect 55548 71544 55554 71596
rect 57422 71544 57428 71596
rect 57480 71544 57486 71596
rect 59630 71544 59636 71596
rect 59688 71544 59694 71596
rect 61562 71544 61568 71596
rect 61620 71544 61626 71596
rect 63126 71544 63132 71596
rect 63184 71584 63190 71596
rect 63221 71587 63279 71593
rect 63221 71584 63233 71587
rect 63184 71556 63233 71584
rect 63184 71544 63190 71556
rect 63221 71553 63233 71556
rect 63267 71553 63279 71587
rect 63221 71547 63279 71553
rect 65426 71544 65432 71596
rect 65484 71584 65490 71596
rect 65797 71587 65855 71593
rect 65797 71584 65809 71587
rect 65484 71556 65809 71584
rect 65484 71544 65490 71556
rect 65797 71553 65809 71556
rect 65843 71553 65855 71587
rect 65797 71547 65855 71553
rect 67358 71544 67364 71596
rect 67416 71584 67422 71596
rect 67729 71587 67787 71593
rect 67729 71584 67741 71587
rect 67416 71556 67741 71584
rect 67416 71544 67422 71556
rect 67729 71553 67741 71556
rect 67775 71553 67787 71587
rect 67729 71547 67787 71553
rect 69934 71544 69940 71596
rect 69992 71544 69998 71596
rect 71866 71544 71872 71596
rect 71924 71544 71930 71596
rect 74166 71544 74172 71596
rect 74224 71544 74230 71596
rect 76098 71544 76104 71596
rect 76156 71584 76162 71596
rect 77389 71587 77447 71593
rect 77389 71584 77401 71587
rect 76156 71556 77401 71584
rect 76156 71544 76162 71556
rect 77389 71553 77401 71556
rect 77435 71553 77447 71587
rect 77389 71547 77447 71553
rect 1104 71290 110860 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 34934 71290
rect 34986 71238 34998 71290
rect 35050 71238 35062 71290
rect 35114 71238 35126 71290
rect 35178 71238 35190 71290
rect 35242 71238 65654 71290
rect 65706 71238 65718 71290
rect 65770 71238 65782 71290
rect 65834 71238 65846 71290
rect 65898 71238 65910 71290
rect 65962 71238 96374 71290
rect 96426 71238 96438 71290
rect 96490 71238 96502 71290
rect 96554 71238 96566 71290
rect 96618 71238 96630 71290
rect 96682 71238 110860 71290
rect 1104 71216 110860 71238
rect 1104 70746 110860 70768
rect 1104 70694 4874 70746
rect 4926 70694 4938 70746
rect 4990 70694 5002 70746
rect 5054 70694 5066 70746
rect 5118 70694 5130 70746
rect 5182 70694 35594 70746
rect 35646 70694 35658 70746
rect 35710 70694 35722 70746
rect 35774 70694 35786 70746
rect 35838 70694 35850 70746
rect 35902 70694 66314 70746
rect 66366 70694 66378 70746
rect 66430 70694 66442 70746
rect 66494 70694 66506 70746
rect 66558 70694 66570 70746
rect 66622 70694 97034 70746
rect 97086 70694 97098 70746
rect 97150 70694 97162 70746
rect 97214 70694 97226 70746
rect 97278 70694 97290 70746
rect 97342 70694 110860 70746
rect 1104 70672 110860 70694
rect 1104 70202 110860 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 34934 70202
rect 34986 70150 34998 70202
rect 35050 70150 35062 70202
rect 35114 70150 35126 70202
rect 35178 70150 35190 70202
rect 35242 70150 65654 70202
rect 65706 70150 65718 70202
rect 65770 70150 65782 70202
rect 65834 70150 65846 70202
rect 65898 70150 65910 70202
rect 65962 70150 96374 70202
rect 96426 70150 96438 70202
rect 96490 70150 96502 70202
rect 96554 70150 96566 70202
rect 96618 70150 96630 70202
rect 96682 70150 110860 70202
rect 1104 70128 110860 70150
rect 1104 69658 110860 69680
rect 1104 69606 4874 69658
rect 4926 69606 4938 69658
rect 4990 69606 5002 69658
rect 5054 69606 5066 69658
rect 5118 69606 5130 69658
rect 5182 69606 35594 69658
rect 35646 69606 35658 69658
rect 35710 69606 35722 69658
rect 35774 69606 35786 69658
rect 35838 69606 35850 69658
rect 35902 69606 66314 69658
rect 66366 69606 66378 69658
rect 66430 69606 66442 69658
rect 66494 69606 66506 69658
rect 66558 69606 66570 69658
rect 66622 69606 97034 69658
rect 97086 69606 97098 69658
rect 97150 69606 97162 69658
rect 97214 69606 97226 69658
rect 97278 69606 97290 69658
rect 97342 69606 110860 69658
rect 1104 69584 110860 69606
rect 1104 69114 110860 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 96374 69114
rect 96426 69062 96438 69114
rect 96490 69062 96502 69114
rect 96554 69062 96566 69114
rect 96618 69062 96630 69114
rect 96682 69062 110860 69114
rect 1104 69040 110860 69062
rect 1104 68570 110860 68592
rect 1104 68518 4874 68570
rect 4926 68518 4938 68570
rect 4990 68518 5002 68570
rect 5054 68518 5066 68570
rect 5118 68518 5130 68570
rect 5182 68518 35594 68570
rect 35646 68518 35658 68570
rect 35710 68518 35722 68570
rect 35774 68518 35786 68570
rect 35838 68518 35850 68570
rect 35902 68518 66314 68570
rect 66366 68518 66378 68570
rect 66430 68518 66442 68570
rect 66494 68518 66506 68570
rect 66558 68518 66570 68570
rect 66622 68518 97034 68570
rect 97086 68518 97098 68570
rect 97150 68518 97162 68570
rect 97214 68518 97226 68570
rect 97278 68518 97290 68570
rect 97342 68518 110860 68570
rect 1104 68496 110860 68518
rect 1104 68026 110860 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 96374 68026
rect 96426 67974 96438 68026
rect 96490 67974 96502 68026
rect 96554 67974 96566 68026
rect 96618 67974 96630 68026
rect 96682 67974 110860 68026
rect 1104 67952 110860 67974
rect 1104 67482 110860 67504
rect 1104 67430 4874 67482
rect 4926 67430 4938 67482
rect 4990 67430 5002 67482
rect 5054 67430 5066 67482
rect 5118 67430 5130 67482
rect 5182 67430 35594 67482
rect 35646 67430 35658 67482
rect 35710 67430 35722 67482
rect 35774 67430 35786 67482
rect 35838 67430 35850 67482
rect 35902 67430 66314 67482
rect 66366 67430 66378 67482
rect 66430 67430 66442 67482
rect 66494 67430 66506 67482
rect 66558 67430 66570 67482
rect 66622 67430 97034 67482
rect 97086 67430 97098 67482
rect 97150 67430 97162 67482
rect 97214 67430 97226 67482
rect 97278 67430 97290 67482
rect 97342 67430 110860 67482
rect 1104 67408 110860 67430
rect 45189 67371 45247 67377
rect 45189 67368 45201 67371
rect 43364 67340 45201 67368
rect 8202 67124 8208 67176
rect 8260 67164 8266 67176
rect 43364 67173 43392 67340
rect 45189 67337 45201 67340
rect 45235 67368 45247 67371
rect 45235 67340 47624 67368
rect 45235 67337 45247 67340
rect 45189 67331 45247 67337
rect 44726 67192 44732 67244
rect 44784 67192 44790 67244
rect 45480 67232 45508 67340
rect 45557 67235 45615 67241
rect 45557 67232 45569 67235
rect 45480 67204 45569 67232
rect 45557 67201 45569 67204
rect 45603 67201 45615 67235
rect 45557 67195 45615 67201
rect 46934 67192 46940 67244
rect 46992 67192 46998 67244
rect 47596 67232 47624 67340
rect 49510 67328 49516 67380
rect 49568 67328 49574 67380
rect 51445 67371 51503 67377
rect 51445 67337 51457 67371
rect 51491 67368 51503 67371
rect 51626 67368 51632 67380
rect 51491 67340 51632 67368
rect 51491 67337 51503 67340
rect 51445 67331 51503 67337
rect 51626 67328 51632 67340
rect 51684 67328 51690 67380
rect 55309 67371 55367 67377
rect 55309 67337 55321 67371
rect 55355 67368 55367 67371
rect 55490 67368 55496 67380
rect 55355 67340 55496 67368
rect 55355 67337 55367 67340
rect 55309 67331 55367 67337
rect 55490 67328 55496 67340
rect 55548 67328 55554 67380
rect 57149 67371 57207 67377
rect 57149 67337 57161 67371
rect 57195 67368 57207 67371
rect 57422 67368 57428 67380
rect 57195 67340 57428 67368
rect 57195 67337 57207 67340
rect 57149 67331 57207 67337
rect 57422 67328 57428 67340
rect 57480 67328 57486 67380
rect 59630 67328 59636 67380
rect 59688 67328 59694 67380
rect 60826 67368 60832 67380
rect 60384 67340 60832 67368
rect 53926 67300 53932 67312
rect 51198 67272 53932 67300
rect 53926 67260 53932 67272
rect 53984 67260 53990 67312
rect 57790 67300 57796 67312
rect 56902 67272 57796 67300
rect 57790 67260 57796 67272
rect 57848 67260 57854 67312
rect 60384 67300 60412 67340
rect 60826 67328 60832 67340
rect 60884 67328 60890 67380
rect 61473 67371 61531 67377
rect 61473 67337 61485 67371
rect 61519 67368 61531 67371
rect 61562 67368 61568 67380
rect 61519 67340 61568 67368
rect 61519 67337 61531 67340
rect 61473 67331 61531 67337
rect 61562 67328 61568 67340
rect 61620 67328 61626 67380
rect 65426 67328 65432 67380
rect 65484 67328 65490 67380
rect 67358 67328 67364 67380
rect 67416 67328 67422 67380
rect 68738 67328 68744 67380
rect 68796 67368 68802 67380
rect 68796 67340 69796 67368
rect 68796 67328 68802 67340
rect 62022 67300 62028 67312
rect 59386 67272 60412 67300
rect 61226 67272 62028 67300
rect 62022 67260 62028 67272
rect 62080 67260 62086 67312
rect 66162 67300 66168 67312
rect 65182 67272 66168 67300
rect 66162 67260 66168 67272
rect 66220 67260 66226 67312
rect 67542 67300 67548 67312
rect 67114 67272 67548 67300
rect 67542 67260 67548 67272
rect 67600 67260 67606 67312
rect 69768 67300 69796 67340
rect 69934 67328 69940 67380
rect 69992 67328 69998 67380
rect 71777 67371 71835 67377
rect 71777 67337 71789 67371
rect 71823 67368 71835 67371
rect 71866 67368 71872 67380
rect 71823 67340 71872 67368
rect 71823 67337 71835 67340
rect 71777 67331 71835 67337
rect 71866 67328 71872 67340
rect 71924 67328 71930 67380
rect 76098 67328 76104 67380
rect 76156 67328 76162 67380
rect 70305 67303 70363 67309
rect 70305 67300 70317 67303
rect 69768 67272 70317 67300
rect 70305 67269 70317 67272
rect 70351 67269 70363 67303
rect 70305 67263 70363 67269
rect 74074 67260 74080 67312
rect 74132 67300 74138 67312
rect 74629 67303 74687 67309
rect 74629 67300 74641 67303
rect 74132 67272 74641 67300
rect 74132 67260 74138 67272
rect 74629 67269 74641 67272
rect 74675 67269 74687 67303
rect 74629 67263 74687 67269
rect 47670 67232 47676 67244
rect 47596 67204 47676 67232
rect 47670 67192 47676 67204
rect 47728 67232 47734 67244
rect 47765 67235 47823 67241
rect 47765 67232 47777 67235
rect 47728 67204 47777 67232
rect 47728 67192 47734 67204
rect 47765 67201 47777 67204
rect 47811 67201 47823 67235
rect 47765 67195 47823 67201
rect 49142 67192 49148 67244
rect 49200 67192 49206 67244
rect 54938 67192 54944 67244
rect 54996 67192 55002 67244
rect 65518 67192 65524 67244
rect 65576 67232 65582 67244
rect 65613 67235 65671 67241
rect 65613 67232 65625 67235
rect 65576 67204 65625 67232
rect 65576 67192 65582 67204
rect 65613 67201 65625 67204
rect 65659 67201 65671 67235
rect 65613 67195 65671 67201
rect 69566 67192 69572 67244
rect 69624 67192 69630 67244
rect 71406 67192 71412 67244
rect 71464 67192 71470 67244
rect 75730 67192 75736 67244
rect 75788 67192 75794 67244
rect 43349 67167 43407 67173
rect 43349 67164 43361 67167
rect 8260 67136 43361 67164
rect 8260 67124 8266 67136
rect 43349 67133 43361 67136
rect 43395 67133 43407 67167
rect 43625 67167 43683 67173
rect 43625 67164 43637 67167
rect 43349 67127 43407 67133
rect 43456 67136 43637 67164
rect 43162 66988 43168 67040
rect 43220 67028 43226 67040
rect 43456 67028 43484 67136
rect 43625 67133 43637 67136
rect 43671 67133 43683 67167
rect 43625 67127 43683 67133
rect 45094 67124 45100 67176
rect 45152 67124 45158 67176
rect 45833 67167 45891 67173
rect 45833 67164 45845 67167
rect 45526 67136 45845 67164
rect 43220 67000 43484 67028
rect 43220 66988 43226 67000
rect 45370 66988 45376 67040
rect 45428 67028 45434 67040
rect 45526 67028 45554 67136
rect 45833 67133 45845 67136
rect 45879 67133 45891 67167
rect 45833 67127 45891 67133
rect 47302 67124 47308 67176
rect 47360 67124 47366 67176
rect 48041 67167 48099 67173
rect 48041 67164 48053 67167
rect 47596 67136 48053 67164
rect 47596 67040 47624 67136
rect 48041 67133 48053 67136
rect 48087 67133 48099 67167
rect 48041 67127 48099 67133
rect 49694 67124 49700 67176
rect 49752 67124 49758 67176
rect 49970 67124 49976 67176
rect 50028 67164 50034 67176
rect 51537 67167 51595 67173
rect 51537 67164 51549 67167
rect 50028 67136 51549 67164
rect 50028 67124 50034 67136
rect 51537 67133 51549 67136
rect 51583 67133 51595 67167
rect 51537 67127 51595 67133
rect 53466 67124 53472 67176
rect 53524 67164 53530 67176
rect 53561 67167 53619 67173
rect 53561 67164 53573 67167
rect 53524 67136 53573 67164
rect 53524 67124 53530 67136
rect 53561 67133 53573 67136
rect 53607 67133 53619 67167
rect 53837 67167 53895 67173
rect 53837 67164 53849 67167
rect 53561 67127 53619 67133
rect 53668 67136 53849 67164
rect 53668 67040 53696 67136
rect 53837 67133 53849 67136
rect 53883 67133 53895 67167
rect 53837 67127 53895 67133
rect 55398 67124 55404 67176
rect 55456 67124 55462 67176
rect 55674 67124 55680 67176
rect 55732 67124 55738 67176
rect 57333 67167 57391 67173
rect 57333 67133 57345 67167
rect 57379 67164 57391 67167
rect 57701 67167 57759 67173
rect 57701 67164 57713 67167
rect 57379 67136 57713 67164
rect 57379 67133 57391 67136
rect 57333 67127 57391 67133
rect 57701 67133 57713 67136
rect 57747 67164 57759 67167
rect 57882 67164 57888 67176
rect 57747 67136 57888 67164
rect 57747 67133 57759 67136
rect 57701 67127 57759 67133
rect 57882 67124 57888 67136
rect 57940 67124 57946 67176
rect 58158 67124 58164 67176
rect 58216 67124 58222 67176
rect 59722 67124 59728 67176
rect 59780 67124 59786 67176
rect 59998 67124 60004 67176
rect 60056 67124 60062 67176
rect 63681 67167 63739 67173
rect 63681 67133 63693 67167
rect 63727 67133 63739 67167
rect 63681 67127 63739 67133
rect 45428 67000 45554 67028
rect 45428 66988 45434 67000
rect 47578 66988 47584 67040
rect 47636 66988 47642 67040
rect 49694 66988 49700 67040
rect 49752 67028 49758 67040
rect 51626 67028 51632 67040
rect 49752 67000 51632 67028
rect 49752 66988 49758 67000
rect 51626 66988 51632 67000
rect 51684 67028 51690 67040
rect 51721 67031 51779 67037
rect 51721 67028 51733 67031
rect 51684 67000 51733 67028
rect 51684 66988 51690 67000
rect 51721 66997 51733 67000
rect 51767 66997 51779 67031
rect 51721 66991 51779 66997
rect 53650 66988 53656 67040
rect 53708 66988 53714 67040
rect 61286 66988 61292 67040
rect 61344 67028 61350 67040
rect 63589 67031 63647 67037
rect 63589 67028 63601 67031
rect 61344 67000 63601 67028
rect 61344 66988 61350 67000
rect 63589 66997 63601 67000
rect 63635 67028 63647 67031
rect 63696 67028 63724 67127
rect 63954 67124 63960 67176
rect 64012 67124 64018 67176
rect 64690 67124 64696 67176
rect 64748 67164 64754 67176
rect 65889 67167 65947 67173
rect 65889 67164 65901 67167
rect 64748 67136 65901 67164
rect 64748 67124 64754 67136
rect 65889 67133 65901 67136
rect 65935 67133 65947 67167
rect 65889 67127 65947 67133
rect 68189 67167 68247 67173
rect 68189 67133 68201 67167
rect 68235 67133 68247 67167
rect 68189 67127 68247 67133
rect 65518 67028 65524 67040
rect 63635 67000 65524 67028
rect 63635 66997 63647 67000
rect 63589 66991 63647 66997
rect 65518 66988 65524 67000
rect 65576 66988 65582 67040
rect 68002 66988 68008 67040
rect 68060 67028 68066 67040
rect 68204 67028 68232 67127
rect 68462 67124 68468 67176
rect 68520 67124 68526 67176
rect 69934 67124 69940 67176
rect 69992 67164 69998 67176
rect 70029 67167 70087 67173
rect 70029 67164 70041 67167
rect 69992 67136 70041 67164
rect 69992 67124 69998 67136
rect 70029 67133 70041 67136
rect 70075 67133 70087 67167
rect 70029 67127 70087 67133
rect 74353 67167 74411 67173
rect 74353 67133 74365 67167
rect 74399 67133 74411 67167
rect 74353 67127 74411 67133
rect 69934 67028 69940 67040
rect 68060 67000 69940 67028
rect 68060 66988 68066 67000
rect 69934 66988 69940 67000
rect 69992 66988 69998 67040
rect 73706 66988 73712 67040
rect 73764 67028 73770 67040
rect 74368 67028 74396 67127
rect 75656 67068 76328 67096
rect 75656 67028 75684 67068
rect 76300 67037 76328 67068
rect 73764 67000 75684 67028
rect 76285 67031 76343 67037
rect 73764 66988 73770 67000
rect 76285 66997 76297 67031
rect 76331 67028 76343 67031
rect 95878 67028 95884 67040
rect 76331 67000 95884 67028
rect 76331 66997 76343 67000
rect 76285 66991 76343 66997
rect 95878 66988 95884 67000
rect 95936 66988 95942 67040
rect 1104 66938 110860 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 96374 66938
rect 96426 66886 96438 66938
rect 96490 66886 96502 66938
rect 96554 66886 96566 66938
rect 96618 66886 96630 66938
rect 96682 66886 110860 66938
rect 1104 66864 110860 66886
rect 47670 66784 47676 66836
rect 47728 66824 47734 66836
rect 49694 66824 49700 66836
rect 47728 66796 49700 66824
rect 47728 66784 47734 66796
rect 49694 66784 49700 66796
rect 49752 66784 49758 66836
rect 53377 66827 53435 66833
rect 53377 66793 53389 66827
rect 53423 66824 53435 66827
rect 53558 66824 53564 66836
rect 53423 66796 53564 66824
rect 53423 66793 53435 66796
rect 53377 66787 53435 66793
rect 53558 66784 53564 66796
rect 53616 66784 53622 66836
rect 54938 66784 54944 66836
rect 54996 66824 55002 66836
rect 57974 66824 57980 66836
rect 54996 66796 57980 66824
rect 54996 66784 55002 66796
rect 57974 66784 57980 66796
rect 58032 66784 58038 66836
rect 59633 66827 59691 66833
rect 59633 66793 59645 66827
rect 59679 66824 59691 66827
rect 59722 66824 59728 66836
rect 59679 66796 59728 66824
rect 59679 66793 59691 66796
rect 59633 66787 59691 66793
rect 59722 66784 59728 66796
rect 59780 66824 59786 66836
rect 61286 66824 61292 66836
rect 59780 66796 61292 66824
rect 59780 66784 59786 66796
rect 61286 66784 61292 66796
rect 61344 66784 61350 66836
rect 65518 66784 65524 66836
rect 65576 66824 65582 66836
rect 65705 66827 65763 66833
rect 65705 66824 65717 66827
rect 65576 66796 65717 66824
rect 65576 66784 65582 66796
rect 65705 66793 65717 66796
rect 65751 66824 65763 66827
rect 68002 66824 68008 66836
rect 65751 66796 68008 66824
rect 65751 66793 65763 66796
rect 65705 66787 65763 66793
rect 68002 66784 68008 66796
rect 68060 66784 68066 66836
rect 69934 66784 69940 66836
rect 69992 66784 69998 66836
rect 73706 66784 73712 66836
rect 73764 66784 73770 66836
rect 44726 66716 44732 66768
rect 44784 66756 44790 66768
rect 48682 66756 48688 66768
rect 44784 66728 48688 66756
rect 44784 66716 44790 66728
rect 48682 66716 48688 66728
rect 48740 66716 48746 66768
rect 46934 66648 46940 66700
rect 46992 66688 46998 66700
rect 50522 66688 50528 66700
rect 46992 66660 50528 66688
rect 46992 66648 46998 66660
rect 50522 66648 50528 66660
rect 50580 66648 50586 66700
rect 51626 66648 51632 66700
rect 51684 66688 51690 66700
rect 53466 66688 53472 66700
rect 51684 66660 53472 66688
rect 51684 66648 51690 66660
rect 53466 66648 53472 66660
rect 53524 66648 53530 66700
rect 61304 66688 61332 66784
rect 63126 66716 63132 66768
rect 63184 66716 63190 66768
rect 61381 66691 61439 66697
rect 61381 66688 61393 66691
rect 61304 66660 61393 66688
rect 61381 66657 61393 66660
rect 61427 66657 61439 66691
rect 61381 66651 61439 66657
rect 71777 66691 71835 66697
rect 71777 66657 71789 66691
rect 71823 66688 71835 66691
rect 73724 66688 73752 66784
rect 71823 66660 73752 66688
rect 71823 66657 71835 66660
rect 71777 66651 71835 66657
rect 53484 66620 53512 66648
rect 55398 66620 55404 66632
rect 53484 66592 55404 66620
rect 55398 66580 55404 66592
rect 55456 66620 55462 66632
rect 55456 66592 55536 66620
rect 55456 66580 55462 66592
rect 49694 66512 49700 66564
rect 49752 66552 49758 66564
rect 51905 66555 51963 66561
rect 51905 66552 51917 66555
rect 49752 66524 51917 66552
rect 49752 66512 49758 66524
rect 51905 66521 51917 66524
rect 51951 66521 51963 66555
rect 55306 66552 55312 66564
rect 53130 66524 55312 66552
rect 51905 66515 51963 66521
rect 55306 66512 55312 66524
rect 55364 66512 55370 66564
rect 55508 66493 55536 66592
rect 61654 66512 61660 66564
rect 61712 66512 61718 66564
rect 64874 66552 64880 66564
rect 62882 66524 64880 66552
rect 64874 66512 64880 66524
rect 64932 66512 64938 66564
rect 71222 66512 71228 66564
rect 71280 66552 71286 66564
rect 72053 66555 72111 66561
rect 72053 66552 72065 66555
rect 71280 66524 72065 66552
rect 71280 66512 71286 66524
rect 72053 66521 72065 66524
rect 72099 66521 72111 66555
rect 73430 66552 73436 66564
rect 73278 66524 73436 66552
rect 72053 66515 72111 66521
rect 73430 66512 73436 66524
rect 73488 66512 73494 66564
rect 55493 66487 55551 66493
rect 55493 66453 55505 66487
rect 55539 66484 55551 66487
rect 56594 66484 56600 66496
rect 55539 66456 56600 66484
rect 55539 66453 55551 66456
rect 55493 66447 55551 66453
rect 56594 66444 56600 66456
rect 56652 66444 56658 66496
rect 73525 66487 73583 66493
rect 73525 66453 73537 66487
rect 73571 66484 73583 66487
rect 74166 66484 74172 66496
rect 73571 66456 74172 66484
rect 73571 66453 73583 66456
rect 73525 66447 73583 66453
rect 74166 66444 74172 66456
rect 74224 66444 74230 66496
rect 1104 66394 110860 66416
rect 1104 66342 4874 66394
rect 4926 66342 4938 66394
rect 4990 66342 5002 66394
rect 5054 66342 5066 66394
rect 5118 66342 5130 66394
rect 5182 66342 35594 66394
rect 35646 66342 35658 66394
rect 35710 66342 35722 66394
rect 35774 66342 35786 66394
rect 35838 66342 35850 66394
rect 35902 66342 66314 66394
rect 66366 66342 66378 66394
rect 66430 66342 66442 66394
rect 66494 66342 66506 66394
rect 66558 66342 66570 66394
rect 66622 66342 97034 66394
rect 97086 66342 97098 66394
rect 97150 66342 97162 66394
rect 97214 66342 97226 66394
rect 97278 66342 97290 66394
rect 97342 66342 107762 66394
rect 107814 66342 107826 66394
rect 107878 66342 107890 66394
rect 107942 66342 107954 66394
rect 108006 66342 108018 66394
rect 108070 66342 110860 66394
rect 1104 66320 110860 66342
rect 49142 66240 49148 66292
rect 49200 66280 49206 66292
rect 56413 66283 56471 66289
rect 49200 66252 52500 66280
rect 49200 66240 49206 66252
rect 48682 66172 48688 66224
rect 48740 66172 48746 66224
rect 50522 66172 50528 66224
rect 50580 66172 50586 66224
rect 52472 66221 52500 66252
rect 56413 66249 56425 66283
rect 56459 66280 56471 66283
rect 56594 66280 56600 66292
rect 56459 66252 56600 66280
rect 56459 66249 56471 66252
rect 56413 66243 56471 66249
rect 56594 66240 56600 66252
rect 56652 66280 56658 66292
rect 57882 66280 57888 66292
rect 56652 66252 57888 66280
rect 56652 66240 56658 66252
rect 57882 66240 57888 66252
rect 57940 66280 57946 66292
rect 59722 66280 59728 66292
rect 57940 66252 59728 66280
rect 57940 66240 57946 66252
rect 52457 66215 52515 66221
rect 52457 66181 52469 66215
rect 52503 66181 52515 66215
rect 52457 66175 52515 66181
rect 53926 66172 53932 66224
rect 53984 66212 53990 66224
rect 54021 66215 54079 66221
rect 54021 66212 54033 66215
rect 53984 66184 54033 66212
rect 53984 66172 53990 66184
rect 54021 66181 54033 66184
rect 54067 66181 54079 66215
rect 54021 66175 54079 66181
rect 55306 66172 55312 66224
rect 55364 66212 55370 66224
rect 58452 66221 58480 66252
rect 59722 66240 59728 66252
rect 59780 66240 59786 66292
rect 75549 66283 75607 66289
rect 75549 66249 75561 66283
rect 75595 66249 75607 66283
rect 75549 66243 75607 66249
rect 55677 66215 55735 66221
rect 55677 66212 55689 66215
rect 55364 66184 55689 66212
rect 55364 66172 55370 66184
rect 55677 66181 55689 66184
rect 55723 66181 55735 66215
rect 58437 66215 58495 66221
rect 55677 66175 55735 66181
rect 55784 66184 58112 66212
rect 55784 66153 55812 66184
rect 48777 66147 48835 66153
rect 48777 66113 48789 66147
rect 48823 66144 48835 66147
rect 50617 66147 50675 66153
rect 50617 66144 50629 66147
rect 48823 66116 50629 66144
rect 48823 66113 48835 66116
rect 48777 66107 48835 66113
rect 50617 66113 50629 66116
rect 50663 66144 50675 66147
rect 52549 66147 52607 66153
rect 52549 66144 52561 66147
rect 50663 66116 52561 66144
rect 50663 66113 50675 66116
rect 50617 66107 50675 66113
rect 52549 66113 52561 66116
rect 52595 66144 52607 66147
rect 54113 66147 54171 66153
rect 54113 66144 54125 66147
rect 52595 66116 54125 66144
rect 52595 66113 52607 66116
rect 52549 66107 52607 66113
rect 54113 66113 54125 66116
rect 54159 66144 54171 66147
rect 55769 66147 55827 66153
rect 55769 66144 55781 66147
rect 54159 66116 55781 66144
rect 54159 66113 54171 66116
rect 54113 66107 54171 66113
rect 55769 66113 55781 66116
rect 55815 66113 55827 66147
rect 55769 66107 55827 66113
rect 57701 66147 57759 66153
rect 57701 66113 57713 66147
rect 57747 66113 57759 66147
rect 57701 66107 57759 66113
rect 57716 66076 57744 66107
rect 57974 66104 57980 66156
rect 58032 66104 58038 66156
rect 58084 66153 58112 66184
rect 58437 66181 58449 66215
rect 58483 66181 58495 66215
rect 58437 66175 58495 66181
rect 60826 66172 60832 66224
rect 60884 66172 60890 66224
rect 60936 66184 63264 66212
rect 60936 66153 60964 66184
rect 63236 66153 63264 66184
rect 64432 66184 64828 66212
rect 64432 66153 64460 66184
rect 58069 66147 58127 66153
rect 58069 66113 58081 66147
rect 58115 66144 58127 66147
rect 59081 66147 59139 66153
rect 59081 66144 59093 66147
rect 58115 66116 59093 66144
rect 58115 66113 58127 66116
rect 58069 66107 58127 66113
rect 59081 66113 59093 66116
rect 59127 66144 59139 66147
rect 60921 66147 60979 66153
rect 60921 66144 60933 66147
rect 59127 66116 60933 66144
rect 59127 66113 59139 66116
rect 59081 66107 59139 66113
rect 60921 66113 60933 66116
rect 60967 66113 60979 66147
rect 60921 66107 60979 66113
rect 62853 66147 62911 66153
rect 62853 66113 62865 66147
rect 62899 66113 62911 66147
rect 62853 66107 62911 66113
rect 63221 66147 63279 66153
rect 63221 66113 63233 66147
rect 63267 66144 63279 66147
rect 64417 66147 64475 66153
rect 64417 66144 64429 66147
rect 63267 66116 64429 66144
rect 63267 66113 63279 66116
rect 63221 66107 63279 66113
rect 64417 66113 64429 66116
rect 64463 66113 64475 66147
rect 64417 66107 64475 66113
rect 62868 66076 62896 66107
rect 64598 66104 64604 66156
rect 64656 66144 64662 66156
rect 64800 66153 64828 66184
rect 64874 66172 64880 66224
rect 64932 66172 64938 66224
rect 66162 66172 66168 66224
rect 66220 66212 66226 66224
rect 66257 66215 66315 66221
rect 66257 66212 66269 66215
rect 66220 66184 66269 66212
rect 66220 66172 66226 66184
rect 66257 66181 66269 66184
rect 66303 66181 66315 66215
rect 66257 66175 66315 66181
rect 67542 66172 67548 66224
rect 67600 66212 67606 66224
rect 67913 66215 67971 66221
rect 67913 66212 67925 66215
rect 67600 66184 67925 66212
rect 67600 66172 67606 66184
rect 67913 66181 67925 66184
rect 67959 66181 67971 66215
rect 67913 66175 67971 66181
rect 69566 66172 69572 66224
rect 69624 66172 69630 66224
rect 71406 66172 71412 66224
rect 71464 66172 71470 66224
rect 73430 66172 73436 66224
rect 73488 66172 73494 66224
rect 75564 66212 75592 66243
rect 75730 66240 75736 66292
rect 75788 66240 75794 66292
rect 73540 66184 75592 66212
rect 75748 66212 75776 66240
rect 76009 66215 76067 66221
rect 76009 66212 76021 66215
rect 75748 66184 76021 66212
rect 73540 66153 73568 66184
rect 64693 66147 64751 66153
rect 64693 66144 64705 66147
rect 64656 66116 64705 66144
rect 64656 66104 64662 66116
rect 64693 66113 64705 66116
rect 64739 66113 64751 66147
rect 64693 66107 64751 66113
rect 64785 66147 64843 66153
rect 64785 66113 64797 66147
rect 64831 66113 64843 66147
rect 64785 66107 64843 66113
rect 66349 66147 66407 66153
rect 66349 66113 66361 66147
rect 66395 66144 66407 66147
rect 68005 66147 68063 66153
rect 68005 66144 68017 66147
rect 66395 66116 68017 66144
rect 66395 66113 66407 66116
rect 66349 66107 66407 66113
rect 68005 66113 68017 66116
rect 68051 66144 68063 66147
rect 69661 66147 69719 66153
rect 69661 66144 69673 66147
rect 68051 66116 69673 66144
rect 68051 66113 68063 66116
rect 68005 66107 68063 66113
rect 69661 66113 69673 66116
rect 69707 66144 69719 66147
rect 71501 66147 71559 66153
rect 71501 66144 71513 66147
rect 69707 66116 71513 66144
rect 69707 66113 69719 66116
rect 69661 66107 69719 66113
rect 71501 66113 71513 66116
rect 71547 66144 71559 66147
rect 73525 66147 73583 66153
rect 73525 66144 73537 66147
rect 71547 66116 73537 66144
rect 71547 66113 71559 66116
rect 71501 66107 71559 66113
rect 73525 66113 73537 66116
rect 73571 66113 73583 66147
rect 73525 66107 73583 66113
rect 75564 66076 75592 66184
rect 76009 66181 76021 66184
rect 76055 66181 76067 66215
rect 76009 66175 76067 66181
rect 95878 66172 95884 66224
rect 95936 66172 95942 66224
rect 75730 66104 75736 66156
rect 75788 66104 75794 66156
rect 75917 66147 75975 66153
rect 75917 66113 75929 66147
rect 75963 66113 75975 66147
rect 91925 66147 91983 66153
rect 91925 66144 91937 66147
rect 75917 66107 75975 66113
rect 76024 66116 76420 66144
rect 75932 66076 75960 66107
rect 57716 66048 58296 66076
rect 62868 66048 63632 66076
rect 58268 66017 58296 66048
rect 63604 66017 63632 66048
rect 64892 66048 70394 66076
rect 75564 66048 75960 66076
rect 58253 66011 58311 66017
rect 58253 65977 58265 66011
rect 58299 66008 58311 66011
rect 61565 66011 61623 66017
rect 61565 66008 61577 66011
rect 58299 65980 61577 66008
rect 58299 65977 58311 65980
rect 58253 65971 58311 65977
rect 61565 65977 61577 65980
rect 61611 66008 61623 66011
rect 63589 66011 63647 66017
rect 61611 65980 63448 66008
rect 61611 65977 61623 65980
rect 61565 65971 61623 65977
rect 63420 65952 63448 65980
rect 63589 65977 63601 66011
rect 63635 66008 63647 66011
rect 64892 66008 64920 66048
rect 63635 65980 64920 66008
rect 70366 66008 70394 66048
rect 76024 66008 76052 66116
rect 70366 65980 76052 66008
rect 63635 65977 63647 65980
rect 63589 65971 63647 65977
rect 57790 65900 57796 65952
rect 57848 65940 57854 65952
rect 58989 65943 59047 65949
rect 58989 65940 59001 65943
rect 57848 65912 59001 65940
rect 57848 65900 57854 65912
rect 58989 65909 59001 65912
rect 59035 65909 59047 65943
rect 58989 65903 59047 65909
rect 62022 65900 62028 65952
rect 62080 65940 62086 65952
rect 63129 65943 63187 65949
rect 63129 65940 63141 65943
rect 62080 65912 63141 65940
rect 62080 65900 62086 65912
rect 63129 65909 63141 65912
rect 63175 65909 63187 65943
rect 63129 65903 63187 65909
rect 63402 65900 63408 65952
rect 63460 65900 63466 65952
rect 64598 65900 64604 65952
rect 64656 65940 64662 65952
rect 65153 65943 65211 65949
rect 65153 65940 65165 65943
rect 64656 65912 65165 65940
rect 64656 65900 64662 65912
rect 65153 65909 65165 65912
rect 65199 65940 65211 65943
rect 75730 65940 75736 65952
rect 65199 65912 75736 65940
rect 65199 65909 65211 65912
rect 65153 65903 65211 65909
rect 75730 65900 75736 65912
rect 75788 65940 75794 65952
rect 76193 65943 76251 65949
rect 76193 65940 76205 65943
rect 75788 65912 76205 65940
rect 75788 65900 75794 65912
rect 76193 65909 76205 65912
rect 76239 65940 76251 65943
rect 76282 65940 76288 65952
rect 76239 65912 76288 65940
rect 76239 65909 76251 65912
rect 76193 65903 76251 65909
rect 76282 65900 76288 65912
rect 76340 65900 76346 65952
rect 76392 65940 76420 66116
rect 84166 66116 91937 66144
rect 76466 66036 76472 66088
rect 76524 66076 76530 66088
rect 84166 66076 84194 66116
rect 91925 66113 91937 66116
rect 91971 66144 91983 66147
rect 92382 66144 92388 66156
rect 91971 66116 92388 66144
rect 91971 66113 91983 66116
rect 91925 66107 91983 66113
rect 92382 66104 92388 66116
rect 92440 66104 92446 66156
rect 76524 66048 77294 66076
rect 76524 66036 76530 66048
rect 77266 66008 77294 66048
rect 80026 66048 84194 66076
rect 80026 66008 80054 66048
rect 102778 66008 102784 66020
rect 77266 65980 80054 66008
rect 82096 65980 102784 66008
rect 82096 65940 82124 65980
rect 102778 65968 102784 65980
rect 102836 65968 102842 66020
rect 76392 65912 82124 65940
rect 86310 65900 86316 65952
rect 86368 65900 86374 65952
rect 87322 65900 87328 65952
rect 87380 65900 87386 65952
rect 92017 65943 92075 65949
rect 92017 65909 92029 65943
rect 92063 65940 92075 65943
rect 92290 65940 92296 65952
rect 92063 65912 92296 65940
rect 92063 65909 92075 65912
rect 92017 65903 92075 65909
rect 92290 65900 92296 65912
rect 92348 65900 92354 65952
rect 1104 65850 110860 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 96374 65850
rect 96426 65798 96438 65850
rect 96490 65798 96502 65850
rect 96554 65798 96566 65850
rect 96618 65798 96630 65850
rect 96682 65798 107026 65850
rect 107078 65798 107090 65850
rect 107142 65798 107154 65850
rect 107206 65798 107218 65850
rect 107270 65798 107282 65850
rect 107334 65798 110860 65850
rect 1104 65776 110860 65798
rect 63402 65696 63408 65748
rect 63460 65736 63466 65748
rect 100754 65736 100760 65748
rect 63460 65708 100760 65736
rect 63460 65696 63466 65708
rect 100754 65696 100760 65708
rect 100812 65696 100818 65748
rect 92290 65628 92296 65680
rect 92348 65668 92354 65680
rect 102962 65668 102968 65680
rect 92348 65640 102968 65668
rect 92348 65628 92354 65640
rect 102962 65628 102968 65640
rect 103020 65628 103026 65680
rect 1104 65306 7912 65328
rect 1104 65254 4874 65306
rect 4926 65254 4938 65306
rect 4990 65254 5002 65306
rect 5054 65254 5066 65306
rect 5118 65254 5130 65306
rect 5182 65254 7912 65306
rect 1104 65232 7912 65254
rect 104052 65306 110860 65328
rect 104052 65254 107762 65306
rect 107814 65254 107826 65306
rect 107878 65254 107890 65306
rect 107942 65254 107954 65306
rect 108006 65254 108018 65306
rect 108070 65254 110860 65306
rect 104052 65232 110860 65254
rect 92382 64880 92388 64932
rect 92440 64920 92446 64932
rect 102870 64920 102876 64932
rect 92440 64892 102876 64920
rect 92440 64880 92446 64892
rect 102870 64880 102876 64892
rect 102928 64880 102934 64932
rect 1104 64762 7912 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 7912 64762
rect 1104 64688 7912 64710
rect 104052 64762 110860 64784
rect 104052 64710 107026 64762
rect 107078 64710 107090 64762
rect 107142 64710 107154 64762
rect 107206 64710 107218 64762
rect 107270 64710 107282 64762
rect 107334 64710 110860 64762
rect 104052 64688 110860 64710
rect 100754 64268 100760 64320
rect 100812 64308 100818 64320
rect 104434 64308 104440 64320
rect 100812 64280 104440 64308
rect 100812 64268 100818 64280
rect 104434 64268 104440 64280
rect 104492 64268 104498 64320
rect 1104 64218 7912 64240
rect 1104 64166 4874 64218
rect 4926 64166 4938 64218
rect 4990 64166 5002 64218
rect 5054 64166 5066 64218
rect 5118 64166 5130 64218
rect 5182 64166 7912 64218
rect 1104 64144 7912 64166
rect 104052 64218 110860 64240
rect 104052 64166 107762 64218
rect 107814 64166 107826 64218
rect 107878 64166 107890 64218
rect 107942 64166 107954 64218
rect 108006 64166 108018 64218
rect 108070 64166 110860 64218
rect 104052 64144 110860 64166
rect 1104 63674 7912 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 7912 63674
rect 1104 63600 7912 63622
rect 104052 63674 110860 63696
rect 104052 63622 107026 63674
rect 107078 63622 107090 63674
rect 107142 63622 107154 63674
rect 107206 63622 107218 63674
rect 107270 63622 107282 63674
rect 107334 63622 110860 63674
rect 104052 63600 110860 63622
rect 1104 63130 7912 63152
rect 1104 63078 4874 63130
rect 4926 63078 4938 63130
rect 4990 63078 5002 63130
rect 5054 63078 5066 63130
rect 5118 63078 5130 63130
rect 5182 63078 7912 63130
rect 1104 63056 7912 63078
rect 104052 63130 110860 63152
rect 104052 63078 107762 63130
rect 107814 63078 107826 63130
rect 107878 63078 107890 63130
rect 107942 63078 107954 63130
rect 108006 63078 108018 63130
rect 108070 63078 110860 63130
rect 104052 63056 110860 63078
rect 1104 62586 7912 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 7912 62586
rect 1104 62512 7912 62534
rect 104052 62586 110860 62608
rect 104052 62534 107026 62586
rect 107078 62534 107090 62586
rect 107142 62534 107154 62586
rect 107206 62534 107218 62586
rect 107270 62534 107282 62586
rect 107334 62534 110860 62586
rect 104052 62512 110860 62534
rect 1104 62042 7912 62064
rect 1104 61990 4874 62042
rect 4926 61990 4938 62042
rect 4990 61990 5002 62042
rect 5054 61990 5066 62042
rect 5118 61990 5130 62042
rect 5182 61990 7912 62042
rect 1104 61968 7912 61990
rect 104052 62042 110860 62064
rect 104052 61990 107762 62042
rect 107814 61990 107826 62042
rect 107878 61990 107890 62042
rect 107942 61990 107954 62042
rect 108006 61990 108018 62042
rect 108070 61990 110860 62042
rect 104052 61968 110860 61990
rect 1104 61498 7912 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 7912 61498
rect 1104 61424 7912 61446
rect 104052 61498 110860 61520
rect 104052 61446 107026 61498
rect 107078 61446 107090 61498
rect 107142 61446 107154 61498
rect 107206 61446 107218 61498
rect 107270 61446 107282 61498
rect 107334 61446 110860 61498
rect 104052 61424 110860 61446
rect 1104 60954 7912 60976
rect 1104 60902 4874 60954
rect 4926 60902 4938 60954
rect 4990 60902 5002 60954
rect 5054 60902 5066 60954
rect 5118 60902 5130 60954
rect 5182 60902 7912 60954
rect 1104 60880 7912 60902
rect 104052 60954 110860 60976
rect 104052 60902 107762 60954
rect 107814 60902 107826 60954
rect 107878 60902 107890 60954
rect 107942 60902 107954 60954
rect 108006 60902 108018 60954
rect 108070 60902 110860 60954
rect 104052 60880 110860 60902
rect 1104 60410 7912 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 7912 60410
rect 1104 60336 7912 60358
rect 104052 60410 110860 60432
rect 104052 60358 107026 60410
rect 107078 60358 107090 60410
rect 107142 60358 107154 60410
rect 107206 60358 107218 60410
rect 107270 60358 107282 60410
rect 107334 60358 110860 60410
rect 104052 60336 110860 60358
rect 103698 60052 103704 60104
rect 103756 60092 103762 60104
rect 104345 60095 104403 60101
rect 104345 60092 104357 60095
rect 103756 60064 104357 60092
rect 103756 60052 103762 60064
rect 104345 60061 104357 60064
rect 104391 60061 104403 60095
rect 104345 60055 104403 60061
rect 1104 59866 7912 59888
rect 1104 59814 4874 59866
rect 4926 59814 4938 59866
rect 4990 59814 5002 59866
rect 5054 59814 5066 59866
rect 5118 59814 5130 59866
rect 5182 59814 7912 59866
rect 1104 59792 7912 59814
rect 104052 59866 110860 59888
rect 104052 59814 107762 59866
rect 107814 59814 107826 59866
rect 107878 59814 107890 59866
rect 107942 59814 107954 59866
rect 108006 59814 108018 59866
rect 108070 59814 110860 59866
rect 104052 59792 110860 59814
rect 1104 59322 7912 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 7912 59322
rect 1104 59248 7912 59270
rect 104052 59322 110860 59344
rect 104052 59270 107026 59322
rect 107078 59270 107090 59322
rect 107142 59270 107154 59322
rect 107206 59270 107218 59322
rect 107270 59270 107282 59322
rect 107334 59270 110860 59322
rect 104052 59248 110860 59270
rect 1104 58778 7912 58800
rect 1104 58726 4874 58778
rect 4926 58726 4938 58778
rect 4990 58726 5002 58778
rect 5054 58726 5066 58778
rect 5118 58726 5130 58778
rect 5182 58726 7912 58778
rect 1104 58704 7912 58726
rect 104052 58778 110860 58800
rect 104052 58726 107762 58778
rect 107814 58726 107826 58778
rect 107878 58726 107890 58778
rect 107942 58726 107954 58778
rect 108006 58726 108018 58778
rect 108070 58726 110860 58778
rect 104052 58704 110860 58726
rect 1104 58234 7912 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 7912 58234
rect 1104 58160 7912 58182
rect 104052 58234 110860 58256
rect 104052 58182 107026 58234
rect 107078 58182 107090 58234
rect 107142 58182 107154 58234
rect 107206 58182 107218 58234
rect 107270 58182 107282 58234
rect 107334 58182 110860 58234
rect 104052 58160 110860 58182
rect 102962 57876 102968 57928
rect 103020 57916 103026 57928
rect 103020 57888 103514 57916
rect 103020 57876 103026 57888
rect 103486 57780 103514 57888
rect 104345 57783 104403 57789
rect 104345 57780 104357 57783
rect 103486 57752 104357 57780
rect 1104 57690 7912 57712
rect 1104 57638 4874 57690
rect 4926 57638 4938 57690
rect 4990 57638 5002 57690
rect 5054 57638 5066 57690
rect 5118 57638 5130 57690
rect 5182 57638 7912 57690
rect 1104 57616 7912 57638
rect 103992 57508 104020 57752
rect 104345 57749 104357 57752
rect 104391 57749 104403 57783
rect 104345 57743 104403 57749
rect 104052 57690 110860 57712
rect 104052 57638 107762 57690
rect 107814 57638 107826 57690
rect 107878 57638 107890 57690
rect 107942 57638 107954 57690
rect 108006 57638 108018 57690
rect 108070 57638 110860 57690
rect 104052 57616 110860 57638
rect 103992 57480 105110 57508
rect 104342 57400 104348 57452
rect 104400 57400 104406 57452
rect 104618 57332 104624 57384
rect 104676 57332 104682 57384
rect 104986 57332 104992 57384
rect 105044 57372 105050 57384
rect 106369 57375 106427 57381
rect 106369 57372 106381 57375
rect 105044 57344 106381 57372
rect 105044 57332 105050 57344
rect 106369 57341 106381 57344
rect 106415 57372 106427 57375
rect 106461 57375 106519 57381
rect 106461 57372 106473 57375
rect 106415 57344 106473 57372
rect 106415 57341 106427 57344
rect 106369 57335 106427 57341
rect 106461 57341 106473 57344
rect 106507 57341 106519 57375
rect 106461 57335 106519 57341
rect 106642 57196 106648 57248
rect 106700 57196 106706 57248
rect 1104 57146 7912 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 7912 57146
rect 1104 57072 7912 57094
rect 104052 57146 110860 57168
rect 104052 57094 107026 57146
rect 107078 57094 107090 57146
rect 107142 57094 107154 57146
rect 107206 57094 107218 57146
rect 107270 57094 107282 57146
rect 107334 57094 110860 57146
rect 104052 57072 110860 57094
rect 104986 56856 104992 56908
rect 105044 56896 105050 56908
rect 105173 56899 105231 56905
rect 105173 56896 105185 56899
rect 105044 56868 105185 56896
rect 105044 56856 105050 56868
rect 105173 56865 105185 56868
rect 105219 56865 105231 56899
rect 105173 56859 105231 56865
rect 104437 56695 104495 56701
rect 104437 56661 104449 56695
rect 104483 56692 104495 56695
rect 104526 56692 104532 56704
rect 104483 56664 104532 56692
rect 104483 56661 104495 56664
rect 104437 56655 104495 56661
rect 104526 56652 104532 56664
rect 104584 56652 104590 56704
rect 1104 56602 7912 56624
rect 1104 56550 4874 56602
rect 4926 56550 4938 56602
rect 4990 56550 5002 56602
rect 5054 56550 5066 56602
rect 5118 56550 5130 56602
rect 5182 56550 7912 56602
rect 1104 56528 7912 56550
rect 104052 56602 110860 56624
rect 104052 56550 107762 56602
rect 107814 56550 107826 56602
rect 107878 56550 107890 56602
rect 107942 56550 107954 56602
rect 108006 56550 108018 56602
rect 108070 56550 110860 56602
rect 104052 56528 110860 56550
rect 1104 56058 7912 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 7912 56058
rect 1104 55984 7912 56006
rect 104052 56058 110860 56080
rect 104052 56006 107026 56058
rect 107078 56006 107090 56058
rect 107142 56006 107154 56058
rect 107206 56006 107218 56058
rect 107270 56006 107282 56058
rect 107334 56006 110860 56058
rect 104052 55984 110860 56006
rect 104437 55947 104495 55953
rect 104437 55913 104449 55947
rect 104483 55944 104495 55947
rect 104618 55944 104624 55956
rect 104483 55916 104624 55944
rect 104483 55913 104495 55916
rect 104437 55907 104495 55913
rect 104618 55904 104624 55916
rect 104676 55904 104682 55956
rect 104526 55700 104532 55752
rect 104584 55700 104590 55752
rect 1104 55514 7912 55536
rect 1104 55462 4874 55514
rect 4926 55462 4938 55514
rect 4990 55462 5002 55514
rect 5054 55462 5066 55514
rect 5118 55462 5130 55514
rect 5182 55462 7912 55514
rect 1104 55440 7912 55462
rect 104052 55514 110860 55536
rect 104052 55462 107762 55514
rect 107814 55462 107826 55514
rect 107878 55462 107890 55514
rect 107942 55462 107954 55514
rect 108006 55462 108018 55514
rect 108070 55462 110860 55514
rect 104052 55440 110860 55462
rect 1104 54970 7912 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 7912 54970
rect 1104 54896 7912 54918
rect 104052 54970 110860 54992
rect 104052 54918 107026 54970
rect 107078 54918 107090 54970
rect 107142 54918 107154 54970
rect 107206 54918 107218 54970
rect 107270 54918 107282 54970
rect 107334 54918 110860 54970
rect 104052 54896 110860 54918
rect 104250 54680 104256 54732
rect 104308 54720 104314 54732
rect 104345 54723 104403 54729
rect 104345 54720 104357 54723
rect 104308 54692 104357 54720
rect 104308 54680 104314 54692
rect 104345 54689 104357 54692
rect 104391 54720 104403 54723
rect 106366 54720 106372 54732
rect 104391 54692 106372 54720
rect 104391 54689 104403 54692
rect 104345 54683 104403 54689
rect 106366 54680 106372 54692
rect 106424 54720 106430 54732
rect 106737 54723 106795 54729
rect 106737 54720 106749 54723
rect 106424 54692 106749 54720
rect 106424 54680 106430 54692
rect 106737 54689 106749 54692
rect 106783 54689 106795 54723
rect 106737 54683 106795 54689
rect 104618 54544 104624 54596
rect 104676 54544 104682 54596
rect 105078 54544 105084 54596
rect 105136 54544 105142 54596
rect 106182 54544 106188 54596
rect 106240 54584 106246 54596
rect 106369 54587 106427 54593
rect 106369 54584 106381 54587
rect 106240 54556 106381 54584
rect 106240 54544 106246 54556
rect 106369 54553 106381 54556
rect 106415 54584 106427 54587
rect 106461 54587 106519 54593
rect 106461 54584 106473 54587
rect 106415 54556 106473 54584
rect 106415 54553 106427 54556
rect 106369 54547 106427 54553
rect 106461 54553 106473 54556
rect 106507 54553 106519 54587
rect 106461 54547 106519 54553
rect 1104 54426 7912 54448
rect 1104 54374 4874 54426
rect 4926 54374 4938 54426
rect 4990 54374 5002 54426
rect 5054 54374 5066 54426
rect 5118 54374 5130 54426
rect 5182 54374 7912 54426
rect 1104 54352 7912 54374
rect 104052 54426 110860 54448
rect 104052 54374 107762 54426
rect 107814 54374 107826 54426
rect 107878 54374 107890 54426
rect 107942 54374 107954 54426
rect 108006 54374 108018 54426
rect 108070 54374 110860 54426
rect 104052 54352 110860 54374
rect 104437 54315 104495 54321
rect 104437 54281 104449 54315
rect 104483 54312 104495 54315
rect 105078 54312 105084 54324
rect 104483 54284 105084 54312
rect 104483 54281 104495 54284
rect 104437 54275 104495 54281
rect 105078 54272 105084 54284
rect 105136 54272 105142 54324
rect 102870 54136 102876 54188
rect 102928 54176 102934 54188
rect 104345 54179 104403 54185
rect 104345 54176 104357 54179
rect 102928 54148 104357 54176
rect 102928 54136 102934 54148
rect 104345 54145 104357 54148
rect 104391 54176 104403 54179
rect 104526 54176 104532 54188
rect 104391 54148 104532 54176
rect 104391 54145 104403 54148
rect 104345 54139 104403 54145
rect 104526 54136 104532 54148
rect 104584 54136 104590 54188
rect 104526 53932 104532 53984
rect 104584 53972 104590 53984
rect 104621 53975 104679 53981
rect 104621 53972 104633 53975
rect 104584 53944 104633 53972
rect 104584 53932 104590 53944
rect 104621 53941 104633 53944
rect 104667 53941 104679 53975
rect 104621 53935 104679 53941
rect 1104 53882 7912 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 7912 53882
rect 1104 53808 7912 53830
rect 104052 53882 110860 53904
rect 104052 53830 107026 53882
rect 107078 53830 107090 53882
rect 107142 53830 107154 53882
rect 107206 53830 107218 53882
rect 107270 53830 107282 53882
rect 107334 53830 110860 53882
rect 104052 53808 110860 53830
rect 104345 53771 104403 53777
rect 104345 53737 104357 53771
rect 104391 53768 104403 53771
rect 104618 53768 104624 53780
rect 104391 53740 104624 53768
rect 104391 53737 104403 53740
rect 104345 53731 104403 53737
rect 104618 53728 104624 53740
rect 104676 53728 104682 53780
rect 104986 53728 104992 53780
rect 105044 53728 105050 53780
rect 104621 53635 104679 53641
rect 104621 53601 104633 53635
rect 104667 53632 104679 53635
rect 104894 53632 104900 53644
rect 104667 53604 104900 53632
rect 104667 53601 104679 53604
rect 104621 53595 104679 53601
rect 104894 53592 104900 53604
rect 104952 53632 104958 53644
rect 105173 53635 105231 53641
rect 105173 53632 105185 53635
rect 104952 53604 105185 53632
rect 104952 53592 104958 53604
rect 105173 53601 105185 53604
rect 105219 53632 105231 53635
rect 106182 53632 106188 53644
rect 105219 53604 106188 53632
rect 105219 53601 105231 53604
rect 105173 53595 105231 53601
rect 106182 53592 106188 53604
rect 106240 53592 106246 53644
rect 104713 53567 104771 53573
rect 104713 53533 104725 53567
rect 104759 53564 104771 53567
rect 104802 53564 104808 53576
rect 104759 53536 104808 53564
rect 104759 53533 104771 53536
rect 104713 53527 104771 53533
rect 104802 53524 104808 53536
rect 104860 53564 104866 53576
rect 104986 53564 104992 53576
rect 104860 53536 104992 53564
rect 104860 53524 104866 53536
rect 104986 53524 104992 53536
rect 105044 53524 105050 53576
rect 1104 53338 7912 53360
rect 1104 53286 4874 53338
rect 4926 53286 4938 53338
rect 4990 53286 5002 53338
rect 5054 53286 5066 53338
rect 5118 53286 5130 53338
rect 5182 53286 7912 53338
rect 1104 53264 7912 53286
rect 104052 53338 110860 53360
rect 104052 53286 107762 53338
rect 107814 53286 107826 53338
rect 107878 53286 107890 53338
rect 107942 53286 107954 53338
rect 108006 53286 108018 53338
rect 108070 53286 110860 53338
rect 104052 53264 110860 53286
rect 1104 52794 7912 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 7912 52794
rect 1104 52720 7912 52742
rect 104052 52794 110860 52816
rect 104052 52742 107026 52794
rect 107078 52742 107090 52794
rect 107142 52742 107154 52794
rect 107206 52742 107218 52794
rect 107270 52742 107282 52794
rect 107334 52742 110860 52794
rect 104052 52720 110860 52742
rect 1104 52250 7912 52272
rect 1104 52198 4874 52250
rect 4926 52198 4938 52250
rect 4990 52198 5002 52250
rect 5054 52198 5066 52250
rect 5118 52198 5130 52250
rect 5182 52198 7912 52250
rect 1104 52176 7912 52198
rect 104052 52250 110860 52272
rect 104052 52198 107762 52250
rect 107814 52198 107826 52250
rect 107878 52198 107890 52250
rect 107942 52198 107954 52250
rect 108006 52198 108018 52250
rect 108070 52198 110860 52250
rect 104052 52176 110860 52198
rect 1104 51706 7912 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 7912 51706
rect 1104 51632 7912 51654
rect 104052 51706 110860 51728
rect 104052 51654 107026 51706
rect 107078 51654 107090 51706
rect 107142 51654 107154 51706
rect 107206 51654 107218 51706
rect 107270 51654 107282 51706
rect 107334 51654 110860 51706
rect 104052 51632 110860 51654
rect 1104 51162 7912 51184
rect 1104 51110 4874 51162
rect 4926 51110 4938 51162
rect 4990 51110 5002 51162
rect 5054 51110 5066 51162
rect 5118 51110 5130 51162
rect 5182 51110 7912 51162
rect 1104 51088 7912 51110
rect 104052 51162 110860 51184
rect 104052 51110 107762 51162
rect 107814 51110 107826 51162
rect 107878 51110 107890 51162
rect 107942 51110 107954 51162
rect 108006 51110 108018 51162
rect 108070 51110 110860 51162
rect 104052 51088 110860 51110
rect 1104 50618 7912 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 7912 50618
rect 1104 50544 7912 50566
rect 104052 50618 110860 50640
rect 104052 50566 107026 50618
rect 107078 50566 107090 50618
rect 107142 50566 107154 50618
rect 107206 50566 107218 50618
rect 107270 50566 107282 50618
rect 107334 50566 110860 50618
rect 104052 50544 110860 50566
rect 1104 50074 7912 50096
rect 1104 50022 4874 50074
rect 4926 50022 4938 50074
rect 4990 50022 5002 50074
rect 5054 50022 5066 50074
rect 5118 50022 5130 50074
rect 5182 50022 7912 50074
rect 1104 50000 7912 50022
rect 104052 50074 110860 50096
rect 104052 50022 107762 50074
rect 107814 50022 107826 50074
rect 107878 50022 107890 50074
rect 107942 50022 107954 50074
rect 108006 50022 108018 50074
rect 108070 50022 110860 50074
rect 104052 50000 110860 50022
rect 1104 49530 7912 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 7912 49530
rect 1104 49456 7912 49478
rect 104052 49530 110860 49552
rect 104052 49478 107026 49530
rect 107078 49478 107090 49530
rect 107142 49478 107154 49530
rect 107206 49478 107218 49530
rect 107270 49478 107282 49530
rect 107334 49478 110860 49530
rect 104052 49456 110860 49478
rect 1104 48986 7912 49008
rect 1104 48934 4874 48986
rect 4926 48934 4938 48986
rect 4990 48934 5002 48986
rect 5054 48934 5066 48986
rect 5118 48934 5130 48986
rect 5182 48934 7912 48986
rect 1104 48912 7912 48934
rect 104052 48986 110860 49008
rect 104052 48934 107762 48986
rect 107814 48934 107826 48986
rect 107878 48934 107890 48986
rect 107942 48934 107954 48986
rect 108006 48934 108018 48986
rect 108070 48934 110860 48986
rect 104052 48912 110860 48934
rect 1104 48442 7912 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 7912 48442
rect 1104 48368 7912 48390
rect 104052 48442 110860 48464
rect 104052 48390 107026 48442
rect 107078 48390 107090 48442
rect 107142 48390 107154 48442
rect 107206 48390 107218 48442
rect 107270 48390 107282 48442
rect 107334 48390 110860 48442
rect 104052 48368 110860 48390
rect 1104 47898 7912 47920
rect 1104 47846 4874 47898
rect 4926 47846 4938 47898
rect 4990 47846 5002 47898
rect 5054 47846 5066 47898
rect 5118 47846 5130 47898
rect 5182 47846 7912 47898
rect 1104 47824 7912 47846
rect 104052 47898 110860 47920
rect 104052 47846 107762 47898
rect 107814 47846 107826 47898
rect 107878 47846 107890 47898
rect 107942 47846 107954 47898
rect 108006 47846 108018 47898
rect 108070 47846 110860 47898
rect 104052 47824 110860 47846
rect 1104 47354 7912 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 7912 47354
rect 1104 47280 7912 47302
rect 104052 47354 110860 47376
rect 104052 47302 107026 47354
rect 107078 47302 107090 47354
rect 107142 47302 107154 47354
rect 107206 47302 107218 47354
rect 107270 47302 107282 47354
rect 107334 47302 110860 47354
rect 104052 47280 110860 47302
rect 1104 46810 7912 46832
rect 1104 46758 4874 46810
rect 4926 46758 4938 46810
rect 4990 46758 5002 46810
rect 5054 46758 5066 46810
rect 5118 46758 5130 46810
rect 5182 46758 7912 46810
rect 1104 46736 7912 46758
rect 104052 46810 110860 46832
rect 104052 46758 107762 46810
rect 107814 46758 107826 46810
rect 107878 46758 107890 46810
rect 107942 46758 107954 46810
rect 108006 46758 108018 46810
rect 108070 46758 110860 46810
rect 104052 46736 110860 46758
rect 1104 46266 7912 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 7912 46266
rect 1104 46192 7912 46214
rect 104052 46266 110860 46288
rect 104052 46214 107026 46266
rect 107078 46214 107090 46266
rect 107142 46214 107154 46266
rect 107206 46214 107218 46266
rect 107270 46214 107282 46266
rect 107334 46214 110860 46266
rect 104052 46192 110860 46214
rect 104802 46152 104808 46164
rect 104544 46124 104808 46152
rect 104250 46044 104256 46096
rect 104308 46084 104314 46096
rect 104345 46087 104403 46093
rect 104345 46084 104357 46087
rect 104308 46056 104357 46084
rect 104308 46044 104314 46056
rect 104345 46053 104357 46056
rect 104391 46053 104403 46087
rect 104345 46047 104403 46053
rect 104544 45957 104572 46124
rect 104802 46112 104808 46124
rect 104860 46112 104866 46164
rect 104529 45951 104587 45957
rect 104529 45917 104541 45951
rect 104575 45917 104587 45951
rect 104529 45911 104587 45917
rect 104621 45951 104679 45957
rect 104621 45917 104633 45951
rect 104667 45948 104679 45951
rect 104894 45948 104900 45960
rect 104667 45920 104900 45948
rect 104667 45917 104679 45920
rect 104621 45911 104679 45917
rect 104894 45908 104900 45920
rect 104952 45908 104958 45960
rect 104345 45883 104403 45889
rect 104345 45849 104357 45883
rect 104391 45880 104403 45883
rect 104391 45852 105216 45880
rect 104391 45849 104403 45852
rect 104345 45843 104403 45849
rect 104894 45772 104900 45824
rect 104952 45772 104958 45824
rect 105188 45821 105216 45852
rect 105173 45815 105231 45821
rect 105173 45781 105185 45815
rect 105219 45812 105231 45815
rect 105446 45812 105452 45824
rect 105219 45784 105452 45812
rect 105219 45781 105231 45784
rect 105173 45775 105231 45781
rect 105446 45772 105452 45784
rect 105504 45772 105510 45824
rect 1104 45722 7912 45744
rect 1104 45670 4874 45722
rect 4926 45670 4938 45722
rect 4990 45670 5002 45722
rect 5054 45670 5066 45722
rect 5118 45670 5130 45722
rect 5182 45670 7912 45722
rect 1104 45648 7912 45670
rect 104052 45722 110860 45744
rect 104052 45670 107762 45722
rect 107814 45670 107826 45722
rect 107878 45670 107890 45722
rect 107942 45670 107954 45722
rect 108006 45670 108018 45722
rect 108070 45670 110860 45722
rect 104052 45648 110860 45670
rect 1104 45178 7912 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 7912 45178
rect 1104 45104 7912 45126
rect 104052 45178 110860 45200
rect 104052 45126 107026 45178
rect 107078 45126 107090 45178
rect 107142 45126 107154 45178
rect 107206 45126 107218 45178
rect 107270 45126 107282 45178
rect 107334 45126 110860 45178
rect 104052 45104 110860 45126
rect 104529 45067 104587 45073
rect 104529 45033 104541 45067
rect 104575 45064 104587 45067
rect 104894 45064 104900 45076
rect 104575 45036 104900 45064
rect 104575 45033 104587 45036
rect 104529 45027 104587 45033
rect 104894 45024 104900 45036
rect 104952 45064 104958 45076
rect 105265 45067 105323 45073
rect 105265 45064 105277 45067
rect 104952 45036 105277 45064
rect 104952 45024 104958 45036
rect 105265 45033 105277 45036
rect 105311 45033 105323 45067
rect 105265 45027 105323 45033
rect 104710 44996 104716 45008
rect 104544 44968 104716 44996
rect 104345 44795 104403 44801
rect 104345 44761 104357 44795
rect 104391 44792 104403 44795
rect 104544 44792 104572 44968
rect 104710 44956 104716 44968
rect 104768 44996 104774 45008
rect 105081 44999 105139 45005
rect 105081 44996 105093 44999
rect 104768 44968 105093 44996
rect 104768 44956 104774 44968
rect 105081 44965 105093 44968
rect 105127 44965 105139 44999
rect 105081 44959 105139 44965
rect 105446 44928 105452 44940
rect 104391 44764 104572 44792
rect 104636 44900 105452 44928
rect 104391 44761 104403 44764
rect 104345 44755 104403 44761
rect 104529 44727 104587 44733
rect 104529 44693 104541 44727
rect 104575 44724 104587 44727
rect 104636 44724 104664 44900
rect 105446 44888 105452 44900
rect 105504 44888 105510 44940
rect 104575 44696 104664 44724
rect 104713 44727 104771 44733
rect 104575 44693 104587 44696
rect 104529 44687 104587 44693
rect 104713 44693 104725 44727
rect 104759 44724 104771 44727
rect 104897 44727 104955 44733
rect 104897 44724 104909 44727
rect 104759 44696 104909 44724
rect 104759 44693 104771 44696
rect 104713 44687 104771 44693
rect 104897 44693 104909 44696
rect 104943 44724 104955 44727
rect 105170 44724 105176 44736
rect 104943 44696 105176 44724
rect 104943 44693 104955 44696
rect 104897 44687 104955 44693
rect 105170 44684 105176 44696
rect 105228 44684 105234 44736
rect 105446 44684 105452 44736
rect 105504 44684 105510 44736
rect 1104 44634 7912 44656
rect 1104 44582 4874 44634
rect 4926 44582 4938 44634
rect 4990 44582 5002 44634
rect 5054 44582 5066 44634
rect 5118 44582 5130 44634
rect 5182 44582 7912 44634
rect 1104 44560 7912 44582
rect 104052 44634 110860 44656
rect 104052 44582 107762 44634
rect 107814 44582 107826 44634
rect 107878 44582 107890 44634
rect 107942 44582 107954 44634
rect 108006 44582 108018 44634
rect 108070 44582 110860 44634
rect 104052 44560 110860 44582
rect 1104 44090 7912 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 7912 44090
rect 1104 44016 7912 44038
rect 104052 44090 110860 44112
rect 104052 44038 107026 44090
rect 107078 44038 107090 44090
rect 107142 44038 107154 44090
rect 107206 44038 107218 44090
rect 107270 44038 107282 44090
rect 107334 44038 110860 44090
rect 104052 44016 110860 44038
rect 104526 43936 104532 43988
rect 104584 43976 104590 43988
rect 104621 43979 104679 43985
rect 104621 43976 104633 43979
rect 104584 43948 104633 43976
rect 104584 43936 104590 43948
rect 104621 43945 104633 43948
rect 104667 43945 104679 43979
rect 104621 43939 104679 43945
rect 104345 43775 104403 43781
rect 104345 43741 104357 43775
rect 104391 43772 104403 43775
rect 104526 43772 104532 43784
rect 104391 43744 104532 43772
rect 104391 43741 104403 43744
rect 104345 43735 104403 43741
rect 104526 43732 104532 43744
rect 104584 43732 104590 43784
rect 104437 43707 104495 43713
rect 104437 43673 104449 43707
rect 104483 43704 104495 43707
rect 105078 43704 105084 43716
rect 104483 43676 105084 43704
rect 104483 43673 104495 43676
rect 104437 43667 104495 43673
rect 105078 43664 105084 43676
rect 105136 43664 105142 43716
rect 1104 43546 7912 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 7912 43546
rect 1104 43472 7912 43494
rect 104052 43546 110860 43568
rect 104052 43494 107762 43546
rect 107814 43494 107826 43546
rect 107878 43494 107890 43546
rect 107942 43494 107954 43546
rect 108006 43494 108018 43546
rect 108070 43494 110860 43546
rect 104052 43472 110860 43494
rect 1104 43002 7912 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 7912 43002
rect 1104 42928 7912 42950
rect 104052 43002 110860 43024
rect 104052 42950 107026 43002
rect 107078 42950 107090 43002
rect 107142 42950 107154 43002
rect 107206 42950 107218 43002
rect 107270 42950 107282 43002
rect 107334 42950 110860 43002
rect 104052 42928 110860 42950
rect 104345 42755 104403 42761
rect 104345 42721 104357 42755
rect 104391 42752 104403 42755
rect 104986 42752 104992 42764
rect 104391 42724 104992 42752
rect 104391 42721 104403 42724
rect 104345 42715 104403 42721
rect 104986 42712 104992 42724
rect 105044 42712 105050 42764
rect 104618 42576 104624 42628
rect 104676 42576 104682 42628
rect 105078 42576 105084 42628
rect 105136 42576 105142 42628
rect 104158 42508 104164 42560
rect 104216 42548 104222 42560
rect 105446 42548 105452 42560
rect 104216 42520 105452 42548
rect 104216 42508 104222 42520
rect 105446 42508 105452 42520
rect 105504 42548 105510 42560
rect 106093 42551 106151 42557
rect 106093 42548 106105 42551
rect 105504 42520 106105 42548
rect 105504 42508 105510 42520
rect 106093 42517 106105 42520
rect 106139 42548 106151 42551
rect 106185 42551 106243 42557
rect 106185 42548 106197 42551
rect 106139 42520 106197 42548
rect 106139 42517 106151 42520
rect 106093 42511 106151 42517
rect 106185 42517 106197 42520
rect 106231 42517 106243 42551
rect 106185 42511 106243 42517
rect 106366 42508 106372 42560
rect 106424 42508 106430 42560
rect 1104 42458 7912 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 7912 42458
rect 1104 42384 7912 42406
rect 104052 42458 110860 42480
rect 104052 42406 107762 42458
rect 107814 42406 107826 42458
rect 107878 42406 107890 42458
rect 107942 42406 107954 42458
rect 108006 42406 108018 42458
rect 108070 42406 110860 42458
rect 104052 42384 110860 42406
rect 104529 42211 104587 42217
rect 104529 42177 104541 42211
rect 104575 42208 104587 42211
rect 104986 42208 104992 42220
rect 104575 42180 104992 42208
rect 104575 42177 104587 42180
rect 104529 42171 104587 42177
rect 104986 42168 104992 42180
rect 105044 42208 105050 42220
rect 106090 42208 106096 42220
rect 105044 42180 106096 42208
rect 105044 42168 105050 42180
rect 106090 42168 106096 42180
rect 106148 42168 106154 42220
rect 106090 41964 106096 42016
rect 106148 42004 106154 42016
rect 106366 42004 106372 42016
rect 106148 41976 106372 42004
rect 106148 41964 106154 41976
rect 106366 41964 106372 41976
rect 106424 42004 106430 42016
rect 106553 42007 106611 42013
rect 106553 42004 106565 42007
rect 106424 41976 106565 42004
rect 106424 41964 106430 41976
rect 106553 41973 106565 41976
rect 106599 41973 106611 42007
rect 106553 41967 106611 41973
rect 1104 41914 7912 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 7912 41914
rect 1104 41840 7912 41862
rect 104052 41914 110860 41936
rect 104052 41862 107026 41914
rect 107078 41862 107090 41914
rect 107142 41862 107154 41914
rect 107206 41862 107218 41914
rect 107270 41862 107282 41914
rect 107334 41862 110860 41914
rect 104052 41840 110860 41862
rect 104342 41556 104348 41608
rect 104400 41596 104406 41608
rect 104894 41596 104900 41608
rect 104400 41568 104900 41596
rect 104400 41556 104406 41568
rect 104894 41556 104900 41568
rect 104952 41556 104958 41608
rect 106090 41488 106096 41540
rect 106148 41528 106154 41540
rect 106185 41531 106243 41537
rect 106185 41528 106197 41531
rect 106148 41500 106197 41528
rect 106148 41488 106154 41500
rect 106185 41497 106197 41500
rect 106231 41497 106243 41531
rect 106185 41491 106243 41497
rect 7558 41420 7564 41472
rect 7616 41420 7622 41472
rect 1104 41370 7912 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 7912 41370
rect 1104 41296 7912 41318
rect 104052 41370 110860 41392
rect 104052 41318 107762 41370
rect 107814 41318 107826 41370
rect 107878 41318 107890 41370
rect 107942 41318 107954 41370
rect 108006 41318 108018 41370
rect 108070 41318 110860 41370
rect 104052 41296 110860 41318
rect 104437 41259 104495 41265
rect 104437 41225 104449 41259
rect 104483 41256 104495 41259
rect 104618 41256 104624 41268
rect 104483 41228 104624 41256
rect 104483 41225 104495 41228
rect 104437 41219 104495 41225
rect 104618 41216 104624 41228
rect 104676 41216 104682 41268
rect 104894 41216 104900 41268
rect 104952 41216 104958 41268
rect 104250 41080 104256 41132
rect 104308 41120 104314 41132
rect 104345 41123 104403 41129
rect 104345 41120 104357 41123
rect 104308 41092 104357 41120
rect 104308 41080 104314 41092
rect 104345 41089 104357 41092
rect 104391 41089 104403 41123
rect 104345 41083 104403 41089
rect 104529 41123 104587 41129
rect 104529 41089 104541 41123
rect 104575 41120 104587 41123
rect 104575 41092 104756 41120
rect 104575 41089 104587 41092
rect 104529 41083 104587 41089
rect 104728 40925 104756 41092
rect 104713 40919 104771 40925
rect 104713 40885 104725 40919
rect 104759 40916 104771 40919
rect 105170 40916 105176 40928
rect 104759 40888 105176 40916
rect 104759 40885 104771 40888
rect 104713 40879 104771 40885
rect 105170 40876 105176 40888
rect 105228 40916 105234 40928
rect 105906 40916 105912 40928
rect 105228 40888 105912 40916
rect 105228 40876 105234 40888
rect 105906 40876 105912 40888
rect 105964 40876 105970 40928
rect 1104 40826 7912 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 7912 40826
rect 1104 40752 7912 40774
rect 104052 40826 110860 40848
rect 104052 40774 107026 40826
rect 107078 40774 107090 40826
rect 107142 40774 107154 40826
rect 107206 40774 107218 40826
rect 107270 40774 107282 40826
rect 107334 40774 110860 40826
rect 104052 40752 110860 40774
rect 1104 40282 7912 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 7912 40282
rect 1104 40208 7912 40230
rect 104052 40282 110860 40304
rect 104052 40230 107762 40282
rect 107814 40230 107826 40282
rect 107878 40230 107890 40282
rect 107942 40230 107954 40282
rect 108006 40230 108018 40282
rect 108070 40230 110860 40282
rect 104052 40208 110860 40230
rect 7558 39788 7564 39840
rect 7616 39788 7622 39840
rect 1104 39738 7912 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 7912 39738
rect 1104 39664 7912 39686
rect 104052 39738 110860 39760
rect 104052 39686 107026 39738
rect 107078 39686 107090 39738
rect 107142 39686 107154 39738
rect 107206 39686 107218 39738
rect 107270 39686 107282 39738
rect 107334 39686 110860 39738
rect 104052 39664 110860 39686
rect 1104 39194 7912 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 7912 39194
rect 1104 39120 7912 39142
rect 104052 39194 110860 39216
rect 104052 39142 107762 39194
rect 107814 39142 107826 39194
rect 107878 39142 107890 39194
rect 107942 39142 107954 39194
rect 108006 39142 108018 39194
rect 108070 39142 110860 39194
rect 104052 39120 110860 39142
rect 7558 38700 7564 38752
rect 7616 38700 7622 38752
rect 1104 38650 7912 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 7912 38650
rect 1104 38576 7912 38598
rect 104052 38650 110860 38672
rect 104052 38598 107026 38650
rect 107078 38598 107090 38650
rect 107142 38598 107154 38650
rect 107206 38598 107218 38650
rect 107270 38598 107282 38650
rect 107334 38598 110860 38650
rect 104052 38576 110860 38598
rect 1104 38106 7912 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 7912 38106
rect 1104 38032 7912 38054
rect 104052 38106 110860 38128
rect 104052 38054 107762 38106
rect 107814 38054 107826 38106
rect 107878 38054 107890 38106
rect 107942 38054 107954 38106
rect 108006 38054 108018 38106
rect 108070 38054 110860 38106
rect 104052 38032 110860 38054
rect 1104 37562 7912 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 7912 37562
rect 1104 37488 7912 37510
rect 104052 37562 110860 37584
rect 104052 37510 107026 37562
rect 107078 37510 107090 37562
rect 107142 37510 107154 37562
rect 107206 37510 107218 37562
rect 107270 37510 107282 37562
rect 107334 37510 110860 37562
rect 104052 37488 110860 37510
rect 1104 37018 7912 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 7912 37018
rect 1104 36944 7912 36966
rect 104052 37018 110860 37040
rect 104052 36966 107762 37018
rect 107814 36966 107826 37018
rect 107878 36966 107890 37018
rect 107942 36966 107954 37018
rect 108006 36966 108018 37018
rect 108070 36966 110860 37018
rect 104052 36944 110860 36966
rect 104526 36864 104532 36916
rect 104584 36904 104590 36916
rect 104621 36907 104679 36913
rect 104621 36904 104633 36907
rect 104584 36876 104633 36904
rect 104584 36864 104590 36876
rect 104621 36873 104633 36876
rect 104667 36873 104679 36907
rect 104621 36867 104679 36873
rect 7558 36728 7564 36780
rect 7616 36728 7622 36780
rect 104345 36771 104403 36777
rect 104345 36737 104357 36771
rect 104391 36768 104403 36771
rect 104544 36768 104572 36864
rect 104391 36740 104572 36768
rect 104391 36737 104403 36740
rect 104345 36731 104403 36737
rect 104437 36567 104495 36573
rect 104437 36533 104449 36567
rect 104483 36564 104495 36567
rect 104526 36564 104532 36576
rect 104483 36536 104532 36564
rect 104483 36533 104495 36536
rect 104437 36527 104495 36533
rect 104526 36524 104532 36536
rect 104584 36524 104590 36576
rect 1104 36474 7912 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 7912 36474
rect 1104 36400 7912 36422
rect 104052 36474 110860 36496
rect 104052 36422 107026 36474
rect 107078 36422 107090 36474
rect 107142 36422 107154 36474
rect 107206 36422 107218 36474
rect 107270 36422 107282 36474
rect 107334 36422 110860 36474
rect 104052 36400 110860 36422
rect 1104 35930 7912 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 7912 35930
rect 1104 35856 7912 35878
rect 104052 35930 110860 35952
rect 104052 35878 107762 35930
rect 107814 35878 107826 35930
rect 107878 35878 107890 35930
rect 107942 35878 107954 35930
rect 108006 35878 108018 35930
rect 108070 35878 110860 35930
rect 104052 35856 110860 35878
rect 104345 35683 104403 35689
rect 104345 35649 104357 35683
rect 104391 35680 104403 35683
rect 104710 35680 104716 35692
rect 104391 35652 104716 35680
rect 104391 35649 104403 35652
rect 104345 35643 104403 35649
rect 104710 35640 104716 35652
rect 104768 35640 104774 35692
rect 7558 35504 7564 35556
rect 7616 35504 7622 35556
rect 104434 35436 104440 35488
rect 104492 35436 104498 35488
rect 104710 35436 104716 35488
rect 104768 35436 104774 35488
rect 1104 35386 7912 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 7912 35386
rect 1104 35312 7912 35334
rect 104052 35386 110860 35408
rect 104052 35334 107026 35386
rect 107078 35334 107090 35386
rect 107142 35334 107154 35386
rect 107206 35334 107218 35386
rect 107270 35334 107282 35386
rect 107334 35334 110860 35386
rect 104052 35312 110860 35334
rect 1104 34842 7912 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 7912 34842
rect 1104 34768 7912 34790
rect 104052 34842 110860 34864
rect 104052 34790 107762 34842
rect 107814 34790 107826 34842
rect 107878 34790 107890 34842
rect 107942 34790 107954 34842
rect 108006 34790 108018 34842
rect 108070 34790 110860 34842
rect 104052 34768 110860 34790
rect 1104 34298 7912 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 7912 34298
rect 1104 34224 7912 34246
rect 104052 34298 110860 34320
rect 104052 34246 107026 34298
rect 107078 34246 107090 34298
rect 107142 34246 107154 34298
rect 107206 34246 107218 34298
rect 107270 34246 107282 34298
rect 107334 34246 110860 34298
rect 104052 34224 110860 34246
rect 7558 34008 7564 34060
rect 7616 34008 7622 34060
rect 106090 33940 106096 33992
rect 106148 33980 106154 33992
rect 106148 33952 106228 33980
rect 106148 33940 106154 33952
rect 104526 33872 104532 33924
rect 104584 33912 104590 33924
rect 104584 33884 104650 33912
rect 104584 33872 104590 33884
rect 105814 33872 105820 33924
rect 105872 33872 105878 33924
rect 106200 33856 106228 33952
rect 104345 33847 104403 33853
rect 104345 33813 104357 33847
rect 104391 33844 104403 33847
rect 104802 33844 104808 33856
rect 104391 33816 104808 33844
rect 104391 33813 104403 33816
rect 104345 33807 104403 33813
rect 104802 33804 104808 33816
rect 104860 33804 104866 33856
rect 106182 33804 106188 33856
rect 106240 33804 106246 33856
rect 1104 33754 7912 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 7912 33754
rect 1104 33680 7912 33702
rect 104052 33754 110860 33776
rect 104052 33702 107762 33754
rect 107814 33702 107826 33754
rect 107878 33702 107890 33754
rect 107942 33702 107954 33754
rect 108006 33702 108018 33754
rect 108070 33702 110860 33754
rect 104052 33680 110860 33702
rect 104802 33396 104808 33448
rect 104860 33396 104866 33448
rect 105357 33303 105415 33309
rect 105357 33269 105369 33303
rect 105403 33300 105415 33303
rect 105630 33300 105636 33312
rect 105403 33272 105636 33300
rect 105403 33269 105415 33272
rect 105357 33263 105415 33269
rect 105630 33260 105636 33272
rect 105688 33260 105694 33312
rect 1104 33210 7912 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 7912 33210
rect 1104 33136 7912 33158
rect 104052 33210 110860 33232
rect 104052 33158 107026 33210
rect 107078 33158 107090 33210
rect 107142 33158 107154 33210
rect 107206 33158 107218 33210
rect 107270 33158 107282 33210
rect 107334 33158 110860 33210
rect 104052 33136 110860 33158
rect 105446 32920 105452 32972
rect 105504 32960 105510 32972
rect 105817 32963 105875 32969
rect 105817 32960 105829 32963
rect 105504 32932 105829 32960
rect 105504 32920 105510 32932
rect 105817 32929 105829 32932
rect 105863 32929 105875 32963
rect 105817 32923 105875 32929
rect 106093 32895 106151 32901
rect 106093 32861 106105 32895
rect 106139 32892 106151 32895
rect 106182 32892 106188 32904
rect 106139 32864 106188 32892
rect 106139 32861 106151 32864
rect 106093 32855 106151 32861
rect 106182 32852 106188 32864
rect 106240 32892 106246 32904
rect 106240 32864 106320 32892
rect 106240 32852 106246 32864
rect 104434 32784 104440 32836
rect 104492 32824 104498 32836
rect 104492 32796 104650 32824
rect 104492 32784 104498 32796
rect 104345 32759 104403 32765
rect 104345 32725 104357 32759
rect 104391 32756 104403 32759
rect 104526 32756 104532 32768
rect 104391 32728 104532 32756
rect 104391 32725 104403 32728
rect 104345 32719 104403 32725
rect 104526 32716 104532 32728
rect 104584 32716 104590 32768
rect 106292 32765 106320 32864
rect 106277 32759 106335 32765
rect 106277 32725 106289 32759
rect 106323 32756 106335 32759
rect 106366 32756 106372 32768
rect 106323 32728 106372 32756
rect 106323 32725 106335 32728
rect 106277 32719 106335 32725
rect 106366 32716 106372 32728
rect 106424 32716 106430 32768
rect 1104 32666 7912 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 7912 32666
rect 1104 32592 7912 32614
rect 104052 32666 110860 32688
rect 104052 32614 107762 32666
rect 107814 32614 107826 32666
rect 107878 32614 107890 32666
rect 107942 32614 107954 32666
rect 108006 32614 108018 32666
rect 108070 32614 110860 32666
rect 104052 32592 110860 32614
rect 105265 32419 105323 32425
rect 105265 32385 105277 32419
rect 105311 32416 105323 32419
rect 110322 32416 110328 32428
rect 105311 32388 110328 32416
rect 105311 32385 105323 32388
rect 105265 32379 105323 32385
rect 110322 32376 110328 32388
rect 110380 32376 110386 32428
rect 104526 32308 104532 32360
rect 104584 32348 104590 32360
rect 104710 32348 104716 32360
rect 104584 32320 104716 32348
rect 104584 32308 104590 32320
rect 104710 32308 104716 32320
rect 104768 32348 104774 32360
rect 105357 32351 105415 32357
rect 105357 32348 105369 32351
rect 104768 32320 105369 32348
rect 104768 32308 104774 32320
rect 105357 32317 105369 32320
rect 105403 32317 105415 32351
rect 105357 32311 105415 32317
rect 1104 32122 7912 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 7912 32122
rect 1104 32048 7912 32070
rect 104052 32122 110860 32144
rect 104052 32070 107026 32122
rect 107078 32070 107090 32122
rect 107142 32070 107154 32122
rect 107206 32070 107218 32122
rect 107270 32070 107282 32122
rect 107334 32070 110860 32122
rect 104052 32048 110860 32070
rect 105814 31968 105820 32020
rect 105872 32008 105878 32020
rect 106001 32011 106059 32017
rect 106001 32008 106013 32011
rect 105872 31980 106013 32008
rect 105872 31968 105878 31980
rect 106001 31977 106013 31980
rect 106047 31977 106059 32011
rect 106001 31971 106059 31977
rect 110322 31968 110328 32020
rect 110380 31968 110386 32020
rect 104437 31943 104495 31949
rect 104437 31909 104449 31943
rect 104483 31940 104495 31943
rect 104710 31940 104716 31952
rect 104483 31912 104716 31940
rect 104483 31909 104495 31912
rect 104437 31903 104495 31909
rect 104710 31900 104716 31912
rect 104768 31900 104774 31952
rect 105906 31940 105912 31952
rect 105740 31912 105912 31940
rect 105740 31881 105768 31912
rect 105906 31900 105912 31912
rect 105964 31940 105970 31952
rect 106093 31943 106151 31949
rect 106093 31940 106105 31943
rect 105964 31912 106105 31940
rect 105964 31900 105970 31912
rect 106093 31909 106105 31912
rect 106139 31909 106151 31943
rect 106093 31903 106151 31909
rect 105725 31875 105783 31881
rect 105725 31841 105737 31875
rect 105771 31841 105783 31875
rect 105725 31835 105783 31841
rect 104345 31807 104403 31813
rect 104345 31773 104357 31807
rect 104391 31804 104403 31807
rect 104526 31804 104532 31816
rect 104391 31776 104532 31804
rect 104391 31773 104403 31776
rect 104345 31767 104403 31773
rect 104526 31764 104532 31776
rect 104584 31764 104590 31816
rect 104618 31764 104624 31816
rect 104676 31804 104682 31816
rect 104713 31807 104771 31813
rect 104713 31804 104725 31807
rect 104676 31776 104725 31804
rect 104676 31764 104682 31776
rect 104713 31773 104725 31776
rect 104759 31773 104771 31807
rect 104713 31767 104771 31773
rect 105354 31764 105360 31816
rect 105412 31764 105418 31816
rect 105630 31764 105636 31816
rect 105688 31764 105694 31816
rect 110233 31807 110291 31813
rect 110233 31773 110245 31807
rect 110279 31804 110291 31807
rect 110506 31804 110512 31816
rect 110279 31776 110512 31804
rect 110279 31773 110291 31776
rect 110233 31767 110291 31773
rect 110506 31764 110512 31776
rect 110564 31764 110570 31816
rect 1104 31578 7912 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 7912 31578
rect 1104 31504 7912 31526
rect 104052 31578 110860 31600
rect 104052 31526 107762 31578
rect 107814 31526 107826 31578
rect 107878 31526 107890 31578
rect 107942 31526 107954 31578
rect 108006 31526 108018 31578
rect 108070 31526 110860 31578
rect 104052 31504 110860 31526
rect 104526 31084 104532 31136
rect 104584 31124 104590 31136
rect 104621 31127 104679 31133
rect 104621 31124 104633 31127
rect 104584 31096 104633 31124
rect 104584 31084 104590 31096
rect 104621 31093 104633 31096
rect 104667 31093 104679 31127
rect 104621 31087 104679 31093
rect 1104 31034 7912 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 7912 31034
rect 1104 30960 7912 30982
rect 104052 31034 110860 31056
rect 104052 30982 107026 31034
rect 107078 30982 107090 31034
rect 107142 30982 107154 31034
rect 107206 30982 107218 31034
rect 107270 30982 107282 31034
rect 107334 30982 110860 31034
rect 104052 30960 110860 30982
rect 1104 30490 7912 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 7912 30490
rect 1104 30416 7912 30438
rect 104052 30490 110860 30512
rect 104052 30438 107762 30490
rect 107814 30438 107826 30490
rect 107878 30438 107890 30490
rect 107942 30438 107954 30490
rect 108006 30438 108018 30490
rect 108070 30438 110860 30490
rect 104052 30416 110860 30438
rect 104434 30268 104440 30320
rect 104492 30308 104498 30320
rect 104802 30308 104808 30320
rect 104492 30280 104808 30308
rect 104492 30268 104498 30280
rect 104802 30268 104808 30280
rect 104860 30308 104866 30320
rect 105817 30311 105875 30317
rect 104860 30280 105492 30308
rect 104860 30268 104866 30280
rect 104989 30243 105047 30249
rect 104989 30209 105001 30243
rect 105035 30240 105047 30243
rect 105354 30240 105360 30252
rect 105035 30212 105360 30240
rect 105035 30209 105047 30212
rect 104989 30203 105047 30209
rect 105354 30200 105360 30212
rect 105412 30200 105418 30252
rect 105464 30249 105492 30280
rect 105817 30277 105829 30311
rect 105863 30308 105875 30311
rect 105906 30308 105912 30320
rect 105863 30280 105912 30308
rect 105863 30277 105875 30280
rect 105817 30271 105875 30277
rect 105449 30243 105507 30249
rect 105449 30209 105461 30243
rect 105495 30209 105507 30243
rect 105449 30203 105507 30209
rect 105633 30243 105691 30249
rect 105633 30209 105645 30243
rect 105679 30240 105691 30243
rect 105832 30240 105860 30271
rect 105906 30268 105912 30280
rect 105964 30268 105970 30320
rect 105679 30212 105860 30240
rect 105679 30209 105691 30212
rect 105633 30203 105691 30209
rect 105081 30175 105139 30181
rect 105081 30141 105093 30175
rect 105127 30172 105139 30175
rect 105541 30175 105599 30181
rect 105541 30172 105553 30175
rect 105127 30144 105553 30172
rect 105127 30141 105139 30144
rect 105081 30135 105139 30141
rect 105541 30141 105553 30144
rect 105587 30141 105599 30175
rect 105541 30135 105599 30141
rect 105357 30107 105415 30113
rect 105357 30073 105369 30107
rect 105403 30104 105415 30107
rect 105446 30104 105452 30116
rect 105403 30076 105452 30104
rect 105403 30073 105415 30076
rect 105357 30067 105415 30073
rect 105446 30064 105452 30076
rect 105504 30064 105510 30116
rect 1104 29946 7912 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 7912 29946
rect 1104 29872 7912 29894
rect 104052 29946 110860 29968
rect 104052 29894 107026 29946
rect 107078 29894 107090 29946
rect 107142 29894 107154 29946
rect 107206 29894 107218 29946
rect 107270 29894 107282 29946
rect 107334 29894 110860 29946
rect 104052 29872 110860 29894
rect 104345 29631 104403 29637
rect 104345 29597 104357 29631
rect 104391 29628 104403 29631
rect 104526 29628 104532 29640
rect 104391 29600 104532 29628
rect 104391 29597 104403 29600
rect 104345 29591 104403 29597
rect 104526 29588 104532 29600
rect 104584 29628 104590 29640
rect 104584 29600 104756 29628
rect 104584 29588 104590 29600
rect 104250 29452 104256 29504
rect 104308 29492 104314 29504
rect 104728 29501 104756 29600
rect 104437 29495 104495 29501
rect 104437 29492 104449 29495
rect 104308 29464 104449 29492
rect 104308 29452 104314 29464
rect 104437 29461 104449 29464
rect 104483 29461 104495 29495
rect 104437 29455 104495 29461
rect 104713 29495 104771 29501
rect 104713 29461 104725 29495
rect 104759 29492 104771 29495
rect 104802 29492 104808 29504
rect 104759 29464 104808 29492
rect 104759 29461 104771 29464
rect 104713 29455 104771 29461
rect 104802 29452 104808 29464
rect 104860 29452 104866 29504
rect 1104 29402 7912 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 7912 29402
rect 1104 29328 7912 29350
rect 104052 29402 110860 29424
rect 104052 29350 107762 29402
rect 107814 29350 107826 29402
rect 107878 29350 107890 29402
rect 107942 29350 107954 29402
rect 108006 29350 108018 29402
rect 108070 29350 110860 29402
rect 104052 29328 110860 29350
rect 1104 28858 7912 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 7912 28858
rect 1104 28784 7912 28806
rect 104052 28858 110860 28880
rect 104052 28806 107026 28858
rect 107078 28806 107090 28858
rect 107142 28806 107154 28858
rect 107206 28806 107218 28858
rect 107270 28806 107282 28858
rect 107334 28806 110860 28858
rect 104052 28784 110860 28806
rect 104345 28611 104403 28617
rect 104345 28577 104357 28611
rect 104391 28608 104403 28611
rect 106366 28608 106372 28620
rect 104391 28580 106372 28608
rect 104391 28577 104403 28580
rect 104345 28571 104403 28577
rect 106366 28568 106372 28580
rect 106424 28568 106430 28620
rect 104526 28432 104532 28484
rect 104584 28472 104590 28484
rect 104621 28475 104679 28481
rect 104621 28472 104633 28475
rect 104584 28444 104633 28472
rect 104584 28432 104590 28444
rect 104621 28441 104633 28444
rect 104667 28441 104679 28475
rect 104621 28435 104679 28441
rect 104710 28432 104716 28484
rect 104768 28472 104774 28484
rect 104768 28444 105110 28472
rect 104768 28432 104774 28444
rect 105446 28364 105452 28416
rect 105504 28404 105510 28416
rect 106093 28407 106151 28413
rect 106093 28404 106105 28407
rect 105504 28376 106105 28404
rect 105504 28364 105510 28376
rect 106093 28373 106105 28376
rect 106139 28404 106151 28407
rect 106277 28407 106335 28413
rect 106277 28404 106289 28407
rect 106139 28376 106289 28404
rect 106139 28373 106151 28376
rect 106093 28367 106151 28373
rect 106277 28373 106289 28376
rect 106323 28373 106335 28407
rect 106277 28367 106335 28373
rect 106366 28364 106372 28416
rect 106424 28404 106430 28416
rect 106461 28407 106519 28413
rect 106461 28404 106473 28407
rect 106424 28376 106473 28404
rect 106424 28364 106430 28376
rect 106461 28373 106473 28376
rect 106507 28373 106519 28407
rect 106461 28367 106519 28373
rect 1104 28314 7912 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 7912 28314
rect 1104 28240 7912 28262
rect 104052 28314 110860 28336
rect 104052 28262 107762 28314
rect 107814 28262 107826 28314
rect 107878 28262 107890 28314
rect 107942 28262 107954 28314
rect 108006 28262 108018 28314
rect 108070 28262 110860 28314
rect 104052 28240 110860 28262
rect 104713 28203 104771 28209
rect 104713 28169 104725 28203
rect 104759 28200 104771 28203
rect 104759 28172 105032 28200
rect 104759 28169 104771 28172
rect 104713 28163 104771 28169
rect 104434 28092 104440 28144
rect 104492 28132 104498 28144
rect 105004 28141 105032 28172
rect 105078 28141 105084 28144
rect 104805 28135 104863 28141
rect 104805 28132 104817 28135
rect 104492 28104 104817 28132
rect 104492 28092 104498 28104
rect 104805 28101 104817 28104
rect 104851 28101 104863 28135
rect 105004 28135 105084 28141
rect 105004 28104 105033 28135
rect 104805 28095 104863 28101
rect 105021 28101 105033 28104
rect 105067 28101 105084 28135
rect 105021 28095 105084 28101
rect 105078 28092 105084 28095
rect 105136 28132 105142 28144
rect 105906 28132 105912 28144
rect 105136 28104 105912 28132
rect 105136 28092 105142 28104
rect 105906 28092 105912 28104
rect 105964 28092 105970 28144
rect 104710 27820 104716 27872
rect 104768 27860 104774 27872
rect 104989 27863 105047 27869
rect 104989 27860 105001 27863
rect 104768 27832 105001 27860
rect 104768 27820 104774 27832
rect 104989 27829 105001 27832
rect 105035 27829 105047 27863
rect 104989 27823 105047 27829
rect 105170 27820 105176 27872
rect 105228 27820 105234 27872
rect 1104 27770 7912 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 7912 27770
rect 1104 27696 7912 27718
rect 104052 27770 110860 27792
rect 104052 27718 107026 27770
rect 107078 27718 107090 27770
rect 107142 27718 107154 27770
rect 107206 27718 107218 27770
rect 107270 27718 107282 27770
rect 107334 27718 110860 27770
rect 104052 27696 110860 27718
rect 1104 27226 7912 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 7912 27226
rect 1104 27152 7912 27174
rect 104052 27226 110860 27248
rect 104052 27174 107762 27226
rect 107814 27174 107826 27226
rect 107878 27174 107890 27226
rect 107942 27174 107954 27226
rect 108006 27174 108018 27226
rect 108070 27174 110860 27226
rect 104052 27152 110860 27174
rect 104437 27115 104495 27121
rect 104437 27081 104449 27115
rect 104483 27112 104495 27115
rect 104526 27112 104532 27124
rect 104483 27084 104532 27112
rect 104483 27081 104495 27084
rect 104437 27075 104495 27081
rect 104526 27072 104532 27084
rect 104584 27072 104590 27124
rect 104621 27115 104679 27121
rect 104621 27081 104633 27115
rect 104667 27112 104679 27115
rect 104710 27112 104716 27124
rect 104667 27084 104716 27112
rect 104667 27081 104679 27084
rect 104621 27075 104679 27081
rect 104710 27072 104716 27084
rect 104768 27072 104774 27124
rect 105078 27112 105084 27124
rect 104912 27084 105084 27112
rect 104618 26979 104676 26985
rect 104618 26945 104630 26979
rect 104664 26976 104676 26979
rect 104912 26976 104940 27084
rect 105078 27072 105084 27084
rect 105136 27112 105142 27124
rect 105173 27115 105231 27121
rect 105173 27112 105185 27115
rect 105136 27084 105185 27112
rect 105136 27072 105142 27084
rect 105173 27081 105185 27084
rect 105219 27081 105231 27115
rect 105173 27075 105231 27081
rect 105446 27072 105452 27124
rect 105504 27072 105510 27124
rect 105262 27044 105268 27056
rect 105004 27016 105268 27044
rect 105004 26985 105032 27016
rect 105262 27004 105268 27016
rect 105320 27044 105326 27056
rect 105464 27044 105492 27072
rect 105320 27016 105492 27044
rect 105320 27004 105326 27016
rect 104664 26948 104940 26976
rect 104989 26979 105047 26985
rect 104664 26945 104676 26948
rect 104618 26939 104676 26945
rect 104989 26945 105001 26979
rect 105035 26945 105047 26979
rect 104989 26939 105047 26945
rect 105081 26979 105139 26985
rect 105081 26945 105093 26979
rect 105127 26976 105139 26979
rect 105170 26976 105176 26988
rect 105127 26948 105176 26976
rect 105127 26945 105139 26948
rect 105081 26939 105139 26945
rect 105170 26936 105176 26948
rect 105228 26936 105234 26988
rect 1104 26682 7912 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 7912 26682
rect 1104 26608 7912 26630
rect 104052 26682 110860 26704
rect 104052 26630 107026 26682
rect 107078 26630 107090 26682
rect 107142 26630 107154 26682
rect 107206 26630 107218 26682
rect 107270 26630 107282 26682
rect 107334 26630 110860 26682
rect 104052 26608 110860 26630
rect 104342 26256 104348 26308
rect 104400 26296 104406 26308
rect 106366 26296 106372 26308
rect 104400 26268 106372 26296
rect 104400 26256 104406 26268
rect 106366 26256 106372 26268
rect 106424 26256 106430 26308
rect 1104 26138 7912 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 7912 26138
rect 1104 26064 7912 26086
rect 104052 26138 110860 26160
rect 104052 26086 107762 26138
rect 107814 26086 107826 26138
rect 107878 26086 107890 26138
rect 107942 26086 107954 26138
rect 108006 26086 108018 26138
rect 108070 26086 110860 26138
rect 104052 26064 110860 26086
rect 104250 25916 104256 25968
rect 104308 25956 104314 25968
rect 104308 25928 105110 25956
rect 104308 25916 104314 25928
rect 104342 25848 104348 25900
rect 104400 25848 104406 25900
rect 104618 25780 104624 25832
rect 104676 25780 104682 25832
rect 105262 25644 105268 25696
rect 105320 25684 105326 25696
rect 106093 25687 106151 25693
rect 106093 25684 106105 25687
rect 105320 25656 106105 25684
rect 105320 25644 105326 25656
rect 106093 25653 106105 25656
rect 106139 25684 106151 25687
rect 106185 25687 106243 25693
rect 106185 25684 106197 25687
rect 106139 25656 106197 25684
rect 106139 25653 106151 25656
rect 106093 25647 106151 25653
rect 106185 25653 106197 25656
rect 106231 25653 106243 25687
rect 106185 25647 106243 25653
rect 106366 25644 106372 25696
rect 106424 25644 106430 25696
rect 1104 25594 7912 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 7912 25594
rect 1104 25520 7912 25542
rect 104052 25594 110860 25616
rect 104052 25542 107026 25594
rect 107078 25542 107090 25594
rect 107142 25542 107154 25594
rect 107206 25542 107218 25594
rect 107270 25542 107282 25594
rect 107334 25542 110860 25594
rect 104052 25520 110860 25542
rect 104526 25440 104532 25492
rect 104584 25440 104590 25492
rect 104710 25440 104716 25492
rect 104768 25440 104774 25492
rect 104802 25236 104808 25288
rect 104860 25276 104866 25288
rect 105081 25279 105139 25285
rect 105081 25276 105093 25279
rect 104860 25248 105093 25276
rect 104860 25236 104866 25248
rect 105081 25245 105093 25248
rect 105127 25245 105139 25279
rect 105081 25239 105139 25245
rect 104342 25168 104348 25220
rect 104400 25168 104406 25220
rect 105170 25208 105176 25220
rect 104820 25180 105176 25208
rect 104250 25100 104256 25152
rect 104308 25140 104314 25152
rect 104545 25143 104603 25149
rect 104545 25140 104557 25143
rect 104308 25112 104557 25140
rect 104308 25100 104314 25112
rect 104545 25109 104557 25112
rect 104591 25140 104603 25143
rect 104820 25140 104848 25180
rect 105170 25168 105176 25180
rect 105228 25208 105234 25220
rect 105265 25211 105323 25217
rect 105265 25208 105277 25211
rect 105228 25180 105277 25208
rect 105228 25168 105234 25180
rect 105265 25177 105277 25180
rect 105311 25177 105323 25211
rect 105265 25171 105323 25177
rect 104591 25112 104848 25140
rect 104591 25109 104603 25112
rect 104545 25103 104603 25109
rect 104894 25100 104900 25152
rect 104952 25100 104958 25152
rect 1104 25050 7912 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 7912 25050
rect 1104 24976 7912 24998
rect 104052 25050 110860 25072
rect 104052 24998 107762 25050
rect 107814 24998 107826 25050
rect 107878 24998 107890 25050
rect 107942 24998 107954 25050
rect 108006 24998 108018 25050
rect 108070 24998 110860 25050
rect 104052 24976 110860 24998
rect 104158 24760 104164 24812
rect 104216 24800 104222 24812
rect 104345 24803 104403 24809
rect 104345 24800 104357 24803
rect 104216 24772 104357 24800
rect 104216 24760 104222 24772
rect 104345 24769 104357 24772
rect 104391 24769 104403 24803
rect 104345 24763 104403 24769
rect 1104 24506 7912 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 7912 24506
rect 1104 24432 7912 24454
rect 104052 24506 110860 24528
rect 104052 24454 107026 24506
rect 107078 24454 107090 24506
rect 107142 24454 107154 24506
rect 107206 24454 107218 24506
rect 107270 24454 107282 24506
rect 107334 24454 110860 24506
rect 104052 24432 110860 24454
rect 104805 24395 104863 24401
rect 104805 24361 104817 24395
rect 104851 24392 104863 24395
rect 104986 24392 104992 24404
rect 104851 24364 104992 24392
rect 104851 24361 104863 24364
rect 104805 24355 104863 24361
rect 104820 24256 104848 24355
rect 104986 24352 104992 24364
rect 105044 24352 105050 24404
rect 104544 24228 104848 24256
rect 104544 24197 104572 24228
rect 104529 24191 104587 24197
rect 104529 24157 104541 24191
rect 104575 24157 104587 24191
rect 104529 24151 104587 24157
rect 104621 24191 104679 24197
rect 104621 24157 104633 24191
rect 104667 24188 104679 24191
rect 104710 24188 104716 24200
rect 104667 24160 104716 24188
rect 104667 24157 104679 24160
rect 104621 24151 104679 24157
rect 104710 24148 104716 24160
rect 104768 24148 104774 24200
rect 104158 24080 104164 24132
rect 104216 24120 104222 24132
rect 104345 24123 104403 24129
rect 104345 24120 104357 24123
rect 104216 24092 104357 24120
rect 104216 24080 104222 24092
rect 104345 24089 104357 24092
rect 104391 24120 104403 24123
rect 104897 24123 104955 24129
rect 104897 24120 104909 24123
rect 104391 24092 104909 24120
rect 104391 24089 104403 24092
rect 104345 24083 104403 24089
rect 104897 24089 104909 24092
rect 104943 24120 104955 24123
rect 105262 24120 105268 24132
rect 104943 24092 105268 24120
rect 104943 24089 104955 24092
rect 104897 24083 104955 24089
rect 105262 24080 105268 24092
rect 105320 24080 105326 24132
rect 104434 24012 104440 24064
rect 104492 24061 104498 24064
rect 104492 24015 104501 24061
rect 104492 24012 104498 24015
rect 1104 23962 7912 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 7912 23962
rect 1104 23888 7912 23910
rect 104052 23962 110860 23984
rect 104052 23910 107762 23962
rect 107814 23910 107826 23962
rect 107878 23910 107890 23962
rect 107942 23910 107954 23962
rect 108006 23910 108018 23962
rect 108070 23910 110860 23962
rect 104052 23888 110860 23910
rect 104555 23851 104613 23857
rect 104555 23817 104567 23851
rect 104601 23848 104613 23851
rect 104710 23848 104716 23860
rect 104601 23820 104716 23848
rect 104601 23817 104613 23820
rect 104555 23811 104613 23817
rect 104710 23808 104716 23820
rect 104768 23808 104774 23860
rect 104986 23808 104992 23860
rect 105044 23848 105050 23860
rect 105081 23851 105139 23857
rect 105081 23848 105093 23851
rect 105044 23820 105093 23848
rect 105044 23808 105050 23820
rect 105081 23817 105093 23820
rect 105127 23817 105139 23851
rect 105081 23811 105139 23817
rect 105262 23808 105268 23860
rect 105320 23808 105326 23860
rect 104158 23740 104164 23792
rect 104216 23780 104222 23792
rect 104345 23783 104403 23789
rect 104345 23780 104357 23783
rect 104216 23752 104357 23780
rect 104216 23740 104222 23752
rect 104345 23749 104357 23752
rect 104391 23749 104403 23783
rect 105004 23780 105032 23808
rect 104345 23743 104403 23749
rect 104912 23752 105032 23780
rect 104434 23672 104440 23724
rect 104492 23712 104498 23724
rect 104805 23715 104863 23721
rect 104805 23712 104817 23715
rect 104492 23684 104817 23712
rect 104492 23672 104498 23684
rect 104805 23681 104817 23684
rect 104851 23681 104863 23715
rect 104805 23675 104863 23681
rect 104912 23644 104940 23752
rect 104989 23715 105047 23721
rect 104989 23681 105001 23715
rect 105035 23681 105047 23715
rect 104989 23675 105047 23681
rect 104544 23616 104940 23644
rect 104544 23517 104572 23616
rect 104618 23536 104624 23588
rect 104676 23576 104682 23588
rect 104805 23579 104863 23585
rect 104805 23576 104817 23579
rect 104676 23548 104817 23576
rect 104676 23536 104682 23548
rect 104805 23545 104817 23548
rect 104851 23545 104863 23579
rect 104805 23539 104863 23545
rect 104529 23511 104587 23517
rect 104529 23477 104541 23511
rect 104575 23477 104587 23511
rect 104529 23471 104587 23477
rect 104710 23468 104716 23520
rect 104768 23508 104774 23520
rect 105004 23508 105032 23675
rect 104768 23480 105032 23508
rect 104768 23468 104774 23480
rect 1104 23418 7912 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 7912 23418
rect 1104 23344 7912 23366
rect 104052 23418 110860 23440
rect 104052 23366 107026 23418
rect 107078 23366 107090 23418
rect 107142 23366 107154 23418
rect 107206 23366 107218 23418
rect 107270 23366 107282 23418
rect 107334 23366 110860 23418
rect 104052 23344 110860 23366
rect 1104 22874 7912 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 7912 22874
rect 1104 22800 7912 22822
rect 104052 22874 110860 22896
rect 104052 22822 107762 22874
rect 107814 22822 107826 22874
rect 107878 22822 107890 22874
rect 107942 22822 107954 22874
rect 108006 22822 108018 22874
rect 108070 22822 110860 22874
rect 104052 22800 110860 22822
rect 1104 22330 7912 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 7912 22330
rect 1104 22256 7912 22278
rect 104052 22330 110860 22352
rect 104052 22278 107026 22330
rect 107078 22278 107090 22330
rect 107142 22278 107154 22330
rect 107206 22278 107218 22330
rect 107270 22278 107282 22330
rect 107334 22278 110860 22330
rect 104052 22256 110860 22278
rect 1104 21786 7912 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 7912 21786
rect 1104 21712 7912 21734
rect 104052 21786 110860 21808
rect 104052 21734 107762 21786
rect 107814 21734 107826 21786
rect 107878 21734 107890 21786
rect 107942 21734 107954 21786
rect 108006 21734 108018 21786
rect 108070 21734 110860 21786
rect 104052 21712 110860 21734
rect 1104 21242 7912 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 7912 21242
rect 1104 21168 7912 21190
rect 104052 21242 110860 21264
rect 104052 21190 107026 21242
rect 107078 21190 107090 21242
rect 107142 21190 107154 21242
rect 107206 21190 107218 21242
rect 107270 21190 107282 21242
rect 107334 21190 110860 21242
rect 104052 21168 110860 21190
rect 104345 20995 104403 21001
rect 104345 20961 104357 20995
rect 104391 20992 104403 20995
rect 106366 20992 106372 21004
rect 104391 20964 106372 20992
rect 104391 20961 104403 20964
rect 104345 20955 104403 20961
rect 106366 20952 106372 20964
rect 106424 20952 106430 21004
rect 104342 20816 104348 20868
rect 104400 20856 104406 20868
rect 104621 20859 104679 20865
rect 104621 20856 104633 20859
rect 104400 20828 104633 20856
rect 104400 20816 104406 20828
rect 104621 20825 104633 20828
rect 104667 20825 104679 20859
rect 104621 20819 104679 20825
rect 104894 20816 104900 20868
rect 104952 20856 104958 20868
rect 104952 20828 105110 20856
rect 104952 20816 104958 20828
rect 106090 20748 106096 20800
rect 106148 20788 106154 20800
rect 106185 20791 106243 20797
rect 106185 20788 106197 20791
rect 106148 20760 106197 20788
rect 106148 20748 106154 20760
rect 106185 20757 106197 20760
rect 106231 20757 106243 20791
rect 106185 20751 106243 20757
rect 1104 20698 7912 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 7912 20698
rect 1104 20624 7912 20646
rect 104052 20698 110860 20720
rect 104052 20646 107762 20698
rect 107814 20646 107826 20698
rect 107878 20646 107890 20698
rect 107942 20646 107954 20698
rect 108006 20646 108018 20698
rect 108070 20646 110860 20698
rect 104052 20624 110860 20646
rect 104250 20340 104256 20392
rect 104308 20380 104314 20392
rect 104989 20383 105047 20389
rect 104989 20380 105001 20383
rect 104308 20352 105001 20380
rect 104308 20340 104314 20352
rect 104989 20349 105001 20352
rect 105035 20380 105047 20383
rect 106090 20380 106096 20392
rect 105035 20352 106096 20380
rect 105035 20349 105047 20352
rect 104989 20343 105047 20349
rect 106090 20340 106096 20352
rect 106148 20340 106154 20392
rect 104437 20247 104495 20253
rect 104437 20213 104449 20247
rect 104483 20244 104495 20247
rect 104710 20244 104716 20256
rect 104483 20216 104716 20244
rect 104483 20213 104495 20216
rect 104437 20207 104495 20213
rect 104710 20204 104716 20216
rect 104768 20204 104774 20256
rect 1104 20154 7912 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 7912 20154
rect 1104 20080 7912 20102
rect 104052 20154 110860 20176
rect 104052 20102 107026 20154
rect 107078 20102 107090 20154
rect 107142 20102 107154 20154
rect 107206 20102 107218 20154
rect 107270 20102 107282 20154
rect 107334 20102 110860 20154
rect 104052 20080 110860 20102
rect 104250 19660 104256 19712
rect 104308 19700 104314 19712
rect 104345 19703 104403 19709
rect 104345 19700 104357 19703
rect 104308 19672 104357 19700
rect 104308 19660 104314 19672
rect 104345 19669 104357 19672
rect 104391 19669 104403 19703
rect 104345 19663 104403 19669
rect 1104 19610 7912 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 7912 19610
rect 1104 19536 7912 19558
rect 104052 19610 110860 19632
rect 104052 19558 107762 19610
rect 107814 19558 107826 19610
rect 107878 19558 107890 19610
rect 107942 19558 107954 19610
rect 108006 19558 108018 19610
rect 108070 19558 110860 19610
rect 104052 19536 110860 19558
rect 104710 19320 104716 19372
rect 104768 19320 104774 19372
rect 104342 19252 104348 19304
rect 104400 19252 104406 19304
rect 104618 19252 104624 19304
rect 104676 19252 104682 19304
rect 1104 19066 7912 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 7912 19066
rect 1104 18992 7912 19014
rect 104052 19066 110860 19088
rect 104052 19014 107026 19066
rect 107078 19014 107090 19066
rect 107142 19014 107154 19066
rect 107206 19014 107218 19066
rect 107270 19014 107282 19066
rect 107334 19014 110860 19066
rect 104052 18992 110860 19014
rect 1104 18522 7912 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 7912 18522
rect 1104 18448 7912 18470
rect 104052 18522 110860 18544
rect 104052 18470 107762 18522
rect 107814 18470 107826 18522
rect 107878 18470 107890 18522
rect 107942 18470 107954 18522
rect 108006 18470 108018 18522
rect 108070 18470 110860 18522
rect 104052 18448 110860 18470
rect 1104 17978 7912 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 7912 17978
rect 1104 17904 7912 17926
rect 104052 17978 110860 18000
rect 104052 17926 107026 17978
rect 107078 17926 107090 17978
rect 107142 17926 107154 17978
rect 107206 17926 107218 17978
rect 107270 17926 107282 17978
rect 107334 17926 110860 17978
rect 104052 17904 110860 17926
rect 1104 17434 7912 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 7912 17434
rect 1104 17360 7912 17382
rect 104052 17434 110860 17456
rect 104052 17382 107762 17434
rect 107814 17382 107826 17434
rect 107878 17382 107890 17434
rect 107942 17382 107954 17434
rect 108006 17382 108018 17434
rect 108070 17382 110860 17434
rect 104052 17360 110860 17382
rect 1104 16890 7912 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 7912 16890
rect 1104 16816 7912 16838
rect 104052 16890 110860 16912
rect 104052 16838 107026 16890
rect 107078 16838 107090 16890
rect 107142 16838 107154 16890
rect 107206 16838 107218 16890
rect 107270 16838 107282 16890
rect 107334 16838 110860 16890
rect 104052 16816 110860 16838
rect 1104 16346 7912 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 7912 16346
rect 1104 16272 7912 16294
rect 104052 16346 110860 16368
rect 104052 16294 107762 16346
rect 107814 16294 107826 16346
rect 107878 16294 107890 16346
rect 107942 16294 107954 16346
rect 108006 16294 108018 16346
rect 108070 16294 110860 16346
rect 104052 16272 110860 16294
rect 1104 15802 7912 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 7912 15802
rect 1104 15728 7912 15750
rect 104052 15802 110860 15824
rect 104052 15750 107026 15802
rect 107078 15750 107090 15802
rect 107142 15750 107154 15802
rect 107206 15750 107218 15802
rect 107270 15750 107282 15802
rect 107334 15750 110860 15802
rect 104052 15728 110860 15750
rect 7558 15512 7564 15564
rect 7616 15512 7622 15564
rect 1104 15258 7912 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 7912 15258
rect 1104 15184 7912 15206
rect 104052 15258 110860 15280
rect 104052 15206 107762 15258
rect 107814 15206 107826 15258
rect 107878 15206 107890 15258
rect 107942 15206 107954 15258
rect 108006 15206 108018 15258
rect 108070 15206 110860 15258
rect 104052 15184 110860 15206
rect 1104 14714 7912 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 7912 14714
rect 1104 14640 7912 14662
rect 104052 14714 110860 14736
rect 104052 14662 107026 14714
rect 107078 14662 107090 14714
rect 107142 14662 107154 14714
rect 107206 14662 107218 14714
rect 107270 14662 107282 14714
rect 107334 14662 110860 14714
rect 104052 14640 110860 14662
rect 1104 14170 7912 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 7912 14170
rect 1104 14096 7912 14118
rect 104052 14170 110860 14192
rect 104052 14118 107762 14170
rect 107814 14118 107826 14170
rect 107878 14118 107890 14170
rect 107942 14118 107954 14170
rect 108006 14118 108018 14170
rect 108070 14118 110860 14170
rect 104052 14096 110860 14118
rect 1104 13626 7912 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 7912 13626
rect 1104 13552 7912 13574
rect 104052 13626 110860 13648
rect 104052 13574 107026 13626
rect 107078 13574 107090 13626
rect 107142 13574 107154 13626
rect 107206 13574 107218 13626
rect 107270 13574 107282 13626
rect 107334 13574 110860 13626
rect 104052 13552 110860 13574
rect 1104 13082 7912 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 7912 13082
rect 1104 13008 7912 13030
rect 104052 13082 110860 13104
rect 104052 13030 107762 13082
rect 107814 13030 107826 13082
rect 107878 13030 107890 13082
rect 107942 13030 107954 13082
rect 108006 13030 108018 13082
rect 108070 13030 110860 13082
rect 104052 13008 110860 13030
rect 1104 12538 7912 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 7912 12538
rect 1104 12464 7912 12486
rect 104052 12538 110860 12560
rect 104052 12486 107026 12538
rect 107078 12486 107090 12538
rect 107142 12486 107154 12538
rect 107206 12486 107218 12538
rect 107270 12486 107282 12538
rect 107334 12486 110860 12538
rect 104052 12464 110860 12486
rect 1104 11994 7912 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 7912 11994
rect 1104 11920 7912 11942
rect 104052 11994 110860 12016
rect 104052 11942 107762 11994
rect 107814 11942 107826 11994
rect 107878 11942 107890 11994
rect 107942 11942 107954 11994
rect 108006 11942 108018 11994
rect 108070 11942 110860 11994
rect 104052 11920 110860 11942
rect 102778 11704 102784 11756
rect 102836 11744 102842 11756
rect 110414 11744 110420 11756
rect 102836 11716 110420 11744
rect 102836 11704 102842 11716
rect 110414 11704 110420 11716
rect 110472 11704 110478 11756
rect 1104 11450 7912 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 7912 11450
rect 1104 11376 7912 11398
rect 104052 11450 110860 11472
rect 104052 11398 107026 11450
rect 107078 11398 107090 11450
rect 107142 11398 107154 11450
rect 107206 11398 107218 11450
rect 107270 11398 107282 11450
rect 107334 11398 110860 11450
rect 104052 11376 110860 11398
rect 1104 10906 7912 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 7912 10906
rect 1104 10832 7912 10854
rect 104052 10906 110860 10928
rect 104052 10854 107762 10906
rect 107814 10854 107826 10906
rect 107878 10854 107890 10906
rect 107942 10854 107954 10906
rect 108006 10854 108018 10906
rect 108070 10854 110860 10906
rect 104052 10832 110860 10854
rect 1104 10362 7912 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 7912 10362
rect 1104 10288 7912 10310
rect 104052 10362 110860 10384
rect 104052 10310 107026 10362
rect 107078 10310 107090 10362
rect 107142 10310 107154 10362
rect 107206 10310 107218 10362
rect 107270 10310 107282 10362
rect 107334 10310 110860 10362
rect 104052 10288 110860 10310
rect 90358 10004 90364 10056
rect 90416 10044 90422 10056
rect 104434 10044 104440 10056
rect 90416 10016 104440 10044
rect 90416 10004 90422 10016
rect 104434 10004 104440 10016
rect 104492 10004 104498 10056
rect 90726 9936 90732 9988
rect 90784 9976 90790 9988
rect 104158 9976 104164 9988
rect 90784 9948 104164 9976
rect 90784 9936 90790 9948
rect 104158 9936 104164 9948
rect 104216 9936 104222 9988
rect 1104 9818 7912 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 7912 9818
rect 1104 9744 7912 9766
rect 104052 9818 110860 9840
rect 104052 9766 107762 9818
rect 107814 9766 107826 9818
rect 107878 9766 107890 9818
rect 107942 9766 107954 9818
rect 108006 9766 108018 9818
rect 108070 9766 110860 9818
rect 104052 9744 110860 9766
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 16022 9636 16028 9648
rect 8260 9608 16028 9636
rect 8260 9596 8266 9608
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 1104 9274 7912 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 7912 9274
rect 1104 9200 7912 9222
rect 104052 9274 110860 9296
rect 104052 9222 107026 9274
rect 107078 9222 107090 9274
rect 107142 9222 107154 9274
rect 107206 9222 107218 9274
rect 107270 9222 107282 9274
rect 107334 9222 110860 9274
rect 104052 9200 110860 9222
rect 1104 8730 7912 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 7912 8730
rect 1104 8656 7912 8678
rect 104052 8730 110860 8752
rect 104052 8678 107762 8730
rect 107814 8678 107826 8730
rect 107878 8678 107890 8730
rect 107942 8678 107954 8730
rect 108006 8678 108018 8730
rect 108070 8678 110860 8730
rect 104052 8656 110860 8678
rect 1104 8186 7912 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 7912 8186
rect 1104 8112 7912 8134
rect 104052 8186 110860 8208
rect 104052 8134 107026 8186
rect 107078 8134 107090 8186
rect 107142 8134 107154 8186
rect 107206 8134 107218 8186
rect 107270 8134 107282 8186
rect 107334 8134 110860 8186
rect 104052 8112 110860 8134
rect 1104 7642 110860 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 66314 7642
rect 66366 7590 66378 7642
rect 66430 7590 66442 7642
rect 66494 7590 66506 7642
rect 66558 7590 66570 7642
rect 66622 7590 97034 7642
rect 97086 7590 97098 7642
rect 97150 7590 97162 7642
rect 97214 7590 97226 7642
rect 97278 7590 97290 7642
rect 97342 7590 107762 7642
rect 107814 7590 107826 7642
rect 107878 7590 107890 7642
rect 107942 7590 107954 7642
rect 108006 7590 108018 7642
rect 108070 7590 110860 7642
rect 1104 7568 110860 7590
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 16080 7500 16129 7528
rect 16080 7488 16086 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16117 7491 16175 7497
rect 23198 7488 23204 7540
rect 23256 7528 23262 7540
rect 23474 7528 23480 7540
rect 23256 7500 23480 7528
rect 23256 7488 23262 7500
rect 23474 7488 23480 7500
rect 23532 7488 23538 7540
rect 24670 7488 24676 7540
rect 24728 7488 24734 7540
rect 25774 7488 25780 7540
rect 25832 7528 25838 7540
rect 25869 7531 25927 7537
rect 25869 7528 25881 7531
rect 25832 7500 25881 7528
rect 25832 7488 25838 7500
rect 25869 7497 25881 7500
rect 25915 7497 25927 7531
rect 25869 7491 25927 7497
rect 26970 7488 26976 7540
rect 27028 7488 27034 7540
rect 28258 7488 28264 7540
rect 28316 7488 28322 7540
rect 28994 7488 29000 7540
rect 29052 7528 29058 7540
rect 29549 7531 29607 7537
rect 29549 7528 29561 7531
rect 29052 7500 29561 7528
rect 29052 7488 29058 7500
rect 29549 7497 29561 7500
rect 29595 7497 29607 7531
rect 29549 7491 29607 7497
rect 30466 7488 30472 7540
rect 30524 7488 30530 7540
rect 31570 7488 31576 7540
rect 31628 7528 31634 7540
rect 31757 7531 31815 7537
rect 31757 7528 31769 7531
rect 31628 7500 31769 7528
rect 31628 7488 31634 7500
rect 31757 7497 31769 7500
rect 31803 7497 31815 7531
rect 31757 7491 31815 7497
rect 32858 7488 32864 7540
rect 32916 7488 32922 7540
rect 33962 7488 33968 7540
rect 34020 7488 34026 7540
rect 35250 7488 35256 7540
rect 35308 7488 35314 7540
rect 36078 7488 36084 7540
rect 36136 7528 36142 7540
rect 36354 7528 36360 7540
rect 36136 7500 36360 7528
rect 36136 7488 36142 7500
rect 36354 7488 36360 7500
rect 36412 7488 36418 7540
rect 37458 7488 37464 7540
rect 37516 7488 37522 7540
rect 38654 7488 38660 7540
rect 38712 7488 38718 7540
rect 39850 7488 39856 7540
rect 39908 7488 39914 7540
rect 41046 7488 41052 7540
rect 41104 7488 41110 7540
rect 41874 7488 41880 7540
rect 41932 7528 41938 7540
rect 42150 7528 42156 7540
rect 41932 7500 42156 7528
rect 41932 7488 41938 7500
rect 42150 7488 42156 7500
rect 42208 7488 42214 7540
rect 43346 7488 43352 7540
rect 43404 7488 43410 7540
rect 90542 7488 90548 7540
rect 90600 7488 90606 7540
rect 90726 7488 90732 7540
rect 90784 7488 90790 7540
rect 91002 7488 91008 7540
rect 91060 7488 91066 7540
rect 1104 7098 110860 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 107026 7098
rect 107078 7046 107090 7098
rect 107142 7046 107154 7098
rect 107206 7046 107218 7098
rect 107270 7046 107282 7098
rect 107334 7046 110860 7098
rect 1104 7024 110860 7046
rect 1104 6554 110860 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 66314 6554
rect 66366 6502 66378 6554
rect 66430 6502 66442 6554
rect 66494 6502 66506 6554
rect 66558 6502 66570 6554
rect 66622 6502 97034 6554
rect 97086 6502 97098 6554
rect 97150 6502 97162 6554
rect 97214 6502 97226 6554
rect 97278 6502 97290 6554
rect 97342 6502 110860 6554
rect 1104 6480 110860 6502
rect 1104 6010 110860 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 110860 6010
rect 1104 5936 110860 5958
rect 1104 5466 110860 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 66314 5466
rect 66366 5414 66378 5466
rect 66430 5414 66442 5466
rect 66494 5414 66506 5466
rect 66558 5414 66570 5466
rect 66622 5414 97034 5466
rect 97086 5414 97098 5466
rect 97150 5414 97162 5466
rect 97214 5414 97226 5466
rect 97278 5414 97290 5466
rect 97342 5414 110860 5466
rect 1104 5392 110860 5414
rect 1104 4922 110860 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 110860 4922
rect 1104 4848 110860 4870
rect 1104 4378 110860 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 66314 4378
rect 66366 4326 66378 4378
rect 66430 4326 66442 4378
rect 66494 4326 66506 4378
rect 66558 4326 66570 4378
rect 66622 4326 97034 4378
rect 97086 4326 97098 4378
rect 97150 4326 97162 4378
rect 97214 4326 97226 4378
rect 97278 4326 97290 4378
rect 97342 4326 110860 4378
rect 1104 4304 110860 4326
rect 1104 3834 110860 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 110860 3834
rect 1104 3760 110860 3782
rect 1104 3290 110860 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 66314 3290
rect 66366 3238 66378 3290
rect 66430 3238 66442 3290
rect 66494 3238 66506 3290
rect 66558 3238 66570 3290
rect 66622 3238 97034 3290
rect 97086 3238 97098 3290
rect 97150 3238 97162 3290
rect 97214 3238 97226 3290
rect 97278 3238 97290 3290
rect 97342 3238 110860 3290
rect 1104 3216 110860 3238
rect 1104 2746 110860 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 110860 2746
rect 1104 2672 110860 2694
rect 1104 2202 110860 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 66314 2202
rect 66366 2150 66378 2202
rect 66430 2150 66442 2202
rect 66494 2150 66506 2202
rect 66558 2150 66570 2202
rect 66622 2150 97034 2202
rect 97086 2150 97098 2202
rect 97150 2150 97162 2202
rect 97214 2150 97226 2202
rect 97278 2150 97290 2202
rect 97342 2150 110860 2202
rect 1104 2128 110860 2150
<< via1 >>
rect 4874 71782 4926 71834
rect 4938 71782 4990 71834
rect 5002 71782 5054 71834
rect 5066 71782 5118 71834
rect 5130 71782 5182 71834
rect 35594 71782 35646 71834
rect 35658 71782 35710 71834
rect 35722 71782 35774 71834
rect 35786 71782 35838 71834
rect 35850 71782 35902 71834
rect 66314 71782 66366 71834
rect 66378 71782 66430 71834
rect 66442 71782 66494 71834
rect 66506 71782 66558 71834
rect 66570 71782 66622 71834
rect 97034 71782 97086 71834
rect 97098 71782 97150 71834
rect 97162 71782 97214 71834
rect 97226 71782 97278 71834
rect 97290 71782 97342 71834
rect 44456 71680 44508 71732
rect 47032 71680 47084 71732
rect 49608 71680 49660 71732
rect 51540 71680 51592 71732
rect 53472 71680 53524 71732
rect 55404 71680 55456 71732
rect 57336 71680 57388 71732
rect 59268 71680 59320 71732
rect 61200 71680 61252 71732
rect 63132 71680 63184 71732
rect 65708 71680 65760 71732
rect 67640 71680 67692 71732
rect 69572 71680 69624 71732
rect 71504 71680 71556 71732
rect 74080 71680 74132 71732
rect 77300 71680 77352 71732
rect 45100 71544 45152 71596
rect 47308 71544 47360 71596
rect 49516 71544 49568 71596
rect 51632 71587 51684 71596
rect 51632 71553 51641 71587
rect 51641 71553 51675 71587
rect 51675 71553 51684 71587
rect 51632 71544 51684 71553
rect 53564 71587 53616 71596
rect 53564 71553 53573 71587
rect 53573 71553 53607 71587
rect 53607 71553 53616 71587
rect 53564 71544 53616 71553
rect 55496 71587 55548 71596
rect 55496 71553 55505 71587
rect 55505 71553 55539 71587
rect 55539 71553 55548 71587
rect 55496 71544 55548 71553
rect 57428 71587 57480 71596
rect 57428 71553 57437 71587
rect 57437 71553 57471 71587
rect 57471 71553 57480 71587
rect 57428 71544 57480 71553
rect 59636 71587 59688 71596
rect 59636 71553 59645 71587
rect 59645 71553 59679 71587
rect 59679 71553 59688 71587
rect 59636 71544 59688 71553
rect 61568 71587 61620 71596
rect 61568 71553 61577 71587
rect 61577 71553 61611 71587
rect 61611 71553 61620 71587
rect 61568 71544 61620 71553
rect 63132 71544 63184 71596
rect 65432 71544 65484 71596
rect 67364 71544 67416 71596
rect 69940 71587 69992 71596
rect 69940 71553 69949 71587
rect 69949 71553 69983 71587
rect 69983 71553 69992 71587
rect 69940 71544 69992 71553
rect 71872 71587 71924 71596
rect 71872 71553 71881 71587
rect 71881 71553 71915 71587
rect 71915 71553 71924 71587
rect 71872 71544 71924 71553
rect 74172 71587 74224 71596
rect 74172 71553 74181 71587
rect 74181 71553 74215 71587
rect 74215 71553 74224 71587
rect 74172 71544 74224 71553
rect 76104 71544 76156 71596
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 34934 71238 34986 71290
rect 34998 71238 35050 71290
rect 35062 71238 35114 71290
rect 35126 71238 35178 71290
rect 35190 71238 35242 71290
rect 65654 71238 65706 71290
rect 65718 71238 65770 71290
rect 65782 71238 65834 71290
rect 65846 71238 65898 71290
rect 65910 71238 65962 71290
rect 96374 71238 96426 71290
rect 96438 71238 96490 71290
rect 96502 71238 96554 71290
rect 96566 71238 96618 71290
rect 96630 71238 96682 71290
rect 4874 70694 4926 70746
rect 4938 70694 4990 70746
rect 5002 70694 5054 70746
rect 5066 70694 5118 70746
rect 5130 70694 5182 70746
rect 35594 70694 35646 70746
rect 35658 70694 35710 70746
rect 35722 70694 35774 70746
rect 35786 70694 35838 70746
rect 35850 70694 35902 70746
rect 66314 70694 66366 70746
rect 66378 70694 66430 70746
rect 66442 70694 66494 70746
rect 66506 70694 66558 70746
rect 66570 70694 66622 70746
rect 97034 70694 97086 70746
rect 97098 70694 97150 70746
rect 97162 70694 97214 70746
rect 97226 70694 97278 70746
rect 97290 70694 97342 70746
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 34934 70150 34986 70202
rect 34998 70150 35050 70202
rect 35062 70150 35114 70202
rect 35126 70150 35178 70202
rect 35190 70150 35242 70202
rect 65654 70150 65706 70202
rect 65718 70150 65770 70202
rect 65782 70150 65834 70202
rect 65846 70150 65898 70202
rect 65910 70150 65962 70202
rect 96374 70150 96426 70202
rect 96438 70150 96490 70202
rect 96502 70150 96554 70202
rect 96566 70150 96618 70202
rect 96630 70150 96682 70202
rect 4874 69606 4926 69658
rect 4938 69606 4990 69658
rect 5002 69606 5054 69658
rect 5066 69606 5118 69658
rect 5130 69606 5182 69658
rect 35594 69606 35646 69658
rect 35658 69606 35710 69658
rect 35722 69606 35774 69658
rect 35786 69606 35838 69658
rect 35850 69606 35902 69658
rect 66314 69606 66366 69658
rect 66378 69606 66430 69658
rect 66442 69606 66494 69658
rect 66506 69606 66558 69658
rect 66570 69606 66622 69658
rect 97034 69606 97086 69658
rect 97098 69606 97150 69658
rect 97162 69606 97214 69658
rect 97226 69606 97278 69658
rect 97290 69606 97342 69658
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 96374 69062 96426 69114
rect 96438 69062 96490 69114
rect 96502 69062 96554 69114
rect 96566 69062 96618 69114
rect 96630 69062 96682 69114
rect 4874 68518 4926 68570
rect 4938 68518 4990 68570
rect 5002 68518 5054 68570
rect 5066 68518 5118 68570
rect 5130 68518 5182 68570
rect 35594 68518 35646 68570
rect 35658 68518 35710 68570
rect 35722 68518 35774 68570
rect 35786 68518 35838 68570
rect 35850 68518 35902 68570
rect 66314 68518 66366 68570
rect 66378 68518 66430 68570
rect 66442 68518 66494 68570
rect 66506 68518 66558 68570
rect 66570 68518 66622 68570
rect 97034 68518 97086 68570
rect 97098 68518 97150 68570
rect 97162 68518 97214 68570
rect 97226 68518 97278 68570
rect 97290 68518 97342 68570
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 96374 67974 96426 68026
rect 96438 67974 96490 68026
rect 96502 67974 96554 68026
rect 96566 67974 96618 68026
rect 96630 67974 96682 68026
rect 4874 67430 4926 67482
rect 4938 67430 4990 67482
rect 5002 67430 5054 67482
rect 5066 67430 5118 67482
rect 5130 67430 5182 67482
rect 35594 67430 35646 67482
rect 35658 67430 35710 67482
rect 35722 67430 35774 67482
rect 35786 67430 35838 67482
rect 35850 67430 35902 67482
rect 66314 67430 66366 67482
rect 66378 67430 66430 67482
rect 66442 67430 66494 67482
rect 66506 67430 66558 67482
rect 66570 67430 66622 67482
rect 97034 67430 97086 67482
rect 97098 67430 97150 67482
rect 97162 67430 97214 67482
rect 97226 67430 97278 67482
rect 97290 67430 97342 67482
rect 8208 67124 8260 67176
rect 44732 67192 44784 67244
rect 46940 67192 46992 67244
rect 49516 67371 49568 67380
rect 49516 67337 49525 67371
rect 49525 67337 49559 67371
rect 49559 67337 49568 67371
rect 49516 67328 49568 67337
rect 51632 67328 51684 67380
rect 55496 67328 55548 67380
rect 57428 67328 57480 67380
rect 59636 67371 59688 67380
rect 59636 67337 59645 67371
rect 59645 67337 59679 67371
rect 59679 67337 59688 67371
rect 59636 67328 59688 67337
rect 53932 67260 53984 67312
rect 57796 67260 57848 67312
rect 60832 67328 60884 67380
rect 61568 67328 61620 67380
rect 65432 67371 65484 67380
rect 65432 67337 65441 67371
rect 65441 67337 65475 67371
rect 65475 67337 65484 67371
rect 65432 67328 65484 67337
rect 67364 67371 67416 67380
rect 67364 67337 67373 67371
rect 67373 67337 67407 67371
rect 67407 67337 67416 67371
rect 67364 67328 67416 67337
rect 68744 67328 68796 67380
rect 62028 67260 62080 67312
rect 66168 67260 66220 67312
rect 67548 67260 67600 67312
rect 69940 67371 69992 67380
rect 69940 67337 69949 67371
rect 69949 67337 69983 67371
rect 69983 67337 69992 67371
rect 69940 67328 69992 67337
rect 71872 67328 71924 67380
rect 76104 67371 76156 67380
rect 76104 67337 76113 67371
rect 76113 67337 76147 67371
rect 76147 67337 76156 67371
rect 76104 67328 76156 67337
rect 74080 67260 74132 67312
rect 47676 67192 47728 67244
rect 49148 67192 49200 67244
rect 54944 67192 54996 67244
rect 65524 67192 65576 67244
rect 69572 67192 69624 67244
rect 71412 67192 71464 67244
rect 75736 67192 75788 67244
rect 43168 67031 43220 67040
rect 43168 66997 43177 67031
rect 43177 66997 43211 67031
rect 43211 66997 43220 67031
rect 45100 67167 45152 67176
rect 45100 67133 45109 67167
rect 45109 67133 45143 67167
rect 45143 67133 45152 67167
rect 45100 67124 45152 67133
rect 43168 66988 43220 66997
rect 45376 67031 45428 67040
rect 45376 66997 45385 67031
rect 45385 66997 45419 67031
rect 45419 66997 45428 67031
rect 47308 67167 47360 67176
rect 47308 67133 47317 67167
rect 47317 67133 47351 67167
rect 47351 67133 47360 67167
rect 47308 67124 47360 67133
rect 49700 67167 49752 67176
rect 49700 67133 49709 67167
rect 49709 67133 49743 67167
rect 49743 67133 49752 67167
rect 49700 67124 49752 67133
rect 49976 67167 50028 67176
rect 49976 67133 49985 67167
rect 49985 67133 50019 67167
rect 50019 67133 50028 67167
rect 49976 67124 50028 67133
rect 53472 67124 53524 67176
rect 55404 67167 55456 67176
rect 55404 67133 55413 67167
rect 55413 67133 55447 67167
rect 55447 67133 55456 67167
rect 55404 67124 55456 67133
rect 55680 67167 55732 67176
rect 55680 67133 55689 67167
rect 55689 67133 55723 67167
rect 55723 67133 55732 67167
rect 55680 67124 55732 67133
rect 57888 67167 57940 67176
rect 57888 67133 57897 67167
rect 57897 67133 57931 67167
rect 57931 67133 57940 67167
rect 57888 67124 57940 67133
rect 58164 67167 58216 67176
rect 58164 67133 58173 67167
rect 58173 67133 58207 67167
rect 58207 67133 58216 67167
rect 58164 67124 58216 67133
rect 59728 67167 59780 67176
rect 59728 67133 59737 67167
rect 59737 67133 59771 67167
rect 59771 67133 59780 67167
rect 59728 67124 59780 67133
rect 60004 67167 60056 67176
rect 60004 67133 60013 67167
rect 60013 67133 60047 67167
rect 60047 67133 60056 67167
rect 60004 67124 60056 67133
rect 45376 66988 45428 66997
rect 47584 67031 47636 67040
rect 47584 66997 47593 67031
rect 47593 66997 47627 67031
rect 47627 66997 47636 67031
rect 47584 66988 47636 66997
rect 49700 66988 49752 67040
rect 51632 66988 51684 67040
rect 53656 66988 53708 67040
rect 61292 66988 61344 67040
rect 63960 67167 64012 67176
rect 63960 67133 63969 67167
rect 63969 67133 64003 67167
rect 64003 67133 64012 67167
rect 63960 67124 64012 67133
rect 64696 67124 64748 67176
rect 65524 66988 65576 67040
rect 68008 67031 68060 67040
rect 68008 66997 68017 67031
rect 68017 66997 68051 67031
rect 68051 66997 68060 67031
rect 68468 67167 68520 67176
rect 68468 67133 68477 67167
rect 68477 67133 68511 67167
rect 68511 67133 68520 67167
rect 68468 67124 68520 67133
rect 69940 67124 69992 67176
rect 68008 66988 68060 66997
rect 69940 66988 69992 67040
rect 73712 66988 73764 67040
rect 95884 66988 95936 67040
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 96374 66886 96426 66938
rect 96438 66886 96490 66938
rect 96502 66886 96554 66938
rect 96566 66886 96618 66938
rect 96630 66886 96682 66938
rect 47676 66827 47728 66836
rect 47676 66793 47685 66827
rect 47685 66793 47719 66827
rect 47719 66793 47728 66827
rect 49700 66827 49752 66836
rect 47676 66784 47728 66793
rect 49700 66793 49709 66827
rect 49709 66793 49743 66827
rect 49743 66793 49752 66827
rect 49700 66784 49752 66793
rect 53564 66784 53616 66836
rect 54944 66784 54996 66836
rect 57980 66784 58032 66836
rect 59728 66784 59780 66836
rect 61292 66827 61344 66836
rect 61292 66793 61301 66827
rect 61301 66793 61335 66827
rect 61335 66793 61344 66827
rect 61292 66784 61344 66793
rect 65524 66784 65576 66836
rect 68008 66784 68060 66836
rect 69940 66827 69992 66836
rect 69940 66793 69949 66827
rect 69949 66793 69983 66827
rect 69983 66793 69992 66827
rect 69940 66784 69992 66793
rect 73712 66827 73764 66836
rect 73712 66793 73721 66827
rect 73721 66793 73755 66827
rect 73755 66793 73764 66827
rect 73712 66784 73764 66793
rect 44732 66716 44784 66768
rect 48688 66716 48740 66768
rect 46940 66648 46992 66700
rect 50528 66648 50580 66700
rect 51632 66691 51684 66700
rect 51632 66657 51641 66691
rect 51641 66657 51675 66691
rect 51675 66657 51684 66691
rect 53472 66691 53524 66700
rect 51632 66648 51684 66657
rect 53472 66657 53481 66691
rect 53481 66657 53515 66691
rect 53515 66657 53524 66691
rect 53472 66648 53524 66657
rect 63132 66759 63184 66768
rect 63132 66725 63141 66759
rect 63141 66725 63175 66759
rect 63175 66725 63184 66759
rect 63132 66716 63184 66725
rect 55404 66580 55456 66632
rect 49700 66512 49752 66564
rect 55312 66512 55364 66564
rect 61660 66555 61712 66564
rect 61660 66521 61669 66555
rect 61669 66521 61703 66555
rect 61703 66521 61712 66555
rect 61660 66512 61712 66521
rect 64880 66512 64932 66564
rect 71228 66512 71280 66564
rect 73436 66512 73488 66564
rect 56600 66444 56652 66496
rect 74172 66444 74224 66496
rect 4874 66342 4926 66394
rect 4938 66342 4990 66394
rect 5002 66342 5054 66394
rect 5066 66342 5118 66394
rect 5130 66342 5182 66394
rect 35594 66342 35646 66394
rect 35658 66342 35710 66394
rect 35722 66342 35774 66394
rect 35786 66342 35838 66394
rect 35850 66342 35902 66394
rect 66314 66342 66366 66394
rect 66378 66342 66430 66394
rect 66442 66342 66494 66394
rect 66506 66342 66558 66394
rect 66570 66342 66622 66394
rect 97034 66342 97086 66394
rect 97098 66342 97150 66394
rect 97162 66342 97214 66394
rect 97226 66342 97278 66394
rect 97290 66342 97342 66394
rect 107762 66342 107814 66394
rect 107826 66342 107878 66394
rect 107890 66342 107942 66394
rect 107954 66342 108006 66394
rect 108018 66342 108070 66394
rect 49148 66240 49200 66292
rect 48688 66215 48740 66224
rect 48688 66181 48697 66215
rect 48697 66181 48731 66215
rect 48731 66181 48740 66215
rect 48688 66172 48740 66181
rect 50528 66215 50580 66224
rect 50528 66181 50537 66215
rect 50537 66181 50571 66215
rect 50571 66181 50580 66215
rect 50528 66172 50580 66181
rect 56600 66240 56652 66292
rect 57888 66240 57940 66292
rect 53932 66172 53984 66224
rect 55312 66172 55364 66224
rect 59728 66240 59780 66292
rect 57980 66147 58032 66156
rect 57980 66113 57989 66147
rect 57989 66113 58023 66147
rect 58023 66113 58032 66147
rect 57980 66104 58032 66113
rect 60832 66215 60884 66224
rect 60832 66181 60841 66215
rect 60841 66181 60875 66215
rect 60875 66181 60884 66215
rect 60832 66172 60884 66181
rect 64604 66104 64656 66156
rect 64880 66215 64932 66224
rect 64880 66181 64889 66215
rect 64889 66181 64923 66215
rect 64923 66181 64932 66215
rect 64880 66172 64932 66181
rect 66168 66172 66220 66224
rect 67548 66172 67600 66224
rect 69572 66215 69624 66224
rect 69572 66181 69581 66215
rect 69581 66181 69615 66215
rect 69615 66181 69624 66215
rect 69572 66172 69624 66181
rect 71412 66215 71464 66224
rect 71412 66181 71421 66215
rect 71421 66181 71455 66215
rect 71455 66181 71464 66215
rect 71412 66172 71464 66181
rect 73436 66215 73488 66224
rect 73436 66181 73445 66215
rect 73445 66181 73479 66215
rect 73479 66181 73488 66215
rect 73436 66172 73488 66181
rect 75736 66240 75788 66292
rect 95884 66215 95936 66224
rect 95884 66181 95893 66215
rect 95893 66181 95927 66215
rect 95927 66181 95936 66215
rect 95884 66172 95936 66181
rect 75736 66147 75788 66156
rect 75736 66113 75745 66147
rect 75745 66113 75779 66147
rect 75779 66113 75788 66147
rect 75736 66104 75788 66113
rect 57796 65900 57848 65952
rect 62028 65900 62080 65952
rect 63408 65943 63460 65952
rect 63408 65909 63417 65943
rect 63417 65909 63451 65943
rect 63451 65909 63460 65943
rect 63408 65900 63460 65909
rect 64604 65900 64656 65952
rect 75736 65900 75788 65952
rect 76288 65900 76340 65952
rect 76472 66036 76524 66088
rect 92388 66147 92440 66156
rect 92388 66113 92397 66147
rect 92397 66113 92431 66147
rect 92431 66113 92440 66147
rect 92388 66104 92440 66113
rect 102784 65968 102836 66020
rect 86316 65943 86368 65952
rect 86316 65909 86325 65943
rect 86325 65909 86359 65943
rect 86359 65909 86368 65943
rect 86316 65900 86368 65909
rect 87328 65943 87380 65952
rect 87328 65909 87337 65943
rect 87337 65909 87371 65943
rect 87371 65909 87380 65943
rect 87328 65900 87380 65909
rect 92296 65943 92348 65952
rect 92296 65909 92305 65943
rect 92305 65909 92339 65943
rect 92339 65909 92348 65943
rect 92296 65900 92348 65909
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 96374 65798 96426 65850
rect 96438 65798 96490 65850
rect 96502 65798 96554 65850
rect 96566 65798 96618 65850
rect 96630 65798 96682 65850
rect 107026 65798 107078 65850
rect 107090 65798 107142 65850
rect 107154 65798 107206 65850
rect 107218 65798 107270 65850
rect 107282 65798 107334 65850
rect 63408 65696 63460 65748
rect 100760 65696 100812 65748
rect 92296 65628 92348 65680
rect 102968 65628 103020 65680
rect 4874 65254 4926 65306
rect 4938 65254 4990 65306
rect 5002 65254 5054 65306
rect 5066 65254 5118 65306
rect 5130 65254 5182 65306
rect 107762 65254 107814 65306
rect 107826 65254 107878 65306
rect 107890 65254 107942 65306
rect 107954 65254 108006 65306
rect 108018 65254 108070 65306
rect 92388 64880 92440 64932
rect 102876 64880 102928 64932
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 107026 64710 107078 64762
rect 107090 64710 107142 64762
rect 107154 64710 107206 64762
rect 107218 64710 107270 64762
rect 107282 64710 107334 64762
rect 100760 64268 100812 64320
rect 104440 64268 104492 64320
rect 4874 64166 4926 64218
rect 4938 64166 4990 64218
rect 5002 64166 5054 64218
rect 5066 64166 5118 64218
rect 5130 64166 5182 64218
rect 107762 64166 107814 64218
rect 107826 64166 107878 64218
rect 107890 64166 107942 64218
rect 107954 64166 108006 64218
rect 108018 64166 108070 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 107026 63622 107078 63674
rect 107090 63622 107142 63674
rect 107154 63622 107206 63674
rect 107218 63622 107270 63674
rect 107282 63622 107334 63674
rect 4874 63078 4926 63130
rect 4938 63078 4990 63130
rect 5002 63078 5054 63130
rect 5066 63078 5118 63130
rect 5130 63078 5182 63130
rect 107762 63078 107814 63130
rect 107826 63078 107878 63130
rect 107890 63078 107942 63130
rect 107954 63078 108006 63130
rect 108018 63078 108070 63130
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 107026 62534 107078 62586
rect 107090 62534 107142 62586
rect 107154 62534 107206 62586
rect 107218 62534 107270 62586
rect 107282 62534 107334 62586
rect 4874 61990 4926 62042
rect 4938 61990 4990 62042
rect 5002 61990 5054 62042
rect 5066 61990 5118 62042
rect 5130 61990 5182 62042
rect 107762 61990 107814 62042
rect 107826 61990 107878 62042
rect 107890 61990 107942 62042
rect 107954 61990 108006 62042
rect 108018 61990 108070 62042
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 107026 61446 107078 61498
rect 107090 61446 107142 61498
rect 107154 61446 107206 61498
rect 107218 61446 107270 61498
rect 107282 61446 107334 61498
rect 4874 60902 4926 60954
rect 4938 60902 4990 60954
rect 5002 60902 5054 60954
rect 5066 60902 5118 60954
rect 5130 60902 5182 60954
rect 107762 60902 107814 60954
rect 107826 60902 107878 60954
rect 107890 60902 107942 60954
rect 107954 60902 108006 60954
rect 108018 60902 108070 60954
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 107026 60358 107078 60410
rect 107090 60358 107142 60410
rect 107154 60358 107206 60410
rect 107218 60358 107270 60410
rect 107282 60358 107334 60410
rect 103704 60052 103756 60104
rect 4874 59814 4926 59866
rect 4938 59814 4990 59866
rect 5002 59814 5054 59866
rect 5066 59814 5118 59866
rect 5130 59814 5182 59866
rect 107762 59814 107814 59866
rect 107826 59814 107878 59866
rect 107890 59814 107942 59866
rect 107954 59814 108006 59866
rect 108018 59814 108070 59866
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 107026 59270 107078 59322
rect 107090 59270 107142 59322
rect 107154 59270 107206 59322
rect 107218 59270 107270 59322
rect 107282 59270 107334 59322
rect 4874 58726 4926 58778
rect 4938 58726 4990 58778
rect 5002 58726 5054 58778
rect 5066 58726 5118 58778
rect 5130 58726 5182 58778
rect 107762 58726 107814 58778
rect 107826 58726 107878 58778
rect 107890 58726 107942 58778
rect 107954 58726 108006 58778
rect 108018 58726 108070 58778
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 107026 58182 107078 58234
rect 107090 58182 107142 58234
rect 107154 58182 107206 58234
rect 107218 58182 107270 58234
rect 107282 58182 107334 58234
rect 102968 57876 103020 57928
rect 4874 57638 4926 57690
rect 4938 57638 4990 57690
rect 5002 57638 5054 57690
rect 5066 57638 5118 57690
rect 5130 57638 5182 57690
rect 107762 57638 107814 57690
rect 107826 57638 107878 57690
rect 107890 57638 107942 57690
rect 107954 57638 108006 57690
rect 108018 57638 108070 57690
rect 104348 57443 104400 57452
rect 104348 57409 104357 57443
rect 104357 57409 104391 57443
rect 104391 57409 104400 57443
rect 104348 57400 104400 57409
rect 104624 57375 104676 57384
rect 104624 57341 104633 57375
rect 104633 57341 104667 57375
rect 104667 57341 104676 57375
rect 104624 57332 104676 57341
rect 104992 57332 105044 57384
rect 106648 57239 106700 57248
rect 106648 57205 106657 57239
rect 106657 57205 106691 57239
rect 106691 57205 106700 57239
rect 106648 57196 106700 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 107026 57094 107078 57146
rect 107090 57094 107142 57146
rect 107154 57094 107206 57146
rect 107218 57094 107270 57146
rect 107282 57094 107334 57146
rect 104992 56899 105044 56908
rect 104992 56865 105001 56899
rect 105001 56865 105035 56899
rect 105035 56865 105044 56899
rect 104992 56856 105044 56865
rect 104532 56652 104584 56704
rect 4874 56550 4926 56602
rect 4938 56550 4990 56602
rect 5002 56550 5054 56602
rect 5066 56550 5118 56602
rect 5130 56550 5182 56602
rect 107762 56550 107814 56602
rect 107826 56550 107878 56602
rect 107890 56550 107942 56602
rect 107954 56550 108006 56602
rect 108018 56550 108070 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 107026 56006 107078 56058
rect 107090 56006 107142 56058
rect 107154 56006 107206 56058
rect 107218 56006 107270 56058
rect 107282 56006 107334 56058
rect 104624 55904 104676 55956
rect 104532 55743 104584 55752
rect 104532 55709 104541 55743
rect 104541 55709 104575 55743
rect 104575 55709 104584 55743
rect 104532 55700 104584 55709
rect 4874 55462 4926 55514
rect 4938 55462 4990 55514
rect 5002 55462 5054 55514
rect 5066 55462 5118 55514
rect 5130 55462 5182 55514
rect 107762 55462 107814 55514
rect 107826 55462 107878 55514
rect 107890 55462 107942 55514
rect 107954 55462 108006 55514
rect 108018 55462 108070 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 107026 54918 107078 54970
rect 107090 54918 107142 54970
rect 107154 54918 107206 54970
rect 107218 54918 107270 54970
rect 107282 54918 107334 54970
rect 104256 54680 104308 54732
rect 106372 54680 106424 54732
rect 104624 54587 104676 54596
rect 104624 54553 104633 54587
rect 104633 54553 104667 54587
rect 104667 54553 104676 54587
rect 104624 54544 104676 54553
rect 105084 54544 105136 54596
rect 106188 54544 106240 54596
rect 4874 54374 4926 54426
rect 4938 54374 4990 54426
rect 5002 54374 5054 54426
rect 5066 54374 5118 54426
rect 5130 54374 5182 54426
rect 107762 54374 107814 54426
rect 107826 54374 107878 54426
rect 107890 54374 107942 54426
rect 107954 54374 108006 54426
rect 108018 54374 108070 54426
rect 105084 54272 105136 54324
rect 102876 54136 102928 54188
rect 104532 54136 104584 54188
rect 104532 53932 104584 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 107026 53830 107078 53882
rect 107090 53830 107142 53882
rect 107154 53830 107206 53882
rect 107218 53830 107270 53882
rect 107282 53830 107334 53882
rect 104624 53728 104676 53780
rect 104992 53771 105044 53780
rect 104992 53737 105001 53771
rect 105001 53737 105035 53771
rect 105035 53737 105044 53771
rect 104992 53728 105044 53737
rect 104900 53592 104952 53644
rect 106188 53592 106240 53644
rect 104808 53524 104860 53576
rect 104992 53524 105044 53576
rect 4874 53286 4926 53338
rect 4938 53286 4990 53338
rect 5002 53286 5054 53338
rect 5066 53286 5118 53338
rect 5130 53286 5182 53338
rect 107762 53286 107814 53338
rect 107826 53286 107878 53338
rect 107890 53286 107942 53338
rect 107954 53286 108006 53338
rect 108018 53286 108070 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 107026 52742 107078 52794
rect 107090 52742 107142 52794
rect 107154 52742 107206 52794
rect 107218 52742 107270 52794
rect 107282 52742 107334 52794
rect 4874 52198 4926 52250
rect 4938 52198 4990 52250
rect 5002 52198 5054 52250
rect 5066 52198 5118 52250
rect 5130 52198 5182 52250
rect 107762 52198 107814 52250
rect 107826 52198 107878 52250
rect 107890 52198 107942 52250
rect 107954 52198 108006 52250
rect 108018 52198 108070 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 107026 51654 107078 51706
rect 107090 51654 107142 51706
rect 107154 51654 107206 51706
rect 107218 51654 107270 51706
rect 107282 51654 107334 51706
rect 4874 51110 4926 51162
rect 4938 51110 4990 51162
rect 5002 51110 5054 51162
rect 5066 51110 5118 51162
rect 5130 51110 5182 51162
rect 107762 51110 107814 51162
rect 107826 51110 107878 51162
rect 107890 51110 107942 51162
rect 107954 51110 108006 51162
rect 108018 51110 108070 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 107026 50566 107078 50618
rect 107090 50566 107142 50618
rect 107154 50566 107206 50618
rect 107218 50566 107270 50618
rect 107282 50566 107334 50618
rect 4874 50022 4926 50074
rect 4938 50022 4990 50074
rect 5002 50022 5054 50074
rect 5066 50022 5118 50074
rect 5130 50022 5182 50074
rect 107762 50022 107814 50074
rect 107826 50022 107878 50074
rect 107890 50022 107942 50074
rect 107954 50022 108006 50074
rect 108018 50022 108070 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 107026 49478 107078 49530
rect 107090 49478 107142 49530
rect 107154 49478 107206 49530
rect 107218 49478 107270 49530
rect 107282 49478 107334 49530
rect 4874 48934 4926 48986
rect 4938 48934 4990 48986
rect 5002 48934 5054 48986
rect 5066 48934 5118 48986
rect 5130 48934 5182 48986
rect 107762 48934 107814 48986
rect 107826 48934 107878 48986
rect 107890 48934 107942 48986
rect 107954 48934 108006 48986
rect 108018 48934 108070 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 107026 48390 107078 48442
rect 107090 48390 107142 48442
rect 107154 48390 107206 48442
rect 107218 48390 107270 48442
rect 107282 48390 107334 48442
rect 4874 47846 4926 47898
rect 4938 47846 4990 47898
rect 5002 47846 5054 47898
rect 5066 47846 5118 47898
rect 5130 47846 5182 47898
rect 107762 47846 107814 47898
rect 107826 47846 107878 47898
rect 107890 47846 107942 47898
rect 107954 47846 108006 47898
rect 108018 47846 108070 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 107026 47302 107078 47354
rect 107090 47302 107142 47354
rect 107154 47302 107206 47354
rect 107218 47302 107270 47354
rect 107282 47302 107334 47354
rect 4874 46758 4926 46810
rect 4938 46758 4990 46810
rect 5002 46758 5054 46810
rect 5066 46758 5118 46810
rect 5130 46758 5182 46810
rect 107762 46758 107814 46810
rect 107826 46758 107878 46810
rect 107890 46758 107942 46810
rect 107954 46758 108006 46810
rect 108018 46758 108070 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 107026 46214 107078 46266
rect 107090 46214 107142 46266
rect 107154 46214 107206 46266
rect 107218 46214 107270 46266
rect 107282 46214 107334 46266
rect 104808 46155 104860 46164
rect 104256 46044 104308 46096
rect 104808 46121 104817 46155
rect 104817 46121 104851 46155
rect 104851 46121 104860 46155
rect 104808 46112 104860 46121
rect 104900 45908 104952 45960
rect 104900 45815 104952 45824
rect 104900 45781 104909 45815
rect 104909 45781 104943 45815
rect 104943 45781 104952 45815
rect 104900 45772 104952 45781
rect 105452 45772 105504 45824
rect 4874 45670 4926 45722
rect 4938 45670 4990 45722
rect 5002 45670 5054 45722
rect 5066 45670 5118 45722
rect 5130 45670 5182 45722
rect 107762 45670 107814 45722
rect 107826 45670 107878 45722
rect 107890 45670 107942 45722
rect 107954 45670 108006 45722
rect 108018 45670 108070 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 107026 45126 107078 45178
rect 107090 45126 107142 45178
rect 107154 45126 107206 45178
rect 107218 45126 107270 45178
rect 107282 45126 107334 45178
rect 104900 45024 104952 45076
rect 104716 44956 104768 45008
rect 105452 44888 105504 44940
rect 105176 44684 105228 44736
rect 105452 44727 105504 44736
rect 105452 44693 105461 44727
rect 105461 44693 105495 44727
rect 105495 44693 105504 44727
rect 105452 44684 105504 44693
rect 4874 44582 4926 44634
rect 4938 44582 4990 44634
rect 5002 44582 5054 44634
rect 5066 44582 5118 44634
rect 5130 44582 5182 44634
rect 107762 44582 107814 44634
rect 107826 44582 107878 44634
rect 107890 44582 107942 44634
rect 107954 44582 108006 44634
rect 108018 44582 108070 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 107026 44038 107078 44090
rect 107090 44038 107142 44090
rect 107154 44038 107206 44090
rect 107218 44038 107270 44090
rect 107282 44038 107334 44090
rect 104532 43936 104584 43988
rect 104532 43732 104584 43784
rect 105084 43664 105136 43716
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 107762 43494 107814 43546
rect 107826 43494 107878 43546
rect 107890 43494 107942 43546
rect 107954 43494 108006 43546
rect 108018 43494 108070 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 107026 42950 107078 43002
rect 107090 42950 107142 43002
rect 107154 42950 107206 43002
rect 107218 42950 107270 43002
rect 107282 42950 107334 43002
rect 104992 42712 105044 42764
rect 104624 42619 104676 42628
rect 104624 42585 104633 42619
rect 104633 42585 104667 42619
rect 104667 42585 104676 42619
rect 104624 42576 104676 42585
rect 105084 42576 105136 42628
rect 104164 42508 104216 42560
rect 105452 42508 105504 42560
rect 106372 42551 106424 42560
rect 106372 42517 106381 42551
rect 106381 42517 106415 42551
rect 106415 42517 106424 42551
rect 106372 42508 106424 42517
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 107762 42406 107814 42458
rect 107826 42406 107878 42458
rect 107890 42406 107942 42458
rect 107954 42406 108006 42458
rect 108018 42406 108070 42458
rect 104992 42168 105044 42220
rect 106096 42168 106148 42220
rect 106096 41964 106148 42016
rect 106372 41964 106424 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 107026 41862 107078 41914
rect 107090 41862 107142 41914
rect 107154 41862 107206 41914
rect 107218 41862 107270 41914
rect 107282 41862 107334 41914
rect 104348 41599 104400 41608
rect 104348 41565 104357 41599
rect 104357 41565 104391 41599
rect 104391 41565 104400 41599
rect 104348 41556 104400 41565
rect 104900 41556 104952 41608
rect 106096 41531 106148 41540
rect 106096 41497 106105 41531
rect 106105 41497 106139 41531
rect 106139 41497 106148 41531
rect 106096 41488 106148 41497
rect 7564 41463 7616 41472
rect 7564 41429 7573 41463
rect 7573 41429 7607 41463
rect 7607 41429 7616 41463
rect 7564 41420 7616 41429
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 107762 41318 107814 41370
rect 107826 41318 107878 41370
rect 107890 41318 107942 41370
rect 107954 41318 108006 41370
rect 108018 41318 108070 41370
rect 104624 41216 104676 41268
rect 104900 41259 104952 41268
rect 104900 41225 104909 41259
rect 104909 41225 104943 41259
rect 104943 41225 104952 41259
rect 104900 41216 104952 41225
rect 104256 41080 104308 41132
rect 105176 40876 105228 40928
rect 105912 40876 105964 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 107026 40774 107078 40826
rect 107090 40774 107142 40826
rect 107154 40774 107206 40826
rect 107218 40774 107270 40826
rect 107282 40774 107334 40826
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 107762 40230 107814 40282
rect 107826 40230 107878 40282
rect 107890 40230 107942 40282
rect 107954 40230 108006 40282
rect 108018 40230 108070 40282
rect 7564 39831 7616 39840
rect 7564 39797 7573 39831
rect 7573 39797 7607 39831
rect 7607 39797 7616 39831
rect 7564 39788 7616 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 107026 39686 107078 39738
rect 107090 39686 107142 39738
rect 107154 39686 107206 39738
rect 107218 39686 107270 39738
rect 107282 39686 107334 39738
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 107762 39142 107814 39194
rect 107826 39142 107878 39194
rect 107890 39142 107942 39194
rect 107954 39142 108006 39194
rect 108018 39142 108070 39194
rect 7564 38743 7616 38752
rect 7564 38709 7573 38743
rect 7573 38709 7607 38743
rect 7607 38709 7616 38743
rect 7564 38700 7616 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 107026 38598 107078 38650
rect 107090 38598 107142 38650
rect 107154 38598 107206 38650
rect 107218 38598 107270 38650
rect 107282 38598 107334 38650
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 107762 38054 107814 38106
rect 107826 38054 107878 38106
rect 107890 38054 107942 38106
rect 107954 38054 108006 38106
rect 108018 38054 108070 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 107026 37510 107078 37562
rect 107090 37510 107142 37562
rect 107154 37510 107206 37562
rect 107218 37510 107270 37562
rect 107282 37510 107334 37562
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 107762 36966 107814 37018
rect 107826 36966 107878 37018
rect 107890 36966 107942 37018
rect 107954 36966 108006 37018
rect 108018 36966 108070 37018
rect 104532 36864 104584 36916
rect 7564 36771 7616 36780
rect 7564 36737 7573 36771
rect 7573 36737 7607 36771
rect 7607 36737 7616 36771
rect 7564 36728 7616 36737
rect 104532 36524 104584 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 107026 36422 107078 36474
rect 107090 36422 107142 36474
rect 107154 36422 107206 36474
rect 107218 36422 107270 36474
rect 107282 36422 107334 36474
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 107762 35878 107814 35930
rect 107826 35878 107878 35930
rect 107890 35878 107942 35930
rect 107954 35878 108006 35930
rect 108018 35878 108070 35930
rect 104716 35640 104768 35692
rect 7564 35547 7616 35556
rect 7564 35513 7573 35547
rect 7573 35513 7607 35547
rect 7607 35513 7616 35547
rect 7564 35504 7616 35513
rect 104440 35479 104492 35488
rect 104440 35445 104449 35479
rect 104449 35445 104483 35479
rect 104483 35445 104492 35479
rect 104440 35436 104492 35445
rect 104716 35479 104768 35488
rect 104716 35445 104725 35479
rect 104725 35445 104759 35479
rect 104759 35445 104768 35479
rect 104716 35436 104768 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 107026 35334 107078 35386
rect 107090 35334 107142 35386
rect 107154 35334 107206 35386
rect 107218 35334 107270 35386
rect 107282 35334 107334 35386
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 107762 34790 107814 34842
rect 107826 34790 107878 34842
rect 107890 34790 107942 34842
rect 107954 34790 108006 34842
rect 108018 34790 108070 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 107026 34246 107078 34298
rect 107090 34246 107142 34298
rect 107154 34246 107206 34298
rect 107218 34246 107270 34298
rect 107282 34246 107334 34298
rect 7564 34051 7616 34060
rect 7564 34017 7573 34051
rect 7573 34017 7607 34051
rect 7607 34017 7616 34051
rect 7564 34008 7616 34017
rect 106096 33983 106148 33992
rect 106096 33949 106105 33983
rect 106105 33949 106139 33983
rect 106139 33949 106148 33983
rect 106096 33940 106148 33949
rect 104532 33872 104584 33924
rect 105820 33915 105872 33924
rect 105820 33881 105829 33915
rect 105829 33881 105863 33915
rect 105863 33881 105872 33915
rect 105820 33872 105872 33881
rect 104808 33804 104860 33856
rect 106188 33847 106240 33856
rect 106188 33813 106197 33847
rect 106197 33813 106231 33847
rect 106231 33813 106240 33847
rect 106188 33804 106240 33813
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 107762 33702 107814 33754
rect 107826 33702 107878 33754
rect 107890 33702 107942 33754
rect 107954 33702 108006 33754
rect 108018 33702 108070 33754
rect 104808 33439 104860 33448
rect 104808 33405 104817 33439
rect 104817 33405 104851 33439
rect 104851 33405 104860 33439
rect 104808 33396 104860 33405
rect 105636 33260 105688 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 107026 33158 107078 33210
rect 107090 33158 107142 33210
rect 107154 33158 107206 33210
rect 107218 33158 107270 33210
rect 107282 33158 107334 33210
rect 105452 32920 105504 32972
rect 106188 32852 106240 32904
rect 104440 32784 104492 32836
rect 104532 32716 104584 32768
rect 106372 32716 106424 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 107762 32614 107814 32666
rect 107826 32614 107878 32666
rect 107890 32614 107942 32666
rect 107954 32614 108006 32666
rect 108018 32614 108070 32666
rect 110328 32376 110380 32428
rect 104532 32351 104584 32360
rect 104532 32317 104541 32351
rect 104541 32317 104575 32351
rect 104575 32317 104584 32351
rect 104532 32308 104584 32317
rect 104716 32308 104768 32360
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 107026 32070 107078 32122
rect 107090 32070 107142 32122
rect 107154 32070 107206 32122
rect 107218 32070 107270 32122
rect 107282 32070 107334 32122
rect 105820 31968 105872 32020
rect 110328 32011 110380 32020
rect 110328 31977 110337 32011
rect 110337 31977 110371 32011
rect 110371 31977 110380 32011
rect 110328 31968 110380 31977
rect 104716 31900 104768 31952
rect 105912 31900 105964 31952
rect 104532 31764 104584 31816
rect 104624 31764 104676 31816
rect 105360 31807 105412 31816
rect 105360 31773 105369 31807
rect 105369 31773 105403 31807
rect 105403 31773 105412 31807
rect 105360 31764 105412 31773
rect 105636 31807 105688 31816
rect 105636 31773 105645 31807
rect 105645 31773 105679 31807
rect 105679 31773 105688 31807
rect 105636 31764 105688 31773
rect 110512 31807 110564 31816
rect 110512 31773 110521 31807
rect 110521 31773 110555 31807
rect 110555 31773 110564 31807
rect 110512 31764 110564 31773
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 107762 31526 107814 31578
rect 107826 31526 107878 31578
rect 107890 31526 107942 31578
rect 107954 31526 108006 31578
rect 108018 31526 108070 31578
rect 104532 31084 104584 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 107026 30982 107078 31034
rect 107090 30982 107142 31034
rect 107154 30982 107206 31034
rect 107218 30982 107270 31034
rect 107282 30982 107334 31034
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 107762 30438 107814 30490
rect 107826 30438 107878 30490
rect 107890 30438 107942 30490
rect 107954 30438 108006 30490
rect 108018 30438 108070 30490
rect 104440 30268 104492 30320
rect 104808 30268 104860 30320
rect 105360 30200 105412 30252
rect 105912 30268 105964 30320
rect 105452 30064 105504 30116
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 107026 29894 107078 29946
rect 107090 29894 107142 29946
rect 107154 29894 107206 29946
rect 107218 29894 107270 29946
rect 107282 29894 107334 29946
rect 104532 29588 104584 29640
rect 104256 29452 104308 29504
rect 104808 29452 104860 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 107762 29350 107814 29402
rect 107826 29350 107878 29402
rect 107890 29350 107942 29402
rect 107954 29350 108006 29402
rect 108018 29350 108070 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 107026 28806 107078 28858
rect 107090 28806 107142 28858
rect 107154 28806 107206 28858
rect 107218 28806 107270 28858
rect 107282 28806 107334 28858
rect 106372 28568 106424 28620
rect 104532 28432 104584 28484
rect 104716 28432 104768 28484
rect 105452 28364 105504 28416
rect 106372 28364 106424 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 107762 28262 107814 28314
rect 107826 28262 107878 28314
rect 107890 28262 107942 28314
rect 107954 28262 108006 28314
rect 108018 28262 108070 28314
rect 104440 28092 104492 28144
rect 105084 28092 105136 28144
rect 105912 28092 105964 28144
rect 104716 27820 104768 27872
rect 105176 27863 105228 27872
rect 105176 27829 105185 27863
rect 105185 27829 105219 27863
rect 105219 27829 105228 27863
rect 105176 27820 105228 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 107026 27718 107078 27770
rect 107090 27718 107142 27770
rect 107154 27718 107206 27770
rect 107218 27718 107270 27770
rect 107282 27718 107334 27770
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 107762 27174 107814 27226
rect 107826 27174 107878 27226
rect 107890 27174 107942 27226
rect 107954 27174 108006 27226
rect 108018 27174 108070 27226
rect 104532 27072 104584 27124
rect 104716 27072 104768 27124
rect 105084 27072 105136 27124
rect 105452 27115 105504 27124
rect 105452 27081 105461 27115
rect 105461 27081 105495 27115
rect 105495 27081 105504 27115
rect 105452 27072 105504 27081
rect 105268 27004 105320 27056
rect 105176 26936 105228 26988
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 107026 26630 107078 26682
rect 107090 26630 107142 26682
rect 107154 26630 107206 26682
rect 107218 26630 107270 26682
rect 107282 26630 107334 26682
rect 104348 26256 104400 26308
rect 106372 26256 106424 26308
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 107762 26086 107814 26138
rect 107826 26086 107878 26138
rect 107890 26086 107942 26138
rect 107954 26086 108006 26138
rect 108018 26086 108070 26138
rect 104256 25916 104308 25968
rect 104348 25891 104400 25900
rect 104348 25857 104357 25891
rect 104357 25857 104391 25891
rect 104391 25857 104400 25891
rect 104348 25848 104400 25857
rect 104624 25823 104676 25832
rect 104624 25789 104633 25823
rect 104633 25789 104667 25823
rect 104667 25789 104676 25823
rect 104624 25780 104676 25789
rect 105268 25644 105320 25696
rect 106372 25687 106424 25696
rect 106372 25653 106381 25687
rect 106381 25653 106415 25687
rect 106415 25653 106424 25687
rect 106372 25644 106424 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 107026 25542 107078 25594
rect 107090 25542 107142 25594
rect 107154 25542 107206 25594
rect 107218 25542 107270 25594
rect 107282 25542 107334 25594
rect 104532 25483 104584 25492
rect 104532 25449 104541 25483
rect 104541 25449 104575 25483
rect 104575 25449 104584 25483
rect 104532 25440 104584 25449
rect 104716 25483 104768 25492
rect 104716 25449 104725 25483
rect 104725 25449 104759 25483
rect 104759 25449 104768 25483
rect 104716 25440 104768 25449
rect 104808 25279 104860 25288
rect 104808 25245 104817 25279
rect 104817 25245 104851 25279
rect 104851 25245 104860 25279
rect 104808 25236 104860 25245
rect 104348 25211 104400 25220
rect 104348 25177 104357 25211
rect 104357 25177 104391 25211
rect 104391 25177 104400 25211
rect 104348 25168 104400 25177
rect 104256 25100 104308 25152
rect 105176 25168 105228 25220
rect 104900 25143 104952 25152
rect 104900 25109 104909 25143
rect 104909 25109 104943 25143
rect 104943 25109 104952 25143
rect 104900 25100 104952 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 107762 24998 107814 25050
rect 107826 24998 107878 25050
rect 107890 24998 107942 25050
rect 107954 24998 108006 25050
rect 108018 24998 108070 25050
rect 104164 24760 104216 24812
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 107026 24454 107078 24506
rect 107090 24454 107142 24506
rect 107154 24454 107206 24506
rect 107218 24454 107270 24506
rect 107282 24454 107334 24506
rect 104992 24352 105044 24404
rect 104716 24148 104768 24200
rect 104164 24080 104216 24132
rect 105268 24080 105320 24132
rect 104440 24055 104492 24064
rect 104440 24021 104455 24055
rect 104455 24021 104489 24055
rect 104489 24021 104492 24055
rect 104440 24012 104492 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 107762 23910 107814 23962
rect 107826 23910 107878 23962
rect 107890 23910 107942 23962
rect 107954 23910 108006 23962
rect 108018 23910 108070 23962
rect 104716 23808 104768 23860
rect 104992 23808 105044 23860
rect 105268 23851 105320 23860
rect 105268 23817 105277 23851
rect 105277 23817 105311 23851
rect 105311 23817 105320 23851
rect 105268 23808 105320 23817
rect 104164 23740 104216 23792
rect 104440 23672 104492 23724
rect 104624 23536 104676 23588
rect 104716 23511 104768 23520
rect 104716 23477 104725 23511
rect 104725 23477 104759 23511
rect 104759 23477 104768 23511
rect 104716 23468 104768 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 107026 23366 107078 23418
rect 107090 23366 107142 23418
rect 107154 23366 107206 23418
rect 107218 23366 107270 23418
rect 107282 23366 107334 23418
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 107762 22822 107814 22874
rect 107826 22822 107878 22874
rect 107890 22822 107942 22874
rect 107954 22822 108006 22874
rect 108018 22822 108070 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 107026 22278 107078 22330
rect 107090 22278 107142 22330
rect 107154 22278 107206 22330
rect 107218 22278 107270 22330
rect 107282 22278 107334 22330
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 107762 21734 107814 21786
rect 107826 21734 107878 21786
rect 107890 21734 107942 21786
rect 107954 21734 108006 21786
rect 108018 21734 108070 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 107026 21190 107078 21242
rect 107090 21190 107142 21242
rect 107154 21190 107206 21242
rect 107218 21190 107270 21242
rect 107282 21190 107334 21242
rect 106372 20995 106424 21004
rect 106372 20961 106381 20995
rect 106381 20961 106415 20995
rect 106415 20961 106424 20995
rect 106372 20952 106424 20961
rect 104348 20816 104400 20868
rect 104900 20816 104952 20868
rect 106096 20791 106148 20800
rect 106096 20757 106105 20791
rect 106105 20757 106139 20791
rect 106139 20757 106148 20791
rect 106096 20748 106148 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 107762 20646 107814 20698
rect 107826 20646 107878 20698
rect 107890 20646 107942 20698
rect 107954 20646 108006 20698
rect 108018 20646 108070 20698
rect 104256 20340 104308 20392
rect 106096 20340 106148 20392
rect 104716 20204 104768 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 107026 20102 107078 20154
rect 107090 20102 107142 20154
rect 107154 20102 107206 20154
rect 107218 20102 107270 20154
rect 107282 20102 107334 20154
rect 104256 19660 104308 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 107762 19558 107814 19610
rect 107826 19558 107878 19610
rect 107890 19558 107942 19610
rect 107954 19558 108006 19610
rect 108018 19558 108070 19610
rect 104716 19363 104768 19372
rect 104716 19329 104725 19363
rect 104725 19329 104759 19363
rect 104759 19329 104768 19363
rect 104716 19320 104768 19329
rect 104348 19295 104400 19304
rect 104348 19261 104357 19295
rect 104357 19261 104391 19295
rect 104391 19261 104400 19295
rect 104348 19252 104400 19261
rect 104624 19295 104676 19304
rect 104624 19261 104633 19295
rect 104633 19261 104667 19295
rect 104667 19261 104676 19295
rect 104624 19252 104676 19261
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 107026 19014 107078 19066
rect 107090 19014 107142 19066
rect 107154 19014 107206 19066
rect 107218 19014 107270 19066
rect 107282 19014 107334 19066
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 107762 18470 107814 18522
rect 107826 18470 107878 18522
rect 107890 18470 107942 18522
rect 107954 18470 108006 18522
rect 108018 18470 108070 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 107026 17926 107078 17978
rect 107090 17926 107142 17978
rect 107154 17926 107206 17978
rect 107218 17926 107270 17978
rect 107282 17926 107334 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 107762 17382 107814 17434
rect 107826 17382 107878 17434
rect 107890 17382 107942 17434
rect 107954 17382 108006 17434
rect 108018 17382 108070 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 107026 16838 107078 16890
rect 107090 16838 107142 16890
rect 107154 16838 107206 16890
rect 107218 16838 107270 16890
rect 107282 16838 107334 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 107762 16294 107814 16346
rect 107826 16294 107878 16346
rect 107890 16294 107942 16346
rect 107954 16294 108006 16346
rect 108018 16294 108070 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 107026 15750 107078 15802
rect 107090 15750 107142 15802
rect 107154 15750 107206 15802
rect 107218 15750 107270 15802
rect 107282 15750 107334 15802
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 7564 15512 7616 15521
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 107762 15206 107814 15258
rect 107826 15206 107878 15258
rect 107890 15206 107942 15258
rect 107954 15206 108006 15258
rect 108018 15206 108070 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 107026 14662 107078 14714
rect 107090 14662 107142 14714
rect 107154 14662 107206 14714
rect 107218 14662 107270 14714
rect 107282 14662 107334 14714
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 107762 14118 107814 14170
rect 107826 14118 107878 14170
rect 107890 14118 107942 14170
rect 107954 14118 108006 14170
rect 108018 14118 108070 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 107026 13574 107078 13626
rect 107090 13574 107142 13626
rect 107154 13574 107206 13626
rect 107218 13574 107270 13626
rect 107282 13574 107334 13626
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 107762 13030 107814 13082
rect 107826 13030 107878 13082
rect 107890 13030 107942 13082
rect 107954 13030 108006 13082
rect 108018 13030 108070 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 107026 12486 107078 12538
rect 107090 12486 107142 12538
rect 107154 12486 107206 12538
rect 107218 12486 107270 12538
rect 107282 12486 107334 12538
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 107762 11942 107814 11994
rect 107826 11942 107878 11994
rect 107890 11942 107942 11994
rect 107954 11942 108006 11994
rect 108018 11942 108070 11994
rect 102784 11704 102836 11756
rect 110420 11704 110472 11756
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 107026 11398 107078 11450
rect 107090 11398 107142 11450
rect 107154 11398 107206 11450
rect 107218 11398 107270 11450
rect 107282 11398 107334 11450
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 107762 10854 107814 10906
rect 107826 10854 107878 10906
rect 107890 10854 107942 10906
rect 107954 10854 108006 10906
rect 108018 10854 108070 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 107026 10310 107078 10362
rect 107090 10310 107142 10362
rect 107154 10310 107206 10362
rect 107218 10310 107270 10362
rect 107282 10310 107334 10362
rect 90364 10004 90416 10056
rect 104440 10004 104492 10056
rect 90732 9936 90784 9988
rect 104164 9936 104216 9988
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 107762 9766 107814 9818
rect 107826 9766 107878 9818
rect 107890 9766 107942 9818
rect 107954 9766 108006 9818
rect 108018 9766 108070 9818
rect 8208 9596 8260 9648
rect 16028 9596 16080 9648
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 107026 9222 107078 9274
rect 107090 9222 107142 9274
rect 107154 9222 107206 9274
rect 107218 9222 107270 9274
rect 107282 9222 107334 9274
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 107762 8678 107814 8730
rect 107826 8678 107878 8730
rect 107890 8678 107942 8730
rect 107954 8678 108006 8730
rect 108018 8678 108070 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 107026 8134 107078 8186
rect 107090 8134 107142 8186
rect 107154 8134 107206 8186
rect 107218 8134 107270 8186
rect 107282 8134 107334 8186
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 66314 7590 66366 7642
rect 66378 7590 66430 7642
rect 66442 7590 66494 7642
rect 66506 7590 66558 7642
rect 66570 7590 66622 7642
rect 97034 7590 97086 7642
rect 97098 7590 97150 7642
rect 97162 7590 97214 7642
rect 97226 7590 97278 7642
rect 97290 7590 97342 7642
rect 107762 7590 107814 7642
rect 107826 7590 107878 7642
rect 107890 7590 107942 7642
rect 107954 7590 108006 7642
rect 108018 7590 108070 7642
rect 16028 7488 16080 7540
rect 23204 7488 23256 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 25780 7488 25832 7540
rect 26976 7531 27028 7540
rect 26976 7497 26985 7531
rect 26985 7497 27019 7531
rect 27019 7497 27028 7531
rect 26976 7488 27028 7497
rect 28264 7531 28316 7540
rect 28264 7497 28273 7531
rect 28273 7497 28307 7531
rect 28307 7497 28316 7531
rect 28264 7488 28316 7497
rect 29000 7488 29052 7540
rect 30472 7531 30524 7540
rect 30472 7497 30481 7531
rect 30481 7497 30515 7531
rect 30515 7497 30524 7531
rect 30472 7488 30524 7497
rect 31576 7488 31628 7540
rect 32864 7531 32916 7540
rect 32864 7497 32873 7531
rect 32873 7497 32907 7531
rect 32907 7497 32916 7531
rect 32864 7488 32916 7497
rect 33968 7531 34020 7540
rect 33968 7497 33977 7531
rect 33977 7497 34011 7531
rect 34011 7497 34020 7531
rect 33968 7488 34020 7497
rect 35256 7531 35308 7540
rect 35256 7497 35265 7531
rect 35265 7497 35299 7531
rect 35299 7497 35308 7531
rect 35256 7488 35308 7497
rect 36084 7488 36136 7540
rect 36360 7531 36412 7540
rect 36360 7497 36369 7531
rect 36369 7497 36403 7531
rect 36403 7497 36412 7531
rect 36360 7488 36412 7497
rect 37464 7531 37516 7540
rect 37464 7497 37473 7531
rect 37473 7497 37507 7531
rect 37507 7497 37516 7531
rect 37464 7488 37516 7497
rect 38660 7531 38712 7540
rect 38660 7497 38669 7531
rect 38669 7497 38703 7531
rect 38703 7497 38712 7531
rect 38660 7488 38712 7497
rect 39856 7531 39908 7540
rect 39856 7497 39865 7531
rect 39865 7497 39899 7531
rect 39899 7497 39908 7531
rect 39856 7488 39908 7497
rect 41052 7531 41104 7540
rect 41052 7497 41061 7531
rect 41061 7497 41095 7531
rect 41095 7497 41104 7531
rect 41052 7488 41104 7497
rect 41880 7488 41932 7540
rect 42156 7531 42208 7540
rect 42156 7497 42165 7531
rect 42165 7497 42199 7531
rect 42199 7497 42208 7531
rect 42156 7488 42208 7497
rect 43352 7531 43404 7540
rect 43352 7497 43361 7531
rect 43361 7497 43395 7531
rect 43395 7497 43404 7531
rect 43352 7488 43404 7497
rect 90548 7531 90600 7540
rect 90548 7497 90557 7531
rect 90557 7497 90591 7531
rect 90591 7497 90600 7531
rect 90548 7488 90600 7497
rect 90732 7531 90784 7540
rect 90732 7497 90741 7531
rect 90741 7497 90775 7531
rect 90775 7497 90784 7531
rect 90732 7488 90784 7497
rect 91008 7531 91060 7540
rect 91008 7497 91017 7531
rect 91017 7497 91051 7531
rect 91051 7497 91060 7531
rect 91008 7488 91060 7497
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 107026 7046 107078 7098
rect 107090 7046 107142 7098
rect 107154 7046 107206 7098
rect 107218 7046 107270 7098
rect 107282 7046 107334 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 66314 6502 66366 6554
rect 66378 6502 66430 6554
rect 66442 6502 66494 6554
rect 66506 6502 66558 6554
rect 66570 6502 66622 6554
rect 97034 6502 97086 6554
rect 97098 6502 97150 6554
rect 97162 6502 97214 6554
rect 97226 6502 97278 6554
rect 97290 6502 97342 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 66314 5414 66366 5466
rect 66378 5414 66430 5466
rect 66442 5414 66494 5466
rect 66506 5414 66558 5466
rect 66570 5414 66622 5466
rect 97034 5414 97086 5466
rect 97098 5414 97150 5466
rect 97162 5414 97214 5466
rect 97226 5414 97278 5466
rect 97290 5414 97342 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 66314 4326 66366 4378
rect 66378 4326 66430 4378
rect 66442 4326 66494 4378
rect 66506 4326 66558 4378
rect 66570 4326 66622 4378
rect 97034 4326 97086 4378
rect 97098 4326 97150 4378
rect 97162 4326 97214 4378
rect 97226 4326 97278 4378
rect 97290 4326 97342 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 66314 3238 66366 3290
rect 66378 3238 66430 3290
rect 66442 3238 66494 3290
rect 66506 3238 66558 3290
rect 66570 3238 66622 3290
rect 97034 3238 97086 3290
rect 97098 3238 97150 3290
rect 97162 3238 97214 3290
rect 97226 3238 97278 3290
rect 97290 3238 97342 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 66314 2150 66366 2202
rect 66378 2150 66430 2202
rect 66442 2150 66494 2202
rect 66506 2150 66558 2202
rect 66570 2150 66622 2202
rect 97034 2150 97086 2202
rect 97098 2150 97150 2202
rect 97162 2150 97214 2202
rect 97226 2150 97278 2202
rect 97290 2150 97342 2202
<< metal2 >>
rect 44454 73200 44510 74000
rect 47030 73200 47086 74000
rect 49606 73200 49662 74000
rect 51538 73200 51594 74000
rect 53470 73200 53526 74000
rect 55402 73200 55458 74000
rect 57334 73200 57390 74000
rect 59266 73200 59322 74000
rect 61198 73200 61254 74000
rect 63130 73200 63186 74000
rect 65706 73200 65762 74000
rect 67638 73200 67694 74000
rect 69570 73200 69626 74000
rect 71502 73200 71558 74000
rect 74078 73200 74134 74000
rect 77298 73200 77354 74000
rect 4874 71836 5182 71845
rect 4874 71834 4880 71836
rect 4936 71834 4960 71836
rect 5016 71834 5040 71836
rect 5096 71834 5120 71836
rect 5176 71834 5182 71836
rect 4936 71782 4938 71834
rect 5118 71782 5120 71834
rect 4874 71780 4880 71782
rect 4936 71780 4960 71782
rect 5016 71780 5040 71782
rect 5096 71780 5120 71782
rect 5176 71780 5182 71782
rect 4874 71771 5182 71780
rect 35594 71836 35902 71845
rect 35594 71834 35600 71836
rect 35656 71834 35680 71836
rect 35736 71834 35760 71836
rect 35816 71834 35840 71836
rect 35896 71834 35902 71836
rect 35656 71782 35658 71834
rect 35838 71782 35840 71834
rect 35594 71780 35600 71782
rect 35656 71780 35680 71782
rect 35736 71780 35760 71782
rect 35816 71780 35840 71782
rect 35896 71780 35902 71782
rect 35594 71771 35902 71780
rect 44468 71738 44496 73200
rect 47044 71738 47072 73200
rect 49620 71738 49648 73200
rect 51552 71738 51580 73200
rect 53484 71738 53512 73200
rect 55416 71738 55444 73200
rect 57348 71738 57376 73200
rect 59280 71738 59308 73200
rect 61212 71738 61240 73200
rect 63144 71738 63172 73200
rect 65720 71738 65748 73200
rect 66314 71836 66622 71845
rect 66314 71834 66320 71836
rect 66376 71834 66400 71836
rect 66456 71834 66480 71836
rect 66536 71834 66560 71836
rect 66616 71834 66622 71836
rect 66376 71782 66378 71834
rect 66558 71782 66560 71834
rect 66314 71780 66320 71782
rect 66376 71780 66400 71782
rect 66456 71780 66480 71782
rect 66536 71780 66560 71782
rect 66616 71780 66622 71782
rect 66314 71771 66622 71780
rect 67652 71738 67680 73200
rect 69584 71738 69612 73200
rect 71516 71738 71544 73200
rect 74092 71738 74120 73200
rect 77312 71738 77340 73200
rect 97034 71836 97342 71845
rect 97034 71834 97040 71836
rect 97096 71834 97120 71836
rect 97176 71834 97200 71836
rect 97256 71834 97280 71836
rect 97336 71834 97342 71836
rect 97096 71782 97098 71834
rect 97278 71782 97280 71834
rect 97034 71780 97040 71782
rect 97096 71780 97120 71782
rect 97176 71780 97200 71782
rect 97256 71780 97280 71782
rect 97336 71780 97342 71782
rect 97034 71771 97342 71780
rect 44456 71732 44508 71738
rect 44456 71674 44508 71680
rect 47032 71732 47084 71738
rect 47032 71674 47084 71680
rect 49608 71732 49660 71738
rect 49608 71674 49660 71680
rect 51540 71732 51592 71738
rect 51540 71674 51592 71680
rect 53472 71732 53524 71738
rect 53472 71674 53524 71680
rect 55404 71732 55456 71738
rect 55404 71674 55456 71680
rect 57336 71732 57388 71738
rect 57336 71674 57388 71680
rect 59268 71732 59320 71738
rect 59268 71674 59320 71680
rect 61200 71732 61252 71738
rect 61200 71674 61252 71680
rect 63132 71732 63184 71738
rect 63132 71674 63184 71680
rect 65708 71732 65760 71738
rect 65708 71674 65760 71680
rect 67640 71732 67692 71738
rect 67640 71674 67692 71680
rect 69572 71732 69624 71738
rect 69572 71674 69624 71680
rect 71504 71732 71556 71738
rect 71504 71674 71556 71680
rect 74080 71732 74132 71738
rect 74080 71674 74132 71680
rect 77300 71732 77352 71738
rect 77300 71674 77352 71680
rect 45100 71596 45152 71602
rect 45100 71538 45152 71544
rect 47308 71596 47360 71602
rect 47308 71538 47360 71544
rect 49516 71596 49568 71602
rect 49516 71538 49568 71544
rect 51632 71596 51684 71602
rect 51632 71538 51684 71544
rect 53564 71596 53616 71602
rect 53564 71538 53616 71544
rect 55496 71596 55548 71602
rect 55496 71538 55548 71544
rect 57428 71596 57480 71602
rect 57428 71538 57480 71544
rect 59636 71596 59688 71602
rect 59636 71538 59688 71544
rect 61568 71596 61620 71602
rect 61568 71538 61620 71544
rect 63132 71596 63184 71602
rect 63132 71538 63184 71544
rect 65432 71596 65484 71602
rect 65432 71538 65484 71544
rect 67364 71596 67416 71602
rect 67364 71538 67416 71544
rect 69940 71596 69992 71602
rect 69940 71538 69992 71544
rect 71872 71596 71924 71602
rect 71872 71538 71924 71544
rect 74172 71596 74224 71602
rect 74172 71538 74224 71544
rect 76104 71596 76156 71602
rect 76104 71538 76156 71544
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 34934 71292 35242 71301
rect 34934 71290 34940 71292
rect 34996 71290 35020 71292
rect 35076 71290 35100 71292
rect 35156 71290 35180 71292
rect 35236 71290 35242 71292
rect 34996 71238 34998 71290
rect 35178 71238 35180 71290
rect 34934 71236 34940 71238
rect 34996 71236 35020 71238
rect 35076 71236 35100 71238
rect 35156 71236 35180 71238
rect 35236 71236 35242 71238
rect 34934 71227 35242 71236
rect 4874 70748 5182 70757
rect 4874 70746 4880 70748
rect 4936 70746 4960 70748
rect 5016 70746 5040 70748
rect 5096 70746 5120 70748
rect 5176 70746 5182 70748
rect 4936 70694 4938 70746
rect 5118 70694 5120 70746
rect 4874 70692 4880 70694
rect 4936 70692 4960 70694
rect 5016 70692 5040 70694
rect 5096 70692 5120 70694
rect 5176 70692 5182 70694
rect 4874 70683 5182 70692
rect 35594 70748 35902 70757
rect 35594 70746 35600 70748
rect 35656 70746 35680 70748
rect 35736 70746 35760 70748
rect 35816 70746 35840 70748
rect 35896 70746 35902 70748
rect 35656 70694 35658 70746
rect 35838 70694 35840 70746
rect 35594 70692 35600 70694
rect 35656 70692 35680 70694
rect 35736 70692 35760 70694
rect 35816 70692 35840 70694
rect 35896 70692 35902 70694
rect 35594 70683 35902 70692
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70139 4522 70148
rect 34934 70204 35242 70213
rect 34934 70202 34940 70204
rect 34996 70202 35020 70204
rect 35076 70202 35100 70204
rect 35156 70202 35180 70204
rect 35236 70202 35242 70204
rect 34996 70150 34998 70202
rect 35178 70150 35180 70202
rect 34934 70148 34940 70150
rect 34996 70148 35020 70150
rect 35076 70148 35100 70150
rect 35156 70148 35180 70150
rect 35236 70148 35242 70150
rect 34934 70139 35242 70148
rect 4874 69660 5182 69669
rect 4874 69658 4880 69660
rect 4936 69658 4960 69660
rect 5016 69658 5040 69660
rect 5096 69658 5120 69660
rect 5176 69658 5182 69660
rect 4936 69606 4938 69658
rect 5118 69606 5120 69658
rect 4874 69604 4880 69606
rect 4936 69604 4960 69606
rect 5016 69604 5040 69606
rect 5096 69604 5120 69606
rect 5176 69604 5182 69606
rect 4874 69595 5182 69604
rect 35594 69660 35902 69669
rect 35594 69658 35600 69660
rect 35656 69658 35680 69660
rect 35736 69658 35760 69660
rect 35816 69658 35840 69660
rect 35896 69658 35902 69660
rect 35656 69606 35658 69658
rect 35838 69606 35840 69658
rect 35594 69604 35600 69606
rect 35656 69604 35680 69606
rect 35736 69604 35760 69606
rect 35816 69604 35840 69606
rect 35896 69604 35902 69606
rect 35594 69595 35902 69604
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 34934 69116 35242 69125
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69051 35242 69060
rect 4874 68572 5182 68581
rect 4874 68570 4880 68572
rect 4936 68570 4960 68572
rect 5016 68570 5040 68572
rect 5096 68570 5120 68572
rect 5176 68570 5182 68572
rect 4936 68518 4938 68570
rect 5118 68518 5120 68570
rect 4874 68516 4880 68518
rect 4936 68516 4960 68518
rect 5016 68516 5040 68518
rect 5096 68516 5120 68518
rect 5176 68516 5182 68518
rect 4874 68507 5182 68516
rect 35594 68572 35902 68581
rect 35594 68570 35600 68572
rect 35656 68570 35680 68572
rect 35736 68570 35760 68572
rect 35816 68570 35840 68572
rect 35896 68570 35902 68572
rect 35656 68518 35658 68570
rect 35838 68518 35840 68570
rect 35594 68516 35600 68518
rect 35656 68516 35680 68518
rect 35736 68516 35760 68518
rect 35816 68516 35840 68518
rect 35896 68516 35902 68518
rect 35594 68507 35902 68516
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 34934 68028 35242 68037
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67963 35242 67972
rect 4874 67484 5182 67493
rect 4874 67482 4880 67484
rect 4936 67482 4960 67484
rect 5016 67482 5040 67484
rect 5096 67482 5120 67484
rect 5176 67482 5182 67484
rect 4936 67430 4938 67482
rect 5118 67430 5120 67482
rect 4874 67428 4880 67430
rect 4936 67428 4960 67430
rect 5016 67428 5040 67430
rect 5096 67428 5120 67430
rect 5176 67428 5182 67430
rect 4874 67419 5182 67428
rect 35594 67484 35902 67493
rect 35594 67482 35600 67484
rect 35656 67482 35680 67484
rect 35736 67482 35760 67484
rect 35816 67482 35840 67484
rect 35896 67482 35902 67484
rect 35656 67430 35658 67482
rect 35838 67430 35840 67482
rect 35594 67428 35600 67430
rect 35656 67428 35680 67430
rect 35736 67428 35760 67430
rect 35816 67428 35840 67430
rect 35896 67428 35902 67430
rect 35594 67419 35902 67428
rect 44732 67244 44784 67250
rect 44732 67186 44784 67192
rect 8208 67176 8260 67182
rect 8208 67118 8260 67124
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 4874 66396 5182 66405
rect 4874 66394 4880 66396
rect 4936 66394 4960 66396
rect 5016 66394 5040 66396
rect 5096 66394 5120 66396
rect 5176 66394 5182 66396
rect 4936 66342 4938 66394
rect 5118 66342 5120 66394
rect 4874 66340 4880 66342
rect 4936 66340 4960 66342
rect 5016 66340 5040 66342
rect 5096 66340 5120 66342
rect 5176 66340 5182 66342
rect 4874 66331 5182 66340
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 4874 65308 5182 65317
rect 4874 65306 4880 65308
rect 4936 65306 4960 65308
rect 5016 65306 5040 65308
rect 5096 65306 5120 65308
rect 5176 65306 5182 65308
rect 4936 65254 4938 65306
rect 5118 65254 5120 65306
rect 4874 65252 4880 65254
rect 4936 65252 4960 65254
rect 5016 65252 5040 65254
rect 5096 65252 5120 65254
rect 5176 65252 5182 65254
rect 4874 65243 5182 65252
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 4874 64220 5182 64229
rect 4874 64218 4880 64220
rect 4936 64218 4960 64220
rect 5016 64218 5040 64220
rect 5096 64218 5120 64220
rect 5176 64218 5182 64220
rect 4936 64166 4938 64218
rect 5118 64166 5120 64218
rect 4874 64164 4880 64166
rect 4936 64164 4960 64166
rect 5016 64164 5040 64166
rect 5096 64164 5120 64166
rect 5176 64164 5182 64166
rect 4874 64155 5182 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 4874 63132 5182 63141
rect 4874 63130 4880 63132
rect 4936 63130 4960 63132
rect 5016 63130 5040 63132
rect 5096 63130 5120 63132
rect 5176 63130 5182 63132
rect 4936 63078 4938 63130
rect 5118 63078 5120 63130
rect 4874 63076 4880 63078
rect 4936 63076 4960 63078
rect 5016 63076 5040 63078
rect 5096 63076 5120 63078
rect 5176 63076 5182 63078
rect 4874 63067 5182 63076
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 4874 62044 5182 62053
rect 4874 62042 4880 62044
rect 4936 62042 4960 62044
rect 5016 62042 5040 62044
rect 5096 62042 5120 62044
rect 5176 62042 5182 62044
rect 4936 61990 4938 62042
rect 5118 61990 5120 62042
rect 4874 61988 4880 61990
rect 4936 61988 4960 61990
rect 5016 61988 5040 61990
rect 5096 61988 5120 61990
rect 5176 61988 5182 61990
rect 4874 61979 5182 61988
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4874 60956 5182 60965
rect 4874 60954 4880 60956
rect 4936 60954 4960 60956
rect 5016 60954 5040 60956
rect 5096 60954 5120 60956
rect 5176 60954 5182 60956
rect 4936 60902 4938 60954
rect 5118 60902 5120 60954
rect 4874 60900 4880 60902
rect 4936 60900 4960 60902
rect 5016 60900 5040 60902
rect 5096 60900 5120 60902
rect 5176 60900 5182 60902
rect 4874 60891 5182 60900
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 4874 59868 5182 59877
rect 4874 59866 4880 59868
rect 4936 59866 4960 59868
rect 5016 59866 5040 59868
rect 5096 59866 5120 59868
rect 5176 59866 5182 59868
rect 4936 59814 4938 59866
rect 5118 59814 5120 59866
rect 4874 59812 4880 59814
rect 4936 59812 4960 59814
rect 5016 59812 5040 59814
rect 5096 59812 5120 59814
rect 5176 59812 5182 59814
rect 4874 59803 5182 59812
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4874 58780 5182 58789
rect 4874 58778 4880 58780
rect 4936 58778 4960 58780
rect 5016 58778 5040 58780
rect 5096 58778 5120 58780
rect 5176 58778 5182 58780
rect 4936 58726 4938 58778
rect 5118 58726 5120 58778
rect 4874 58724 4880 58726
rect 4936 58724 4960 58726
rect 5016 58724 5040 58726
rect 5096 58724 5120 58726
rect 5176 58724 5182 58726
rect 4874 58715 5182 58724
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4874 57692 5182 57701
rect 4874 57690 4880 57692
rect 4936 57690 4960 57692
rect 5016 57690 5040 57692
rect 5096 57690 5120 57692
rect 5176 57690 5182 57692
rect 4936 57638 4938 57690
rect 5118 57638 5120 57690
rect 4874 57636 4880 57638
rect 4936 57636 4960 57638
rect 5016 57636 5040 57638
rect 5096 57636 5120 57638
rect 5176 57636 5182 57638
rect 4874 57627 5182 57636
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4874 56604 5182 56613
rect 4874 56602 4880 56604
rect 4936 56602 4960 56604
rect 5016 56602 5040 56604
rect 5096 56602 5120 56604
rect 5176 56602 5182 56604
rect 4936 56550 4938 56602
rect 5118 56550 5120 56602
rect 4874 56548 4880 56550
rect 4936 56548 4960 56550
rect 5016 56548 5040 56550
rect 5096 56548 5120 56550
rect 5176 56548 5182 56550
rect 4874 56539 5182 56548
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4874 55516 5182 55525
rect 4874 55514 4880 55516
rect 4936 55514 4960 55516
rect 5016 55514 5040 55516
rect 5096 55514 5120 55516
rect 5176 55514 5182 55516
rect 4936 55462 4938 55514
rect 5118 55462 5120 55514
rect 4874 55460 4880 55462
rect 4936 55460 4960 55462
rect 5016 55460 5040 55462
rect 5096 55460 5120 55462
rect 5176 55460 5182 55462
rect 4874 55451 5182 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4874 54428 5182 54437
rect 4874 54426 4880 54428
rect 4936 54426 4960 54428
rect 5016 54426 5040 54428
rect 5096 54426 5120 54428
rect 5176 54426 5182 54428
rect 4936 54374 4938 54426
rect 5118 54374 5120 54426
rect 4874 54372 4880 54374
rect 4936 54372 4960 54374
rect 5016 54372 5040 54374
rect 5096 54372 5120 54374
rect 5176 54372 5182 54374
rect 4874 54363 5182 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4874 53340 5182 53349
rect 4874 53338 4880 53340
rect 4936 53338 4960 53340
rect 5016 53338 5040 53340
rect 5096 53338 5120 53340
rect 5176 53338 5182 53340
rect 4936 53286 4938 53338
rect 5118 53286 5120 53338
rect 4874 53284 4880 53286
rect 4936 53284 4960 53286
rect 5016 53284 5040 53286
rect 5096 53284 5120 53286
rect 5176 53284 5182 53286
rect 4874 53275 5182 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4874 52252 5182 52261
rect 4874 52250 4880 52252
rect 4936 52250 4960 52252
rect 5016 52250 5040 52252
rect 5096 52250 5120 52252
rect 5176 52250 5182 52252
rect 4936 52198 4938 52250
rect 5118 52198 5120 52250
rect 4874 52196 4880 52198
rect 4936 52196 4960 52198
rect 5016 52196 5040 52198
rect 5096 52196 5120 52198
rect 5176 52196 5182 52198
rect 4874 52187 5182 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4874 51164 5182 51173
rect 4874 51162 4880 51164
rect 4936 51162 4960 51164
rect 5016 51162 5040 51164
rect 5096 51162 5120 51164
rect 5176 51162 5182 51164
rect 4936 51110 4938 51162
rect 5118 51110 5120 51162
rect 4874 51108 4880 51110
rect 4936 51108 4960 51110
rect 5016 51108 5040 51110
rect 5096 51108 5120 51110
rect 5176 51108 5182 51110
rect 4874 51099 5182 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4874 50076 5182 50085
rect 4874 50074 4880 50076
rect 4936 50074 4960 50076
rect 5016 50074 5040 50076
rect 5096 50074 5120 50076
rect 5176 50074 5182 50076
rect 4936 50022 4938 50074
rect 5118 50022 5120 50074
rect 4874 50020 4880 50022
rect 4936 50020 4960 50022
rect 5016 50020 5040 50022
rect 5096 50020 5120 50022
rect 5176 50020 5182 50022
rect 4874 50011 5182 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4874 48988 5182 48997
rect 4874 48986 4880 48988
rect 4936 48986 4960 48988
rect 5016 48986 5040 48988
rect 5096 48986 5120 48988
rect 5176 48986 5182 48988
rect 4936 48934 4938 48986
rect 5118 48934 5120 48986
rect 4874 48932 4880 48934
rect 4936 48932 4960 48934
rect 5016 48932 5040 48934
rect 5096 48932 5120 48934
rect 5176 48932 5182 48934
rect 4874 48923 5182 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4874 47900 5182 47909
rect 4874 47898 4880 47900
rect 4936 47898 4960 47900
rect 5016 47898 5040 47900
rect 5096 47898 5120 47900
rect 5176 47898 5182 47900
rect 4936 47846 4938 47898
rect 5118 47846 5120 47898
rect 4874 47844 4880 47846
rect 4936 47844 4960 47846
rect 5016 47844 5040 47846
rect 5096 47844 5120 47846
rect 5176 47844 5182 47846
rect 4874 47835 5182 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4874 46812 5182 46821
rect 4874 46810 4880 46812
rect 4936 46810 4960 46812
rect 5016 46810 5040 46812
rect 5096 46810 5120 46812
rect 5176 46810 5182 46812
rect 4936 46758 4938 46810
rect 5118 46758 5120 46810
rect 4874 46756 4880 46758
rect 4936 46756 4960 46758
rect 5016 46756 5040 46758
rect 5096 46756 5120 46758
rect 5176 46756 5182 46758
rect 4874 46747 5182 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4874 45724 5182 45733
rect 4874 45722 4880 45724
rect 4936 45722 4960 45724
rect 5016 45722 5040 45724
rect 5096 45722 5120 45724
rect 5176 45722 5182 45724
rect 4936 45670 4938 45722
rect 5118 45670 5120 45722
rect 4874 45668 4880 45670
rect 4936 45668 4960 45670
rect 5016 45668 5040 45670
rect 5096 45668 5120 45670
rect 5176 45668 5182 45670
rect 4874 45659 5182 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4874 44636 5182 44645
rect 4874 44634 4880 44636
rect 4936 44634 4960 44636
rect 5016 44634 5040 44636
rect 5096 44634 5120 44636
rect 5176 44634 5182 44636
rect 4936 44582 4938 44634
rect 5118 44582 5120 44634
rect 4874 44580 4880 44582
rect 4936 44580 4960 44582
rect 5016 44580 5040 44582
rect 5096 44580 5120 44582
rect 5176 44580 5182 44582
rect 4874 44571 5182 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 7564 41472 7616 41478
rect 7564 41414 7616 41420
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 7576 41313 7604 41414
rect 7562 41304 7618 41313
rect 7562 41239 7618 41248
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 7564 39840 7616 39846
rect 7564 39782 7616 39788
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 7576 39545 7604 39782
rect 7562 39536 7618 39545
rect 7562 39471 7618 39480
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 7564 38752 7616 38758
rect 7564 38694 7616 38700
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 7576 38321 7604 38694
rect 7562 38312 7618 38321
rect 7562 38247 7618 38256
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 7562 36816 7618 36825
rect 7562 36751 7564 36760
rect 7616 36751 7618 36760
rect 7564 36722 7616 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 7562 35592 7618 35601
rect 7562 35527 7564 35536
rect 7616 35527 7618 35536
rect 7564 35498 7616 35504
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 7562 34096 7618 34105
rect 7562 34031 7564 34040
rect 7616 34031 7618 34040
rect 7564 34002 7616 34008
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 7562 15600 7618 15609
rect 7562 15535 7564 15544
rect 7616 15535 7618 15544
rect 7564 15506 7616 15512
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 8220 9654 8248 67118
rect 43168 67040 43220 67046
rect 43168 66982 43220 66988
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 35594 66396 35902 66405
rect 35594 66394 35600 66396
rect 35656 66394 35680 66396
rect 35736 66394 35760 66396
rect 35816 66394 35840 66396
rect 35896 66394 35902 66396
rect 35656 66342 35658 66394
rect 35838 66342 35840 66394
rect 35594 66340 35600 66342
rect 35656 66340 35680 66342
rect 35736 66340 35760 66342
rect 35816 66340 35840 66342
rect 35896 66340 35902 66342
rect 35594 66331 35902 66340
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 43180 64161 43208 66982
rect 44744 66774 44772 67186
rect 45112 67182 45140 71538
rect 46940 67244 46992 67250
rect 46940 67186 46992 67192
rect 45100 67176 45152 67182
rect 45100 67118 45152 67124
rect 45376 67040 45428 67046
rect 45376 66982 45428 66988
rect 44732 66768 44784 66774
rect 44732 66710 44784 66716
rect 43166 64152 43222 64161
rect 43166 64087 43222 64096
rect 45388 63889 45416 66982
rect 46952 66706 46980 67186
rect 47320 67182 47348 71538
rect 49528 67386 49556 71538
rect 51644 67386 51672 71538
rect 49516 67380 49568 67386
rect 49516 67322 49568 67328
rect 51632 67380 51684 67386
rect 51632 67322 51684 67328
rect 47676 67244 47728 67250
rect 47676 67186 47728 67192
rect 49148 67244 49200 67250
rect 49148 67186 49200 67192
rect 47308 67176 47360 67182
rect 47308 67118 47360 67124
rect 47584 67040 47636 67046
rect 47584 66982 47636 66988
rect 46940 66700 46992 66706
rect 46940 66642 46992 66648
rect 47596 64025 47624 66982
rect 47688 66842 47716 67186
rect 47676 66836 47728 66842
rect 47676 66778 47728 66784
rect 48688 66768 48740 66774
rect 48688 66710 48740 66716
rect 48700 66230 48728 66710
rect 49160 66298 49188 67186
rect 49700 67176 49752 67182
rect 49700 67118 49752 67124
rect 49976 67176 50028 67182
rect 49976 67118 50028 67124
rect 53472 67176 53524 67182
rect 53472 67118 53524 67124
rect 49712 67046 49740 67118
rect 49700 67040 49752 67046
rect 49700 66982 49752 66988
rect 49712 66842 49740 66982
rect 49700 66836 49752 66842
rect 49700 66778 49752 66784
rect 49700 66564 49752 66570
rect 49700 66506 49752 66512
rect 49712 66337 49740 66506
rect 49698 66328 49754 66337
rect 49148 66292 49200 66298
rect 49698 66263 49754 66272
rect 49148 66234 49200 66240
rect 48688 66224 48740 66230
rect 48688 66166 48740 66172
rect 49988 64161 50016 67118
rect 51632 67040 51684 67046
rect 51632 66982 51684 66988
rect 51644 66706 51672 66982
rect 53484 66706 53512 67118
rect 53576 66842 53604 71538
rect 55508 67386 55536 71538
rect 57440 67386 57468 71538
rect 59648 67386 59676 71538
rect 61580 67386 61608 71538
rect 55496 67380 55548 67386
rect 55496 67322 55548 67328
rect 57428 67380 57480 67386
rect 57428 67322 57480 67328
rect 59636 67380 59688 67386
rect 59636 67322 59688 67328
rect 60832 67380 60884 67386
rect 60832 67322 60884 67328
rect 61568 67380 61620 67386
rect 61568 67322 61620 67328
rect 53932 67312 53984 67318
rect 53932 67254 53984 67260
rect 57796 67312 57848 67318
rect 57796 67254 57848 67260
rect 53656 67040 53708 67046
rect 53656 66982 53708 66988
rect 53564 66836 53616 66842
rect 53564 66778 53616 66784
rect 50528 66700 50580 66706
rect 50528 66642 50580 66648
rect 51632 66700 51684 66706
rect 51632 66642 51684 66648
rect 53472 66700 53524 66706
rect 53472 66642 53524 66648
rect 50540 66230 50568 66642
rect 53668 66473 53696 66982
rect 53654 66464 53710 66473
rect 53654 66399 53710 66408
rect 53944 66230 53972 67254
rect 54944 67244 54996 67250
rect 54944 67186 54996 67192
rect 54956 66842 54984 67186
rect 55404 67176 55456 67182
rect 55404 67118 55456 67124
rect 55680 67176 55732 67182
rect 55680 67118 55732 67124
rect 54944 66836 54996 66842
rect 54944 66778 54996 66784
rect 55416 66638 55444 67118
rect 55692 66745 55720 67118
rect 55678 66736 55734 66745
rect 55678 66671 55734 66680
rect 55404 66632 55456 66638
rect 55404 66574 55456 66580
rect 55312 66564 55364 66570
rect 55312 66506 55364 66512
rect 55324 66230 55352 66506
rect 56600 66496 56652 66502
rect 56600 66438 56652 66444
rect 56612 66298 56640 66438
rect 56600 66292 56652 66298
rect 56600 66234 56652 66240
rect 50528 66224 50580 66230
rect 50528 66166 50580 66172
rect 53932 66224 53984 66230
rect 53932 66166 53984 66172
rect 55312 66224 55364 66230
rect 55312 66166 55364 66172
rect 57808 65958 57836 67254
rect 57888 67176 57940 67182
rect 57888 67118 57940 67124
rect 58164 67176 58216 67182
rect 58164 67118 58216 67124
rect 59728 67176 59780 67182
rect 59728 67118 59780 67124
rect 60004 67176 60056 67182
rect 60004 67118 60056 67124
rect 57900 66298 57928 67118
rect 57980 66836 58032 66842
rect 57980 66778 58032 66784
rect 57888 66292 57940 66298
rect 57888 66234 57940 66240
rect 57992 66162 58020 66778
rect 57980 66156 58032 66162
rect 57980 66098 58032 66104
rect 57796 65952 57848 65958
rect 57796 65894 57848 65900
rect 49974 64152 50030 64161
rect 49974 64087 50030 64096
rect 47582 64016 47638 64025
rect 47582 63951 47638 63960
rect 58176 63889 58204 67118
rect 59740 66842 59768 67118
rect 59728 66836 59780 66842
rect 59728 66778 59780 66784
rect 59740 66298 59768 66778
rect 60016 66473 60044 67118
rect 60002 66464 60058 66473
rect 60002 66399 60058 66408
rect 59728 66292 59780 66298
rect 59728 66234 59780 66240
rect 60844 66230 60872 67322
rect 62028 67312 62080 67318
rect 62028 67254 62080 67260
rect 61292 67040 61344 67046
rect 61292 66982 61344 66988
rect 61304 66842 61332 66982
rect 61292 66836 61344 66842
rect 61292 66778 61344 66784
rect 61660 66564 61712 66570
rect 61660 66506 61712 66512
rect 61672 66337 61700 66506
rect 61658 66328 61714 66337
rect 61658 66263 61714 66272
rect 60832 66224 60884 66230
rect 60832 66166 60884 66172
rect 62040 65958 62068 67254
rect 63144 66774 63172 71538
rect 65444 67386 65472 71538
rect 65654 71292 65962 71301
rect 65654 71290 65660 71292
rect 65716 71290 65740 71292
rect 65796 71290 65820 71292
rect 65876 71290 65900 71292
rect 65956 71290 65962 71292
rect 65716 71238 65718 71290
rect 65898 71238 65900 71290
rect 65654 71236 65660 71238
rect 65716 71236 65740 71238
rect 65796 71236 65820 71238
rect 65876 71236 65900 71238
rect 65956 71236 65962 71238
rect 65654 71227 65962 71236
rect 66314 70748 66622 70757
rect 66314 70746 66320 70748
rect 66376 70746 66400 70748
rect 66456 70746 66480 70748
rect 66536 70746 66560 70748
rect 66616 70746 66622 70748
rect 66376 70694 66378 70746
rect 66558 70694 66560 70746
rect 66314 70692 66320 70694
rect 66376 70692 66400 70694
rect 66456 70692 66480 70694
rect 66536 70692 66560 70694
rect 66616 70692 66622 70694
rect 66314 70683 66622 70692
rect 65654 70204 65962 70213
rect 65654 70202 65660 70204
rect 65716 70202 65740 70204
rect 65796 70202 65820 70204
rect 65876 70202 65900 70204
rect 65956 70202 65962 70204
rect 65716 70150 65718 70202
rect 65898 70150 65900 70202
rect 65654 70148 65660 70150
rect 65716 70148 65740 70150
rect 65796 70148 65820 70150
rect 65876 70148 65900 70150
rect 65956 70148 65962 70150
rect 65654 70139 65962 70148
rect 66314 69660 66622 69669
rect 66314 69658 66320 69660
rect 66376 69658 66400 69660
rect 66456 69658 66480 69660
rect 66536 69658 66560 69660
rect 66616 69658 66622 69660
rect 66376 69606 66378 69658
rect 66558 69606 66560 69658
rect 66314 69604 66320 69606
rect 66376 69604 66400 69606
rect 66456 69604 66480 69606
rect 66536 69604 66560 69606
rect 66616 69604 66622 69606
rect 66314 69595 66622 69604
rect 65654 69116 65962 69125
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69051 65962 69060
rect 66314 68572 66622 68581
rect 66314 68570 66320 68572
rect 66376 68570 66400 68572
rect 66456 68570 66480 68572
rect 66536 68570 66560 68572
rect 66616 68570 66622 68572
rect 66376 68518 66378 68570
rect 66558 68518 66560 68570
rect 66314 68516 66320 68518
rect 66376 68516 66400 68518
rect 66456 68516 66480 68518
rect 66536 68516 66560 68518
rect 66616 68516 66622 68518
rect 66314 68507 66622 68516
rect 65654 68028 65962 68037
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67963 65962 67972
rect 66314 67484 66622 67493
rect 66314 67482 66320 67484
rect 66376 67482 66400 67484
rect 66456 67482 66480 67484
rect 66536 67482 66560 67484
rect 66616 67482 66622 67484
rect 66376 67430 66378 67482
rect 66558 67430 66560 67482
rect 66314 67428 66320 67430
rect 66376 67428 66400 67430
rect 66456 67428 66480 67430
rect 66536 67428 66560 67430
rect 66616 67428 66622 67430
rect 66314 67419 66622 67428
rect 67376 67386 67404 71538
rect 69952 67386 69980 71538
rect 71884 67386 71912 71538
rect 65432 67380 65484 67386
rect 65432 67322 65484 67328
rect 67364 67380 67416 67386
rect 67364 67322 67416 67328
rect 68744 67380 68796 67386
rect 68744 67322 68796 67328
rect 69940 67380 69992 67386
rect 69940 67322 69992 67328
rect 71872 67380 71924 67386
rect 71872 67322 71924 67328
rect 66168 67312 66220 67318
rect 66168 67254 66220 67260
rect 67548 67312 67600 67318
rect 67548 67254 67600 67260
rect 65524 67244 65576 67250
rect 65524 67186 65576 67192
rect 63960 67176 64012 67182
rect 63960 67118 64012 67124
rect 64696 67176 64748 67182
rect 64696 67118 64748 67124
rect 63132 66768 63184 66774
rect 63132 66710 63184 66716
rect 63972 66473 64000 67118
rect 63958 66464 64014 66473
rect 63958 66399 64014 66408
rect 64604 66156 64656 66162
rect 64604 66098 64656 66104
rect 64616 65958 64644 66098
rect 62028 65952 62080 65958
rect 62028 65894 62080 65900
rect 63408 65952 63460 65958
rect 63408 65894 63460 65900
rect 64604 65952 64656 65958
rect 64604 65894 64656 65900
rect 63420 65754 63448 65894
rect 63408 65748 63460 65754
rect 63408 65690 63460 65696
rect 64708 65521 64736 67118
rect 65536 67046 65564 67186
rect 65524 67040 65576 67046
rect 65524 66982 65576 66988
rect 65536 66842 65564 66982
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 65524 66836 65576 66842
rect 65524 66778 65576 66784
rect 64880 66564 64932 66570
rect 64880 66506 64932 66512
rect 64892 66230 64920 66506
rect 66180 66230 66208 67254
rect 66314 66396 66622 66405
rect 66314 66394 66320 66396
rect 66376 66394 66400 66396
rect 66456 66394 66480 66396
rect 66536 66394 66560 66396
rect 66616 66394 66622 66396
rect 66376 66342 66378 66394
rect 66558 66342 66560 66394
rect 66314 66340 66320 66342
rect 66376 66340 66400 66342
rect 66456 66340 66480 66342
rect 66536 66340 66560 66342
rect 66616 66340 66622 66342
rect 66314 66331 66622 66340
rect 67560 66230 67588 67254
rect 68468 67176 68520 67182
rect 68468 67118 68520 67124
rect 68008 67040 68060 67046
rect 68008 66982 68060 66988
rect 68020 66842 68048 66982
rect 68008 66836 68060 66842
rect 68008 66778 68060 66784
rect 68480 66609 68508 67118
rect 68466 66600 68522 66609
rect 68466 66535 68522 66544
rect 64880 66224 64932 66230
rect 64880 66166 64932 66172
rect 66168 66224 66220 66230
rect 66168 66166 66220 66172
rect 67548 66224 67600 66230
rect 67548 66166 67600 66172
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 64694 65512 64750 65521
rect 64694 65447 64750 65456
rect 68756 65385 68784 67322
rect 74080 67312 74132 67318
rect 74080 67254 74132 67260
rect 69572 67244 69624 67250
rect 69572 67186 69624 67192
rect 71412 67244 71464 67250
rect 71412 67186 71464 67192
rect 69584 66230 69612 67186
rect 69940 67176 69992 67182
rect 69940 67118 69992 67124
rect 69952 67046 69980 67118
rect 69940 67040 69992 67046
rect 69940 66982 69992 66988
rect 69952 66842 69980 66982
rect 69940 66836 69992 66842
rect 69940 66778 69992 66784
rect 71228 66564 71280 66570
rect 71228 66506 71280 66512
rect 69572 66224 69624 66230
rect 69572 66166 69624 66172
rect 68742 65376 68798 65385
rect 68742 65311 68798 65320
rect 71240 65113 71268 66506
rect 71424 66230 71452 67186
rect 73712 67040 73764 67046
rect 73712 66982 73764 66988
rect 73724 66842 73752 66982
rect 73712 66836 73764 66842
rect 73712 66778 73764 66784
rect 73436 66564 73488 66570
rect 73436 66506 73488 66512
rect 73448 66230 73476 66506
rect 71412 66224 71464 66230
rect 71412 66166 71464 66172
rect 73436 66224 73488 66230
rect 73436 66166 73488 66172
rect 74092 65385 74120 67254
rect 74184 66502 74212 71538
rect 76116 67386 76144 71538
rect 96374 71292 96682 71301
rect 96374 71290 96380 71292
rect 96436 71290 96460 71292
rect 96516 71290 96540 71292
rect 96596 71290 96620 71292
rect 96676 71290 96682 71292
rect 96436 71238 96438 71290
rect 96618 71238 96620 71290
rect 96374 71236 96380 71238
rect 96436 71236 96460 71238
rect 96516 71236 96540 71238
rect 96596 71236 96620 71238
rect 96676 71236 96682 71238
rect 96374 71227 96682 71236
rect 97034 70748 97342 70757
rect 97034 70746 97040 70748
rect 97096 70746 97120 70748
rect 97176 70746 97200 70748
rect 97256 70746 97280 70748
rect 97336 70746 97342 70748
rect 97096 70694 97098 70746
rect 97278 70694 97280 70746
rect 97034 70692 97040 70694
rect 97096 70692 97120 70694
rect 97176 70692 97200 70694
rect 97256 70692 97280 70694
rect 97336 70692 97342 70694
rect 97034 70683 97342 70692
rect 96374 70204 96682 70213
rect 96374 70202 96380 70204
rect 96436 70202 96460 70204
rect 96516 70202 96540 70204
rect 96596 70202 96620 70204
rect 96676 70202 96682 70204
rect 96436 70150 96438 70202
rect 96618 70150 96620 70202
rect 96374 70148 96380 70150
rect 96436 70148 96460 70150
rect 96516 70148 96540 70150
rect 96596 70148 96620 70150
rect 96676 70148 96682 70150
rect 96374 70139 96682 70148
rect 97034 69660 97342 69669
rect 97034 69658 97040 69660
rect 97096 69658 97120 69660
rect 97176 69658 97200 69660
rect 97256 69658 97280 69660
rect 97336 69658 97342 69660
rect 97096 69606 97098 69658
rect 97278 69606 97280 69658
rect 97034 69604 97040 69606
rect 97096 69604 97120 69606
rect 97176 69604 97200 69606
rect 97256 69604 97280 69606
rect 97336 69604 97342 69606
rect 97034 69595 97342 69604
rect 96374 69116 96682 69125
rect 96374 69114 96380 69116
rect 96436 69114 96460 69116
rect 96516 69114 96540 69116
rect 96596 69114 96620 69116
rect 96676 69114 96682 69116
rect 96436 69062 96438 69114
rect 96618 69062 96620 69114
rect 96374 69060 96380 69062
rect 96436 69060 96460 69062
rect 96516 69060 96540 69062
rect 96596 69060 96620 69062
rect 96676 69060 96682 69062
rect 96374 69051 96682 69060
rect 97034 68572 97342 68581
rect 97034 68570 97040 68572
rect 97096 68570 97120 68572
rect 97176 68570 97200 68572
rect 97256 68570 97280 68572
rect 97336 68570 97342 68572
rect 97096 68518 97098 68570
rect 97278 68518 97280 68570
rect 97034 68516 97040 68518
rect 97096 68516 97120 68518
rect 97176 68516 97200 68518
rect 97256 68516 97280 68518
rect 97336 68516 97342 68518
rect 97034 68507 97342 68516
rect 96374 68028 96682 68037
rect 96374 68026 96380 68028
rect 96436 68026 96460 68028
rect 96516 68026 96540 68028
rect 96596 68026 96620 68028
rect 96676 68026 96682 68028
rect 96436 67974 96438 68026
rect 96618 67974 96620 68026
rect 96374 67972 96380 67974
rect 96436 67972 96460 67974
rect 96516 67972 96540 67974
rect 96596 67972 96620 67974
rect 96676 67972 96682 67974
rect 96374 67963 96682 67972
rect 97034 67484 97342 67493
rect 97034 67482 97040 67484
rect 97096 67482 97120 67484
rect 97176 67482 97200 67484
rect 97256 67482 97280 67484
rect 97336 67482 97342 67484
rect 97096 67430 97098 67482
rect 97278 67430 97280 67482
rect 97034 67428 97040 67430
rect 97096 67428 97120 67430
rect 97176 67428 97200 67430
rect 97256 67428 97280 67430
rect 97336 67428 97342 67430
rect 97034 67419 97342 67428
rect 76104 67380 76156 67386
rect 76104 67322 76156 67328
rect 75736 67244 75788 67250
rect 75736 67186 75788 67192
rect 74172 66496 74224 66502
rect 74172 66438 74224 66444
rect 75748 66298 75776 67186
rect 95884 67040 95936 67046
rect 95884 66982 95936 66988
rect 75736 66292 75788 66298
rect 75736 66234 75788 66240
rect 95896 66230 95924 66982
rect 96374 66940 96682 66949
rect 96374 66938 96380 66940
rect 96436 66938 96460 66940
rect 96516 66938 96540 66940
rect 96596 66938 96620 66940
rect 96676 66938 96682 66940
rect 96436 66886 96438 66938
rect 96618 66886 96620 66938
rect 96374 66884 96380 66886
rect 96436 66884 96460 66886
rect 96516 66884 96540 66886
rect 96596 66884 96620 66886
rect 96676 66884 96682 66886
rect 96374 66875 96682 66884
rect 97034 66396 97342 66405
rect 97034 66394 97040 66396
rect 97096 66394 97120 66396
rect 97176 66394 97200 66396
rect 97256 66394 97280 66396
rect 97336 66394 97342 66396
rect 97096 66342 97098 66394
rect 97278 66342 97280 66394
rect 97034 66340 97040 66342
rect 97096 66340 97120 66342
rect 97176 66340 97200 66342
rect 97256 66340 97280 66342
rect 97336 66340 97342 66342
rect 97034 66331 97342 66340
rect 107762 66396 108070 66405
rect 107762 66394 107768 66396
rect 107824 66394 107848 66396
rect 107904 66394 107928 66396
rect 107984 66394 108008 66396
rect 108064 66394 108070 66396
rect 107824 66342 107826 66394
rect 108006 66342 108008 66394
rect 107762 66340 107768 66342
rect 107824 66340 107848 66342
rect 107904 66340 107928 66342
rect 107984 66340 108008 66342
rect 108064 66340 108070 66342
rect 107762 66331 108070 66340
rect 95884 66224 95936 66230
rect 95884 66166 95936 66172
rect 75736 66156 75788 66162
rect 75736 66098 75788 66104
rect 92388 66156 92440 66162
rect 92388 66098 92440 66104
rect 75748 65958 75776 66098
rect 76472 66088 76524 66094
rect 76472 66030 76524 66036
rect 75736 65952 75788 65958
rect 75736 65894 75788 65900
rect 76288 65952 76340 65958
rect 76484 65940 76512 66030
rect 76340 65912 76512 65940
rect 86316 65952 86368 65958
rect 76288 65894 76340 65900
rect 86316 65894 86368 65900
rect 87328 65952 87380 65958
rect 87328 65894 87380 65900
rect 92296 65952 92348 65958
rect 92296 65894 92348 65900
rect 74078 65376 74134 65385
rect 74078 65311 74134 65320
rect 71226 65104 71282 65113
rect 71226 65039 71282 65048
rect 86328 64025 86356 65894
rect 87340 65385 87368 65894
rect 92308 65686 92336 65894
rect 92296 65680 92348 65686
rect 92296 65622 92348 65628
rect 87326 65376 87382 65385
rect 87326 65311 87382 65320
rect 92400 64938 92428 66098
rect 92388 64932 92440 64938
rect 92388 64874 92440 64880
rect 86314 64016 86370 64025
rect 86314 63951 86370 63960
rect 95896 63889 95924 66166
rect 102784 66020 102836 66026
rect 102784 65962 102836 65968
rect 96374 65852 96682 65861
rect 96374 65850 96380 65852
rect 96436 65850 96460 65852
rect 96516 65850 96540 65852
rect 96596 65850 96620 65852
rect 96676 65850 96682 65852
rect 96436 65798 96438 65850
rect 96618 65798 96620 65850
rect 96374 65796 96380 65798
rect 96436 65796 96460 65798
rect 96516 65796 96540 65798
rect 96596 65796 96620 65798
rect 96676 65796 96682 65798
rect 96374 65787 96682 65796
rect 100760 65748 100812 65754
rect 100760 65690 100812 65696
rect 100772 64326 100800 65690
rect 100760 64320 100812 64326
rect 100760 64262 100812 64268
rect 45374 63880 45430 63889
rect 45374 63815 45430 63824
rect 58162 63880 58218 63889
rect 58162 63815 58218 63824
rect 95882 63880 95938 63889
rect 95882 63815 95938 63824
rect 102796 11762 102824 65962
rect 107026 65852 107334 65861
rect 107026 65850 107032 65852
rect 107088 65850 107112 65852
rect 107168 65850 107192 65852
rect 107248 65850 107272 65852
rect 107328 65850 107334 65852
rect 107088 65798 107090 65850
rect 107270 65798 107272 65850
rect 107026 65796 107032 65798
rect 107088 65796 107112 65798
rect 107168 65796 107192 65798
rect 107248 65796 107272 65798
rect 107328 65796 107334 65798
rect 107026 65787 107334 65796
rect 102968 65680 103020 65686
rect 102968 65622 103020 65628
rect 102876 64932 102928 64938
rect 102876 64874 102928 64880
rect 102888 54194 102916 64874
rect 102980 57934 103008 65622
rect 107762 65308 108070 65317
rect 107762 65306 107768 65308
rect 107824 65306 107848 65308
rect 107904 65306 107928 65308
rect 107984 65306 108008 65308
rect 108064 65306 108070 65308
rect 107824 65254 107826 65306
rect 108006 65254 108008 65306
rect 107762 65252 107768 65254
rect 107824 65252 107848 65254
rect 107904 65252 107928 65254
rect 107984 65252 108008 65254
rect 108064 65252 108070 65254
rect 107762 65243 108070 65252
rect 107026 64764 107334 64773
rect 107026 64762 107032 64764
rect 107088 64762 107112 64764
rect 107168 64762 107192 64764
rect 107248 64762 107272 64764
rect 107328 64762 107334 64764
rect 107088 64710 107090 64762
rect 107270 64710 107272 64762
rect 107026 64708 107032 64710
rect 107088 64708 107112 64710
rect 107168 64708 107192 64710
rect 107248 64708 107272 64710
rect 107328 64708 107334 64710
rect 107026 64699 107334 64708
rect 104440 64320 104492 64326
rect 104440 64262 104492 64268
rect 104346 63880 104402 63889
rect 104346 63815 104402 63824
rect 103704 60104 103756 60110
rect 103704 60046 103756 60052
rect 103716 59809 103744 60046
rect 103702 59800 103758 59809
rect 103702 59735 103758 59744
rect 102968 57928 103020 57934
rect 102968 57870 103020 57876
rect 104360 57458 104388 63815
rect 104348 57452 104400 57458
rect 104348 57394 104400 57400
rect 104360 57338 104388 57394
rect 104268 57310 104388 57338
rect 104268 54738 104296 57310
rect 104256 54732 104308 54738
rect 104256 54674 104308 54680
rect 102876 54188 102928 54194
rect 102876 54130 102928 54136
rect 104256 46096 104308 46102
rect 104256 46038 104308 46044
rect 104164 42560 104216 42566
rect 104164 42502 104216 42508
rect 104176 25129 104204 42502
rect 104268 41138 104296 46038
rect 104452 45554 104480 64262
rect 107762 64220 108070 64229
rect 107762 64218 107768 64220
rect 107824 64218 107848 64220
rect 107904 64218 107928 64220
rect 107984 64218 108008 64220
rect 108064 64218 108070 64220
rect 107824 64166 107826 64218
rect 108006 64166 108008 64218
rect 107762 64164 107768 64166
rect 107824 64164 107848 64166
rect 107904 64164 107928 64166
rect 107984 64164 108008 64166
rect 108064 64164 108070 64166
rect 104990 64152 105046 64161
rect 107762 64155 108070 64164
rect 104990 64087 105046 64096
rect 105004 57390 105032 64087
rect 106186 64016 106242 64025
rect 106186 63951 106242 63960
rect 104624 57384 104676 57390
rect 104624 57326 104676 57332
rect 104992 57384 105044 57390
rect 104992 57326 105044 57332
rect 104532 56704 104584 56710
rect 104532 56646 104584 56652
rect 104544 55758 104572 56646
rect 104636 55962 104664 57326
rect 105004 56914 105032 57326
rect 104992 56908 105044 56914
rect 104992 56850 105044 56856
rect 104624 55956 104676 55962
rect 104624 55898 104676 55904
rect 104532 55752 104584 55758
rect 104532 55694 104584 55700
rect 104624 54596 104676 54602
rect 104624 54538 104676 54544
rect 104532 54188 104584 54194
rect 104532 54130 104584 54136
rect 104544 53990 104572 54130
rect 104532 53984 104584 53990
rect 104532 53926 104584 53932
rect 104360 45526 104480 45554
rect 104360 41614 104388 45526
rect 104544 43994 104572 53926
rect 104636 53786 104664 54538
rect 105004 53786 105032 56850
rect 106200 54602 106228 63951
rect 107026 63676 107334 63685
rect 107026 63674 107032 63676
rect 107088 63674 107112 63676
rect 107168 63674 107192 63676
rect 107248 63674 107272 63676
rect 107328 63674 107334 63676
rect 107088 63622 107090 63674
rect 107270 63622 107272 63674
rect 107026 63620 107032 63622
rect 107088 63620 107112 63622
rect 107168 63620 107192 63622
rect 107248 63620 107272 63622
rect 107328 63620 107334 63622
rect 107026 63611 107334 63620
rect 107762 63132 108070 63141
rect 107762 63130 107768 63132
rect 107824 63130 107848 63132
rect 107904 63130 107928 63132
rect 107984 63130 108008 63132
rect 108064 63130 108070 63132
rect 107824 63078 107826 63130
rect 108006 63078 108008 63130
rect 107762 63076 107768 63078
rect 107824 63076 107848 63078
rect 107904 63076 107928 63078
rect 107984 63076 108008 63078
rect 108064 63076 108070 63078
rect 107762 63067 108070 63076
rect 107026 62588 107334 62597
rect 107026 62586 107032 62588
rect 107088 62586 107112 62588
rect 107168 62586 107192 62588
rect 107248 62586 107272 62588
rect 107328 62586 107334 62588
rect 107088 62534 107090 62586
rect 107270 62534 107272 62586
rect 107026 62532 107032 62534
rect 107088 62532 107112 62534
rect 107168 62532 107192 62534
rect 107248 62532 107272 62534
rect 107328 62532 107334 62534
rect 107026 62523 107334 62532
rect 107762 62044 108070 62053
rect 107762 62042 107768 62044
rect 107824 62042 107848 62044
rect 107904 62042 107928 62044
rect 107984 62042 108008 62044
rect 108064 62042 108070 62044
rect 107824 61990 107826 62042
rect 108006 61990 108008 62042
rect 107762 61988 107768 61990
rect 107824 61988 107848 61990
rect 107904 61988 107928 61990
rect 107984 61988 108008 61990
rect 108064 61988 108070 61990
rect 107762 61979 108070 61988
rect 107026 61500 107334 61509
rect 107026 61498 107032 61500
rect 107088 61498 107112 61500
rect 107168 61498 107192 61500
rect 107248 61498 107272 61500
rect 107328 61498 107334 61500
rect 107088 61446 107090 61498
rect 107270 61446 107272 61498
rect 107026 61444 107032 61446
rect 107088 61444 107112 61446
rect 107168 61444 107192 61446
rect 107248 61444 107272 61446
rect 107328 61444 107334 61446
rect 107026 61435 107334 61444
rect 107762 60956 108070 60965
rect 107762 60954 107768 60956
rect 107824 60954 107848 60956
rect 107904 60954 107928 60956
rect 107984 60954 108008 60956
rect 108064 60954 108070 60956
rect 107824 60902 107826 60954
rect 108006 60902 108008 60954
rect 107762 60900 107768 60902
rect 107824 60900 107848 60902
rect 107904 60900 107928 60902
rect 107984 60900 108008 60902
rect 108064 60900 108070 60902
rect 107762 60891 108070 60900
rect 107026 60412 107334 60421
rect 107026 60410 107032 60412
rect 107088 60410 107112 60412
rect 107168 60410 107192 60412
rect 107248 60410 107272 60412
rect 107328 60410 107334 60412
rect 107088 60358 107090 60410
rect 107270 60358 107272 60410
rect 107026 60356 107032 60358
rect 107088 60356 107112 60358
rect 107168 60356 107192 60358
rect 107248 60356 107272 60358
rect 107328 60356 107334 60358
rect 107026 60347 107334 60356
rect 107762 59868 108070 59877
rect 107762 59866 107768 59868
rect 107824 59866 107848 59868
rect 107904 59866 107928 59868
rect 107984 59866 108008 59868
rect 108064 59866 108070 59868
rect 107824 59814 107826 59866
rect 108006 59814 108008 59866
rect 107762 59812 107768 59814
rect 107824 59812 107848 59814
rect 107904 59812 107928 59814
rect 107984 59812 108008 59814
rect 108064 59812 108070 59814
rect 107762 59803 108070 59812
rect 107026 59324 107334 59333
rect 107026 59322 107032 59324
rect 107088 59322 107112 59324
rect 107168 59322 107192 59324
rect 107248 59322 107272 59324
rect 107328 59322 107334 59324
rect 107088 59270 107090 59322
rect 107270 59270 107272 59322
rect 107026 59268 107032 59270
rect 107088 59268 107112 59270
rect 107168 59268 107192 59270
rect 107248 59268 107272 59270
rect 107328 59268 107334 59270
rect 107026 59259 107334 59268
rect 107762 58780 108070 58789
rect 107762 58778 107768 58780
rect 107824 58778 107848 58780
rect 107904 58778 107928 58780
rect 107984 58778 108008 58780
rect 108064 58778 108070 58780
rect 107824 58726 107826 58778
rect 108006 58726 108008 58778
rect 107762 58724 107768 58726
rect 107824 58724 107848 58726
rect 107904 58724 107928 58726
rect 107984 58724 108008 58726
rect 108064 58724 108070 58726
rect 107762 58715 108070 58724
rect 107026 58236 107334 58245
rect 107026 58234 107032 58236
rect 107088 58234 107112 58236
rect 107168 58234 107192 58236
rect 107248 58234 107272 58236
rect 107328 58234 107334 58236
rect 107088 58182 107090 58234
rect 107270 58182 107272 58234
rect 107026 58180 107032 58182
rect 107088 58180 107112 58182
rect 107168 58180 107192 58182
rect 107248 58180 107272 58182
rect 107328 58180 107334 58182
rect 107026 58171 107334 58180
rect 107762 57692 108070 57701
rect 107762 57690 107768 57692
rect 107824 57690 107848 57692
rect 107904 57690 107928 57692
rect 107984 57690 108008 57692
rect 108064 57690 108070 57692
rect 107824 57638 107826 57690
rect 108006 57638 108008 57690
rect 107762 57636 107768 57638
rect 107824 57636 107848 57638
rect 107904 57636 107928 57638
rect 107984 57636 108008 57638
rect 108064 57636 108070 57638
rect 107762 57627 108070 57636
rect 106648 57248 106700 57254
rect 106648 57190 106700 57196
rect 106660 55214 106688 57190
rect 107026 57148 107334 57157
rect 107026 57146 107032 57148
rect 107088 57146 107112 57148
rect 107168 57146 107192 57148
rect 107248 57146 107272 57148
rect 107328 57146 107334 57148
rect 107088 57094 107090 57146
rect 107270 57094 107272 57146
rect 107026 57092 107032 57094
rect 107088 57092 107112 57094
rect 107168 57092 107192 57094
rect 107248 57092 107272 57094
rect 107328 57092 107334 57094
rect 107026 57083 107334 57092
rect 107762 56604 108070 56613
rect 107762 56602 107768 56604
rect 107824 56602 107848 56604
rect 107904 56602 107928 56604
rect 107984 56602 108008 56604
rect 108064 56602 108070 56604
rect 107824 56550 107826 56602
rect 108006 56550 108008 56602
rect 107762 56548 107768 56550
rect 107824 56548 107848 56550
rect 107904 56548 107928 56550
rect 107984 56548 108008 56550
rect 108064 56548 108070 56550
rect 107762 56539 108070 56548
rect 107026 56060 107334 56069
rect 107026 56058 107032 56060
rect 107088 56058 107112 56060
rect 107168 56058 107192 56060
rect 107248 56058 107272 56060
rect 107328 56058 107334 56060
rect 107088 56006 107090 56058
rect 107270 56006 107272 56058
rect 107026 56004 107032 56006
rect 107088 56004 107112 56006
rect 107168 56004 107192 56006
rect 107248 56004 107272 56006
rect 107328 56004 107334 56006
rect 107026 55995 107334 56004
rect 107762 55516 108070 55525
rect 107762 55514 107768 55516
rect 107824 55514 107848 55516
rect 107904 55514 107928 55516
rect 107984 55514 108008 55516
rect 108064 55514 108070 55516
rect 107824 55462 107826 55514
rect 108006 55462 108008 55514
rect 107762 55460 107768 55462
rect 107824 55460 107848 55462
rect 107904 55460 107928 55462
rect 107984 55460 108008 55462
rect 108064 55460 108070 55462
rect 107762 55451 108070 55460
rect 106384 55186 106688 55214
rect 106384 54738 106412 55186
rect 107026 54972 107334 54981
rect 107026 54970 107032 54972
rect 107088 54970 107112 54972
rect 107168 54970 107192 54972
rect 107248 54970 107272 54972
rect 107328 54970 107334 54972
rect 107088 54918 107090 54970
rect 107270 54918 107272 54970
rect 107026 54916 107032 54918
rect 107088 54916 107112 54918
rect 107168 54916 107192 54918
rect 107248 54916 107272 54918
rect 107328 54916 107334 54918
rect 107026 54907 107334 54916
rect 106372 54732 106424 54738
rect 106372 54674 106424 54680
rect 105084 54596 105136 54602
rect 105084 54538 105136 54544
rect 106188 54596 106240 54602
rect 106188 54538 106240 54544
rect 105096 54330 105124 54538
rect 105084 54324 105136 54330
rect 105084 54266 105136 54272
rect 104624 53780 104676 53786
rect 104624 53722 104676 53728
rect 104992 53780 105044 53786
rect 104992 53722 105044 53728
rect 104900 53644 104952 53650
rect 104900 53586 104952 53592
rect 104808 53576 104860 53582
rect 104808 53518 104860 53524
rect 104820 46170 104848 53518
rect 104808 46164 104860 46170
rect 104808 46106 104860 46112
rect 104820 45554 104848 46106
rect 104912 45966 104940 53586
rect 105004 53582 105032 53722
rect 106200 53650 106228 54538
rect 106188 53644 106240 53650
rect 106188 53586 106240 53592
rect 104992 53576 105044 53582
rect 104992 53518 105044 53524
rect 104900 45960 104952 45966
rect 104900 45902 104952 45908
rect 104912 45830 104940 45902
rect 104900 45824 104952 45830
rect 104900 45766 104952 45772
rect 105452 45824 105504 45830
rect 105452 45766 105504 45772
rect 104728 45526 104848 45554
rect 104728 45014 104756 45526
rect 104912 45082 104940 45766
rect 104900 45076 104952 45082
rect 104900 45018 104952 45024
rect 104716 45008 104768 45014
rect 104716 44950 104768 44956
rect 105464 44946 105492 45766
rect 105452 44940 105504 44946
rect 105452 44882 105504 44888
rect 105464 44742 105492 44882
rect 105176 44736 105228 44742
rect 105176 44678 105228 44684
rect 105452 44736 105504 44742
rect 105452 44678 105504 44684
rect 104532 43988 104584 43994
rect 104532 43930 104584 43936
rect 104544 43790 104572 43930
rect 104532 43784 104584 43790
rect 104532 43726 104584 43732
rect 104348 41608 104400 41614
rect 104348 41550 104400 41556
rect 104256 41132 104308 41138
rect 104256 41074 104308 41080
rect 104544 36922 104572 43726
rect 105084 43716 105136 43722
rect 105084 43658 105136 43664
rect 104992 42764 105044 42770
rect 104992 42706 105044 42712
rect 104624 42628 104676 42634
rect 104624 42570 104676 42576
rect 104636 41274 104664 42570
rect 105004 42226 105032 42706
rect 105096 42634 105124 43658
rect 105084 42628 105136 42634
rect 105084 42570 105136 42576
rect 104992 42220 105044 42226
rect 104992 42162 105044 42168
rect 104900 41608 104952 41614
rect 104900 41550 104952 41556
rect 104912 41274 104940 41550
rect 104624 41268 104676 41274
rect 104624 41210 104676 41216
rect 104900 41268 104952 41274
rect 104900 41210 104952 41216
rect 105188 40934 105216 44678
rect 105464 42566 105492 44678
rect 106384 42566 106412 54674
rect 107762 54428 108070 54437
rect 107762 54426 107768 54428
rect 107824 54426 107848 54428
rect 107904 54426 107928 54428
rect 107984 54426 108008 54428
rect 108064 54426 108070 54428
rect 107824 54374 107826 54426
rect 108006 54374 108008 54426
rect 107762 54372 107768 54374
rect 107824 54372 107848 54374
rect 107904 54372 107928 54374
rect 107984 54372 108008 54374
rect 108064 54372 108070 54374
rect 107762 54363 108070 54372
rect 107026 53884 107334 53893
rect 107026 53882 107032 53884
rect 107088 53882 107112 53884
rect 107168 53882 107192 53884
rect 107248 53882 107272 53884
rect 107328 53882 107334 53884
rect 107088 53830 107090 53882
rect 107270 53830 107272 53882
rect 107026 53828 107032 53830
rect 107088 53828 107112 53830
rect 107168 53828 107192 53830
rect 107248 53828 107272 53830
rect 107328 53828 107334 53830
rect 107026 53819 107334 53828
rect 107762 53340 108070 53349
rect 107762 53338 107768 53340
rect 107824 53338 107848 53340
rect 107904 53338 107928 53340
rect 107984 53338 108008 53340
rect 108064 53338 108070 53340
rect 107824 53286 107826 53338
rect 108006 53286 108008 53338
rect 107762 53284 107768 53286
rect 107824 53284 107848 53286
rect 107904 53284 107928 53286
rect 107984 53284 108008 53286
rect 108064 53284 108070 53286
rect 107762 53275 108070 53284
rect 107026 52796 107334 52805
rect 107026 52794 107032 52796
rect 107088 52794 107112 52796
rect 107168 52794 107192 52796
rect 107248 52794 107272 52796
rect 107328 52794 107334 52796
rect 107088 52742 107090 52794
rect 107270 52742 107272 52794
rect 107026 52740 107032 52742
rect 107088 52740 107112 52742
rect 107168 52740 107192 52742
rect 107248 52740 107272 52742
rect 107328 52740 107334 52742
rect 107026 52731 107334 52740
rect 107762 52252 108070 52261
rect 107762 52250 107768 52252
rect 107824 52250 107848 52252
rect 107904 52250 107928 52252
rect 107984 52250 108008 52252
rect 108064 52250 108070 52252
rect 107824 52198 107826 52250
rect 108006 52198 108008 52250
rect 107762 52196 107768 52198
rect 107824 52196 107848 52198
rect 107904 52196 107928 52198
rect 107984 52196 108008 52198
rect 108064 52196 108070 52198
rect 107762 52187 108070 52196
rect 107026 51708 107334 51717
rect 107026 51706 107032 51708
rect 107088 51706 107112 51708
rect 107168 51706 107192 51708
rect 107248 51706 107272 51708
rect 107328 51706 107334 51708
rect 107088 51654 107090 51706
rect 107270 51654 107272 51706
rect 107026 51652 107032 51654
rect 107088 51652 107112 51654
rect 107168 51652 107192 51654
rect 107248 51652 107272 51654
rect 107328 51652 107334 51654
rect 107026 51643 107334 51652
rect 107762 51164 108070 51173
rect 107762 51162 107768 51164
rect 107824 51162 107848 51164
rect 107904 51162 107928 51164
rect 107984 51162 108008 51164
rect 108064 51162 108070 51164
rect 107824 51110 107826 51162
rect 108006 51110 108008 51162
rect 107762 51108 107768 51110
rect 107824 51108 107848 51110
rect 107904 51108 107928 51110
rect 107984 51108 108008 51110
rect 108064 51108 108070 51110
rect 107762 51099 108070 51108
rect 107026 50620 107334 50629
rect 107026 50618 107032 50620
rect 107088 50618 107112 50620
rect 107168 50618 107192 50620
rect 107248 50618 107272 50620
rect 107328 50618 107334 50620
rect 107088 50566 107090 50618
rect 107270 50566 107272 50618
rect 107026 50564 107032 50566
rect 107088 50564 107112 50566
rect 107168 50564 107192 50566
rect 107248 50564 107272 50566
rect 107328 50564 107334 50566
rect 107026 50555 107334 50564
rect 107762 50076 108070 50085
rect 107762 50074 107768 50076
rect 107824 50074 107848 50076
rect 107904 50074 107928 50076
rect 107984 50074 108008 50076
rect 108064 50074 108070 50076
rect 107824 50022 107826 50074
rect 108006 50022 108008 50074
rect 107762 50020 107768 50022
rect 107824 50020 107848 50022
rect 107904 50020 107928 50022
rect 107984 50020 108008 50022
rect 108064 50020 108070 50022
rect 107762 50011 108070 50020
rect 107026 49532 107334 49541
rect 107026 49530 107032 49532
rect 107088 49530 107112 49532
rect 107168 49530 107192 49532
rect 107248 49530 107272 49532
rect 107328 49530 107334 49532
rect 107088 49478 107090 49530
rect 107270 49478 107272 49530
rect 107026 49476 107032 49478
rect 107088 49476 107112 49478
rect 107168 49476 107192 49478
rect 107248 49476 107272 49478
rect 107328 49476 107334 49478
rect 107026 49467 107334 49476
rect 107762 48988 108070 48997
rect 107762 48986 107768 48988
rect 107824 48986 107848 48988
rect 107904 48986 107928 48988
rect 107984 48986 108008 48988
rect 108064 48986 108070 48988
rect 107824 48934 107826 48986
rect 108006 48934 108008 48986
rect 107762 48932 107768 48934
rect 107824 48932 107848 48934
rect 107904 48932 107928 48934
rect 107984 48932 108008 48934
rect 108064 48932 108070 48934
rect 107762 48923 108070 48932
rect 107026 48444 107334 48453
rect 107026 48442 107032 48444
rect 107088 48442 107112 48444
rect 107168 48442 107192 48444
rect 107248 48442 107272 48444
rect 107328 48442 107334 48444
rect 107088 48390 107090 48442
rect 107270 48390 107272 48442
rect 107026 48388 107032 48390
rect 107088 48388 107112 48390
rect 107168 48388 107192 48390
rect 107248 48388 107272 48390
rect 107328 48388 107334 48390
rect 107026 48379 107334 48388
rect 107762 47900 108070 47909
rect 107762 47898 107768 47900
rect 107824 47898 107848 47900
rect 107904 47898 107928 47900
rect 107984 47898 108008 47900
rect 108064 47898 108070 47900
rect 107824 47846 107826 47898
rect 108006 47846 108008 47898
rect 107762 47844 107768 47846
rect 107824 47844 107848 47846
rect 107904 47844 107928 47846
rect 107984 47844 108008 47846
rect 108064 47844 108070 47846
rect 107762 47835 108070 47844
rect 107026 47356 107334 47365
rect 107026 47354 107032 47356
rect 107088 47354 107112 47356
rect 107168 47354 107192 47356
rect 107248 47354 107272 47356
rect 107328 47354 107334 47356
rect 107088 47302 107090 47354
rect 107270 47302 107272 47354
rect 107026 47300 107032 47302
rect 107088 47300 107112 47302
rect 107168 47300 107192 47302
rect 107248 47300 107272 47302
rect 107328 47300 107334 47302
rect 107026 47291 107334 47300
rect 107762 46812 108070 46821
rect 107762 46810 107768 46812
rect 107824 46810 107848 46812
rect 107904 46810 107928 46812
rect 107984 46810 108008 46812
rect 108064 46810 108070 46812
rect 107824 46758 107826 46810
rect 108006 46758 108008 46810
rect 107762 46756 107768 46758
rect 107824 46756 107848 46758
rect 107904 46756 107928 46758
rect 107984 46756 108008 46758
rect 108064 46756 108070 46758
rect 107762 46747 108070 46756
rect 107026 46268 107334 46277
rect 107026 46266 107032 46268
rect 107088 46266 107112 46268
rect 107168 46266 107192 46268
rect 107248 46266 107272 46268
rect 107328 46266 107334 46268
rect 107088 46214 107090 46266
rect 107270 46214 107272 46266
rect 107026 46212 107032 46214
rect 107088 46212 107112 46214
rect 107168 46212 107192 46214
rect 107248 46212 107272 46214
rect 107328 46212 107334 46214
rect 107026 46203 107334 46212
rect 107762 45724 108070 45733
rect 107762 45722 107768 45724
rect 107824 45722 107848 45724
rect 107904 45722 107928 45724
rect 107984 45722 108008 45724
rect 108064 45722 108070 45724
rect 107824 45670 107826 45722
rect 108006 45670 108008 45722
rect 107762 45668 107768 45670
rect 107824 45668 107848 45670
rect 107904 45668 107928 45670
rect 107984 45668 108008 45670
rect 108064 45668 108070 45670
rect 107762 45659 108070 45668
rect 107026 45180 107334 45189
rect 107026 45178 107032 45180
rect 107088 45178 107112 45180
rect 107168 45178 107192 45180
rect 107248 45178 107272 45180
rect 107328 45178 107334 45180
rect 107088 45126 107090 45178
rect 107270 45126 107272 45178
rect 107026 45124 107032 45126
rect 107088 45124 107112 45126
rect 107168 45124 107192 45126
rect 107248 45124 107272 45126
rect 107328 45124 107334 45126
rect 107026 45115 107334 45124
rect 107762 44636 108070 44645
rect 107762 44634 107768 44636
rect 107824 44634 107848 44636
rect 107904 44634 107928 44636
rect 107984 44634 108008 44636
rect 108064 44634 108070 44636
rect 107824 44582 107826 44634
rect 108006 44582 108008 44634
rect 107762 44580 107768 44582
rect 107824 44580 107848 44582
rect 107904 44580 107928 44582
rect 107984 44580 108008 44582
rect 108064 44580 108070 44582
rect 107762 44571 108070 44580
rect 107026 44092 107334 44101
rect 107026 44090 107032 44092
rect 107088 44090 107112 44092
rect 107168 44090 107192 44092
rect 107248 44090 107272 44092
rect 107328 44090 107334 44092
rect 107088 44038 107090 44090
rect 107270 44038 107272 44090
rect 107026 44036 107032 44038
rect 107088 44036 107112 44038
rect 107168 44036 107192 44038
rect 107248 44036 107272 44038
rect 107328 44036 107334 44038
rect 107026 44027 107334 44036
rect 107762 43548 108070 43557
rect 107762 43546 107768 43548
rect 107824 43546 107848 43548
rect 107904 43546 107928 43548
rect 107984 43546 108008 43548
rect 108064 43546 108070 43548
rect 107824 43494 107826 43546
rect 108006 43494 108008 43546
rect 107762 43492 107768 43494
rect 107824 43492 107848 43494
rect 107904 43492 107928 43494
rect 107984 43492 108008 43494
rect 108064 43492 108070 43494
rect 107762 43483 108070 43492
rect 107026 43004 107334 43013
rect 107026 43002 107032 43004
rect 107088 43002 107112 43004
rect 107168 43002 107192 43004
rect 107248 43002 107272 43004
rect 107328 43002 107334 43004
rect 107088 42950 107090 43002
rect 107270 42950 107272 43002
rect 107026 42948 107032 42950
rect 107088 42948 107112 42950
rect 107168 42948 107192 42950
rect 107248 42948 107272 42950
rect 107328 42948 107334 42950
rect 107026 42939 107334 42948
rect 105452 42560 105504 42566
rect 105452 42502 105504 42508
rect 106372 42560 106424 42566
rect 106372 42502 106424 42508
rect 106096 42220 106148 42226
rect 106096 42162 106148 42168
rect 106108 42022 106136 42162
rect 106384 42022 106412 42502
rect 107762 42460 108070 42469
rect 107762 42458 107768 42460
rect 107824 42458 107848 42460
rect 107904 42458 107928 42460
rect 107984 42458 108008 42460
rect 108064 42458 108070 42460
rect 107824 42406 107826 42458
rect 108006 42406 108008 42458
rect 107762 42404 107768 42406
rect 107824 42404 107848 42406
rect 107904 42404 107928 42406
rect 107984 42404 108008 42406
rect 108064 42404 108070 42406
rect 107762 42395 108070 42404
rect 106096 42016 106148 42022
rect 106096 41958 106148 41964
rect 106372 42016 106424 42022
rect 106372 41958 106424 41964
rect 106108 41546 106136 41958
rect 107026 41916 107334 41925
rect 107026 41914 107032 41916
rect 107088 41914 107112 41916
rect 107168 41914 107192 41916
rect 107248 41914 107272 41916
rect 107328 41914 107334 41916
rect 107088 41862 107090 41914
rect 107270 41862 107272 41914
rect 107026 41860 107032 41862
rect 107088 41860 107112 41862
rect 107168 41860 107192 41862
rect 107248 41860 107272 41862
rect 107328 41860 107334 41862
rect 107026 41851 107334 41860
rect 106096 41540 106148 41546
rect 106096 41482 106148 41488
rect 105176 40928 105228 40934
rect 105176 40870 105228 40876
rect 105912 40928 105964 40934
rect 105912 40870 105964 40876
rect 104532 36916 104584 36922
rect 104532 36858 104584 36864
rect 104544 36802 104572 36858
rect 104544 36774 104664 36802
rect 104532 36576 104584 36582
rect 104532 36518 104584 36524
rect 104440 35488 104492 35494
rect 104440 35430 104492 35436
rect 104452 32842 104480 35430
rect 104544 33930 104572 36518
rect 104636 35894 104664 36774
rect 104636 35866 104756 35894
rect 104728 35698 104756 35866
rect 104716 35692 104768 35698
rect 104716 35634 104768 35640
rect 104728 35494 104756 35634
rect 104716 35488 104768 35494
rect 104716 35430 104768 35436
rect 104532 33924 104584 33930
rect 104532 33866 104584 33872
rect 104440 32836 104492 32842
rect 104440 32778 104492 32784
rect 104532 32768 104584 32774
rect 104584 32716 104664 32722
rect 104532 32710 104664 32716
rect 104544 32694 104664 32710
rect 104532 32360 104584 32366
rect 104532 32302 104584 32308
rect 104544 31822 104572 32302
rect 104636 31822 104664 32694
rect 104728 32366 104756 35430
rect 105820 33924 105872 33930
rect 105820 33866 105872 33872
rect 104808 33856 104860 33862
rect 104808 33798 104860 33804
rect 104820 33454 104848 33798
rect 104808 33448 104860 33454
rect 104808 33390 104860 33396
rect 104716 32360 104768 32366
rect 104716 32302 104768 32308
rect 104716 31952 104768 31958
rect 104716 31894 104768 31900
rect 104532 31816 104584 31822
rect 104532 31758 104584 31764
rect 104624 31816 104676 31822
rect 104624 31758 104676 31764
rect 104544 31142 104572 31758
rect 104532 31136 104584 31142
rect 104532 31078 104584 31084
rect 104440 30320 104492 30326
rect 104440 30262 104492 30268
rect 104256 29504 104308 29510
rect 104256 29446 104308 29452
rect 104268 25974 104296 29446
rect 104452 28150 104480 30262
rect 104544 29646 104572 31078
rect 104532 29640 104584 29646
rect 104532 29582 104584 29588
rect 104532 28484 104584 28490
rect 104532 28426 104584 28432
rect 104440 28144 104492 28150
rect 104440 28086 104492 28092
rect 104348 26308 104400 26314
rect 104348 26250 104400 26256
rect 104256 25968 104308 25974
rect 104256 25910 104308 25916
rect 104360 25906 104388 26250
rect 104348 25900 104400 25906
rect 104348 25842 104400 25848
rect 104452 25242 104480 28086
rect 104544 27130 104572 28426
rect 104636 27826 104664 31758
rect 104728 28490 104756 31894
rect 104820 30326 104848 33390
rect 105636 33312 105688 33318
rect 105636 33254 105688 33260
rect 105452 32972 105504 32978
rect 105452 32914 105504 32920
rect 105360 31816 105412 31822
rect 105360 31758 105412 31764
rect 104808 30320 104860 30326
rect 104808 30262 104860 30268
rect 105372 30258 105400 31758
rect 105360 30252 105412 30258
rect 105360 30194 105412 30200
rect 105464 30122 105492 32914
rect 105648 31822 105676 33254
rect 105832 32026 105860 33866
rect 105820 32020 105872 32026
rect 105820 31962 105872 31968
rect 105924 31958 105952 40870
rect 106108 33998 106136 41482
rect 107762 41372 108070 41381
rect 107762 41370 107768 41372
rect 107824 41370 107848 41372
rect 107904 41370 107928 41372
rect 107984 41370 108008 41372
rect 108064 41370 108070 41372
rect 107824 41318 107826 41370
rect 108006 41318 108008 41370
rect 107762 41316 107768 41318
rect 107824 41316 107848 41318
rect 107904 41316 107928 41318
rect 107984 41316 108008 41318
rect 108064 41316 108070 41318
rect 107762 41307 108070 41316
rect 107026 40828 107334 40837
rect 107026 40826 107032 40828
rect 107088 40826 107112 40828
rect 107168 40826 107192 40828
rect 107248 40826 107272 40828
rect 107328 40826 107334 40828
rect 107088 40774 107090 40826
rect 107270 40774 107272 40826
rect 107026 40772 107032 40774
rect 107088 40772 107112 40774
rect 107168 40772 107192 40774
rect 107248 40772 107272 40774
rect 107328 40772 107334 40774
rect 107026 40763 107334 40772
rect 107762 40284 108070 40293
rect 107762 40282 107768 40284
rect 107824 40282 107848 40284
rect 107904 40282 107928 40284
rect 107984 40282 108008 40284
rect 108064 40282 108070 40284
rect 107824 40230 107826 40282
rect 108006 40230 108008 40282
rect 107762 40228 107768 40230
rect 107824 40228 107848 40230
rect 107904 40228 107928 40230
rect 107984 40228 108008 40230
rect 108064 40228 108070 40230
rect 107762 40219 108070 40228
rect 107026 39740 107334 39749
rect 107026 39738 107032 39740
rect 107088 39738 107112 39740
rect 107168 39738 107192 39740
rect 107248 39738 107272 39740
rect 107328 39738 107334 39740
rect 107088 39686 107090 39738
rect 107270 39686 107272 39738
rect 107026 39684 107032 39686
rect 107088 39684 107112 39686
rect 107168 39684 107192 39686
rect 107248 39684 107272 39686
rect 107328 39684 107334 39686
rect 107026 39675 107334 39684
rect 107762 39196 108070 39205
rect 107762 39194 107768 39196
rect 107824 39194 107848 39196
rect 107904 39194 107928 39196
rect 107984 39194 108008 39196
rect 108064 39194 108070 39196
rect 107824 39142 107826 39194
rect 108006 39142 108008 39194
rect 107762 39140 107768 39142
rect 107824 39140 107848 39142
rect 107904 39140 107928 39142
rect 107984 39140 108008 39142
rect 108064 39140 108070 39142
rect 107762 39131 108070 39140
rect 107026 38652 107334 38661
rect 107026 38650 107032 38652
rect 107088 38650 107112 38652
rect 107168 38650 107192 38652
rect 107248 38650 107272 38652
rect 107328 38650 107334 38652
rect 107088 38598 107090 38650
rect 107270 38598 107272 38650
rect 107026 38596 107032 38598
rect 107088 38596 107112 38598
rect 107168 38596 107192 38598
rect 107248 38596 107272 38598
rect 107328 38596 107334 38598
rect 107026 38587 107334 38596
rect 107762 38108 108070 38117
rect 107762 38106 107768 38108
rect 107824 38106 107848 38108
rect 107904 38106 107928 38108
rect 107984 38106 108008 38108
rect 108064 38106 108070 38108
rect 107824 38054 107826 38106
rect 108006 38054 108008 38106
rect 107762 38052 107768 38054
rect 107824 38052 107848 38054
rect 107904 38052 107928 38054
rect 107984 38052 108008 38054
rect 108064 38052 108070 38054
rect 107762 38043 108070 38052
rect 107026 37564 107334 37573
rect 107026 37562 107032 37564
rect 107088 37562 107112 37564
rect 107168 37562 107192 37564
rect 107248 37562 107272 37564
rect 107328 37562 107334 37564
rect 107088 37510 107090 37562
rect 107270 37510 107272 37562
rect 107026 37508 107032 37510
rect 107088 37508 107112 37510
rect 107168 37508 107192 37510
rect 107248 37508 107272 37510
rect 107328 37508 107334 37510
rect 107026 37499 107334 37508
rect 107762 37020 108070 37029
rect 107762 37018 107768 37020
rect 107824 37018 107848 37020
rect 107904 37018 107928 37020
rect 107984 37018 108008 37020
rect 108064 37018 108070 37020
rect 107824 36966 107826 37018
rect 108006 36966 108008 37018
rect 107762 36964 107768 36966
rect 107824 36964 107848 36966
rect 107904 36964 107928 36966
rect 107984 36964 108008 36966
rect 108064 36964 108070 36966
rect 107762 36955 108070 36964
rect 107026 36476 107334 36485
rect 107026 36474 107032 36476
rect 107088 36474 107112 36476
rect 107168 36474 107192 36476
rect 107248 36474 107272 36476
rect 107328 36474 107334 36476
rect 107088 36422 107090 36474
rect 107270 36422 107272 36474
rect 107026 36420 107032 36422
rect 107088 36420 107112 36422
rect 107168 36420 107192 36422
rect 107248 36420 107272 36422
rect 107328 36420 107334 36422
rect 107026 36411 107334 36420
rect 107762 35932 108070 35941
rect 107762 35930 107768 35932
rect 107824 35930 107848 35932
rect 107904 35930 107928 35932
rect 107984 35930 108008 35932
rect 108064 35930 108070 35932
rect 107824 35878 107826 35930
rect 108006 35878 108008 35930
rect 107762 35876 107768 35878
rect 107824 35876 107848 35878
rect 107904 35876 107928 35878
rect 107984 35876 108008 35878
rect 108064 35876 108070 35878
rect 107762 35867 108070 35876
rect 107026 35388 107334 35397
rect 107026 35386 107032 35388
rect 107088 35386 107112 35388
rect 107168 35386 107192 35388
rect 107248 35386 107272 35388
rect 107328 35386 107334 35388
rect 107088 35334 107090 35386
rect 107270 35334 107272 35386
rect 107026 35332 107032 35334
rect 107088 35332 107112 35334
rect 107168 35332 107192 35334
rect 107248 35332 107272 35334
rect 107328 35332 107334 35334
rect 107026 35323 107334 35332
rect 107762 34844 108070 34853
rect 107762 34842 107768 34844
rect 107824 34842 107848 34844
rect 107904 34842 107928 34844
rect 107984 34842 108008 34844
rect 108064 34842 108070 34844
rect 107824 34790 107826 34842
rect 108006 34790 108008 34842
rect 107762 34788 107768 34790
rect 107824 34788 107848 34790
rect 107904 34788 107928 34790
rect 107984 34788 108008 34790
rect 108064 34788 108070 34790
rect 107762 34779 108070 34788
rect 107026 34300 107334 34309
rect 107026 34298 107032 34300
rect 107088 34298 107112 34300
rect 107168 34298 107192 34300
rect 107248 34298 107272 34300
rect 107328 34298 107334 34300
rect 107088 34246 107090 34298
rect 107270 34246 107272 34298
rect 107026 34244 107032 34246
rect 107088 34244 107112 34246
rect 107168 34244 107192 34246
rect 107248 34244 107272 34246
rect 107328 34244 107334 34246
rect 107026 34235 107334 34244
rect 106096 33992 106148 33998
rect 106096 33934 106148 33940
rect 106188 33856 106240 33862
rect 106188 33798 106240 33804
rect 106200 32910 106228 33798
rect 107762 33756 108070 33765
rect 107762 33754 107768 33756
rect 107824 33754 107848 33756
rect 107904 33754 107928 33756
rect 107984 33754 108008 33756
rect 108064 33754 108070 33756
rect 107824 33702 107826 33754
rect 108006 33702 108008 33754
rect 107762 33700 107768 33702
rect 107824 33700 107848 33702
rect 107904 33700 107928 33702
rect 107984 33700 108008 33702
rect 108064 33700 108070 33702
rect 107762 33691 108070 33700
rect 107026 33212 107334 33221
rect 107026 33210 107032 33212
rect 107088 33210 107112 33212
rect 107168 33210 107192 33212
rect 107248 33210 107272 33212
rect 107328 33210 107334 33212
rect 107088 33158 107090 33210
rect 107270 33158 107272 33210
rect 107026 33156 107032 33158
rect 107088 33156 107112 33158
rect 107168 33156 107192 33158
rect 107248 33156 107272 33158
rect 107328 33156 107334 33158
rect 107026 33147 107334 33156
rect 106188 32904 106240 32910
rect 106188 32846 106240 32852
rect 106372 32768 106424 32774
rect 106372 32710 106424 32716
rect 105912 31952 105964 31958
rect 105912 31894 105964 31900
rect 105636 31816 105688 31822
rect 105636 31758 105688 31764
rect 105924 30326 105952 31894
rect 105912 30320 105964 30326
rect 105912 30262 105964 30268
rect 105452 30116 105504 30122
rect 105452 30058 105504 30064
rect 104808 29504 104860 29510
rect 104808 29446 104860 29452
rect 104716 28484 104768 28490
rect 104716 28426 104768 28432
rect 104716 27872 104768 27878
rect 104636 27820 104716 27826
rect 104636 27814 104768 27820
rect 104636 27798 104756 27814
rect 104532 27124 104584 27130
rect 104532 27066 104584 27072
rect 104636 26234 104664 27798
rect 104716 27124 104768 27130
rect 104716 27066 104768 27072
rect 104544 26206 104664 26234
rect 104544 25498 104572 26206
rect 104624 25832 104676 25838
rect 104624 25774 104676 25780
rect 104532 25492 104584 25498
rect 104532 25434 104584 25440
rect 104360 25226 104480 25242
rect 104348 25220 104480 25226
rect 104400 25214 104480 25220
rect 104348 25162 104400 25168
rect 104256 25152 104308 25158
rect 104162 25120 104218 25129
rect 104256 25094 104308 25100
rect 104162 25055 104218 25064
rect 104176 24818 104204 25055
rect 104164 24812 104216 24818
rect 104164 24754 104216 24760
rect 104164 24132 104216 24138
rect 104164 24074 104216 24080
rect 104176 23798 104204 24074
rect 104164 23792 104216 23798
rect 104164 23734 104216 23740
rect 102784 11756 102836 11762
rect 102784 11698 102836 11704
rect 90364 10056 90416 10062
rect 90364 9998 90416 10004
rect 90376 9897 90404 9998
rect 104176 9994 104204 23734
rect 104268 23202 104296 25094
rect 104360 23361 104388 25162
rect 104440 24064 104492 24070
rect 104440 24006 104492 24012
rect 104452 23730 104480 24006
rect 104440 23724 104492 23730
rect 104440 23666 104492 23672
rect 104346 23352 104402 23361
rect 104346 23287 104402 23296
rect 104268 23174 104480 23202
rect 104348 20868 104400 20874
rect 104348 20810 104400 20816
rect 104256 20392 104308 20398
rect 104256 20334 104308 20340
rect 104268 19718 104296 20334
rect 104256 19712 104308 19718
rect 104256 19654 104308 19660
rect 90732 9988 90784 9994
rect 90732 9930 90784 9936
rect 104164 9988 104216 9994
rect 104164 9930 104216 9936
rect 16026 9888 16082 9897
rect 16026 9823 16082 9832
rect 90362 9888 90418 9897
rect 90362 9823 90418 9832
rect 16040 9654 16068 9823
rect 31574 9752 31630 9761
rect 31574 9687 31630 9696
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 23478 9616 23534 9625
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 16040 7546 16068 9590
rect 23478 9551 23534 9560
rect 30470 9616 30526 9625
rect 30470 9551 30526 9560
rect 23492 7546 23520 9551
rect 25778 8120 25834 8129
rect 25778 8055 25834 8064
rect 28998 8120 29054 8129
rect 28998 8055 29054 8064
rect 24674 7576 24730 7585
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23480 7540 23532 7546
rect 25792 7546 25820 8055
rect 26974 7576 27030 7585
rect 24674 7511 24676 7520
rect 23480 7482 23532 7488
rect 24728 7511 24730 7520
rect 25780 7540 25832 7546
rect 24676 7482 24728 7488
rect 26974 7511 26976 7520
rect 25780 7482 25832 7488
rect 27028 7511 27030 7520
rect 28262 7576 28318 7585
rect 29012 7546 29040 8055
rect 30484 7546 30512 9551
rect 31588 7546 31616 9687
rect 90744 9489 90772 9930
rect 104268 9897 104296 19654
rect 104360 19310 104388 20810
rect 104348 19304 104400 19310
rect 104348 19246 104400 19252
rect 104452 10062 104480 23174
rect 104544 22273 104572 25434
rect 104636 23594 104664 25774
rect 104728 25498 104756 27066
rect 104716 25492 104768 25498
rect 104716 25434 104768 25440
rect 104728 24206 104756 25434
rect 104820 25294 104848 29446
rect 105452 28416 105504 28422
rect 105452 28358 105504 28364
rect 105084 28144 105136 28150
rect 105084 28086 105136 28092
rect 105096 27130 105124 28086
rect 105176 27872 105228 27878
rect 105176 27814 105228 27820
rect 105084 27124 105136 27130
rect 105084 27066 105136 27072
rect 105096 26234 105124 27066
rect 105188 26994 105216 27814
rect 105464 27130 105492 28358
rect 105924 28150 105952 30262
rect 106384 28626 106412 32710
rect 107762 32668 108070 32677
rect 107762 32666 107768 32668
rect 107824 32666 107848 32668
rect 107904 32666 107928 32668
rect 107984 32666 108008 32668
rect 108064 32666 108070 32668
rect 107824 32614 107826 32666
rect 108006 32614 108008 32666
rect 107762 32612 107768 32614
rect 107824 32612 107848 32614
rect 107904 32612 107928 32614
rect 107984 32612 108008 32614
rect 108064 32612 108070 32614
rect 107762 32603 108070 32612
rect 110328 32428 110380 32434
rect 110328 32370 110380 32376
rect 107026 32124 107334 32133
rect 107026 32122 107032 32124
rect 107088 32122 107112 32124
rect 107168 32122 107192 32124
rect 107248 32122 107272 32124
rect 107328 32122 107334 32124
rect 107088 32070 107090 32122
rect 107270 32070 107272 32122
rect 107026 32068 107032 32070
rect 107088 32068 107112 32070
rect 107168 32068 107192 32070
rect 107248 32068 107272 32070
rect 107328 32068 107334 32070
rect 107026 32059 107334 32068
rect 110340 32026 110368 32370
rect 110328 32020 110380 32026
rect 110328 31962 110380 31968
rect 110512 31816 110564 31822
rect 110512 31758 110564 31764
rect 107762 31580 108070 31589
rect 107762 31578 107768 31580
rect 107824 31578 107848 31580
rect 107904 31578 107928 31580
rect 107984 31578 108008 31580
rect 108064 31578 108070 31580
rect 107824 31526 107826 31578
rect 108006 31526 108008 31578
rect 107762 31524 107768 31526
rect 107824 31524 107848 31526
rect 107904 31524 107928 31526
rect 107984 31524 108008 31526
rect 108064 31524 108070 31526
rect 107762 31515 108070 31524
rect 110524 31385 110552 31758
rect 110510 31376 110566 31385
rect 110510 31311 110566 31320
rect 107026 31036 107334 31045
rect 107026 31034 107032 31036
rect 107088 31034 107112 31036
rect 107168 31034 107192 31036
rect 107248 31034 107272 31036
rect 107328 31034 107334 31036
rect 107088 30982 107090 31034
rect 107270 30982 107272 31034
rect 107026 30980 107032 30982
rect 107088 30980 107112 30982
rect 107168 30980 107192 30982
rect 107248 30980 107272 30982
rect 107328 30980 107334 30982
rect 107026 30971 107334 30980
rect 107762 30492 108070 30501
rect 107762 30490 107768 30492
rect 107824 30490 107848 30492
rect 107904 30490 107928 30492
rect 107984 30490 108008 30492
rect 108064 30490 108070 30492
rect 107824 30438 107826 30490
rect 108006 30438 108008 30490
rect 107762 30436 107768 30438
rect 107824 30436 107848 30438
rect 107904 30436 107928 30438
rect 107984 30436 108008 30438
rect 108064 30436 108070 30438
rect 107762 30427 108070 30436
rect 107026 29948 107334 29957
rect 107026 29946 107032 29948
rect 107088 29946 107112 29948
rect 107168 29946 107192 29948
rect 107248 29946 107272 29948
rect 107328 29946 107334 29948
rect 107088 29894 107090 29946
rect 107270 29894 107272 29946
rect 107026 29892 107032 29894
rect 107088 29892 107112 29894
rect 107168 29892 107192 29894
rect 107248 29892 107272 29894
rect 107328 29892 107334 29894
rect 107026 29883 107334 29892
rect 107762 29404 108070 29413
rect 107762 29402 107768 29404
rect 107824 29402 107848 29404
rect 107904 29402 107928 29404
rect 107984 29402 108008 29404
rect 108064 29402 108070 29404
rect 107824 29350 107826 29402
rect 108006 29350 108008 29402
rect 107762 29348 107768 29350
rect 107824 29348 107848 29350
rect 107904 29348 107928 29350
rect 107984 29348 108008 29350
rect 108064 29348 108070 29350
rect 107762 29339 108070 29348
rect 107026 28860 107334 28869
rect 107026 28858 107032 28860
rect 107088 28858 107112 28860
rect 107168 28858 107192 28860
rect 107248 28858 107272 28860
rect 107328 28858 107334 28860
rect 107088 28806 107090 28858
rect 107270 28806 107272 28858
rect 107026 28804 107032 28806
rect 107088 28804 107112 28806
rect 107168 28804 107192 28806
rect 107248 28804 107272 28806
rect 107328 28804 107334 28806
rect 107026 28795 107334 28804
rect 106372 28620 106424 28626
rect 106372 28562 106424 28568
rect 106384 28422 106412 28562
rect 106372 28416 106424 28422
rect 106372 28358 106424 28364
rect 105912 28144 105964 28150
rect 105912 28086 105964 28092
rect 105452 27124 105504 27130
rect 105452 27066 105504 27072
rect 105268 27056 105320 27062
rect 105268 26998 105320 27004
rect 105176 26988 105228 26994
rect 105176 26930 105228 26936
rect 105280 26234 105308 26998
rect 106384 26314 106412 28358
rect 107762 28316 108070 28325
rect 107762 28314 107768 28316
rect 107824 28314 107848 28316
rect 107904 28314 107928 28316
rect 107984 28314 108008 28316
rect 108064 28314 108070 28316
rect 107824 28262 107826 28314
rect 108006 28262 108008 28314
rect 107762 28260 107768 28262
rect 107824 28260 107848 28262
rect 107904 28260 107928 28262
rect 107984 28260 108008 28262
rect 108064 28260 108070 28262
rect 107762 28251 108070 28260
rect 107026 27772 107334 27781
rect 107026 27770 107032 27772
rect 107088 27770 107112 27772
rect 107168 27770 107192 27772
rect 107248 27770 107272 27772
rect 107328 27770 107334 27772
rect 107088 27718 107090 27770
rect 107270 27718 107272 27770
rect 107026 27716 107032 27718
rect 107088 27716 107112 27718
rect 107168 27716 107192 27718
rect 107248 27716 107272 27718
rect 107328 27716 107334 27718
rect 107026 27707 107334 27716
rect 107762 27228 108070 27237
rect 107762 27226 107768 27228
rect 107824 27226 107848 27228
rect 107904 27226 107928 27228
rect 107984 27226 108008 27228
rect 108064 27226 108070 27228
rect 107824 27174 107826 27226
rect 108006 27174 108008 27226
rect 107762 27172 107768 27174
rect 107824 27172 107848 27174
rect 107904 27172 107928 27174
rect 107984 27172 108008 27174
rect 108064 27172 108070 27174
rect 107762 27163 108070 27172
rect 107026 26684 107334 26693
rect 107026 26682 107032 26684
rect 107088 26682 107112 26684
rect 107168 26682 107192 26684
rect 107248 26682 107272 26684
rect 107328 26682 107334 26684
rect 107088 26630 107090 26682
rect 107270 26630 107272 26682
rect 107026 26628 107032 26630
rect 107088 26628 107112 26630
rect 107168 26628 107192 26630
rect 107248 26628 107272 26630
rect 107328 26628 107334 26630
rect 107026 26619 107334 26628
rect 106372 26308 106424 26314
rect 106372 26250 106424 26256
rect 105004 26206 105124 26234
rect 105188 26206 105308 26234
rect 104808 25288 104860 25294
rect 104808 25230 104860 25236
rect 104900 25152 104952 25158
rect 104900 25094 104952 25100
rect 104716 24200 104768 24206
rect 104716 24142 104768 24148
rect 104728 23866 104756 24142
rect 104716 23860 104768 23866
rect 104716 23802 104768 23808
rect 104624 23588 104676 23594
rect 104624 23530 104676 23536
rect 104716 23520 104768 23526
rect 104716 23462 104768 23468
rect 104530 22264 104586 22273
rect 104530 22199 104586 22208
rect 104728 22114 104756 23462
rect 104636 22086 104756 22114
rect 104636 19310 104664 22086
rect 104912 20874 104940 25094
rect 105004 24410 105032 26206
rect 105188 25226 105216 26206
rect 106384 25702 106412 26250
rect 107762 26140 108070 26149
rect 107762 26138 107768 26140
rect 107824 26138 107848 26140
rect 107904 26138 107928 26140
rect 107984 26138 108008 26140
rect 108064 26138 108070 26140
rect 107824 26086 107826 26138
rect 108006 26086 108008 26138
rect 107762 26084 107768 26086
rect 107824 26084 107848 26086
rect 107904 26084 107928 26086
rect 107984 26084 108008 26086
rect 108064 26084 108070 26086
rect 107762 26075 108070 26084
rect 105268 25696 105320 25702
rect 105268 25638 105320 25644
rect 106372 25696 106424 25702
rect 106372 25638 106424 25644
rect 105176 25220 105228 25226
rect 105176 25162 105228 25168
rect 104992 24404 105044 24410
rect 104992 24346 105044 24352
rect 105004 23866 105032 24346
rect 105280 24138 105308 25638
rect 105268 24132 105320 24138
rect 105268 24074 105320 24080
rect 105280 23866 105308 24074
rect 104992 23860 105044 23866
rect 104992 23802 105044 23808
rect 105268 23860 105320 23866
rect 105268 23802 105320 23808
rect 106384 21010 106412 25638
rect 107026 25596 107334 25605
rect 107026 25594 107032 25596
rect 107088 25594 107112 25596
rect 107168 25594 107192 25596
rect 107248 25594 107272 25596
rect 107328 25594 107334 25596
rect 107088 25542 107090 25594
rect 107270 25542 107272 25594
rect 107026 25540 107032 25542
rect 107088 25540 107112 25542
rect 107168 25540 107192 25542
rect 107248 25540 107272 25542
rect 107328 25540 107334 25542
rect 107026 25531 107334 25540
rect 107762 25052 108070 25061
rect 107762 25050 107768 25052
rect 107824 25050 107848 25052
rect 107904 25050 107928 25052
rect 107984 25050 108008 25052
rect 108064 25050 108070 25052
rect 107824 24998 107826 25050
rect 108006 24998 108008 25050
rect 107762 24996 107768 24998
rect 107824 24996 107848 24998
rect 107904 24996 107928 24998
rect 107984 24996 108008 24998
rect 108064 24996 108070 24998
rect 107762 24987 108070 24996
rect 107026 24508 107334 24517
rect 107026 24506 107032 24508
rect 107088 24506 107112 24508
rect 107168 24506 107192 24508
rect 107248 24506 107272 24508
rect 107328 24506 107334 24508
rect 107088 24454 107090 24506
rect 107270 24454 107272 24506
rect 107026 24452 107032 24454
rect 107088 24452 107112 24454
rect 107168 24452 107192 24454
rect 107248 24452 107272 24454
rect 107328 24452 107334 24454
rect 107026 24443 107334 24452
rect 107762 23964 108070 23973
rect 107762 23962 107768 23964
rect 107824 23962 107848 23964
rect 107904 23962 107928 23964
rect 107984 23962 108008 23964
rect 108064 23962 108070 23964
rect 107824 23910 107826 23962
rect 108006 23910 108008 23962
rect 107762 23908 107768 23910
rect 107824 23908 107848 23910
rect 107904 23908 107928 23910
rect 107984 23908 108008 23910
rect 108064 23908 108070 23910
rect 107762 23899 108070 23908
rect 107026 23420 107334 23429
rect 107026 23418 107032 23420
rect 107088 23418 107112 23420
rect 107168 23418 107192 23420
rect 107248 23418 107272 23420
rect 107328 23418 107334 23420
rect 107088 23366 107090 23418
rect 107270 23366 107272 23418
rect 107026 23364 107032 23366
rect 107088 23364 107112 23366
rect 107168 23364 107192 23366
rect 107248 23364 107272 23366
rect 107328 23364 107334 23366
rect 107026 23355 107334 23364
rect 107762 22876 108070 22885
rect 107762 22874 107768 22876
rect 107824 22874 107848 22876
rect 107904 22874 107928 22876
rect 107984 22874 108008 22876
rect 108064 22874 108070 22876
rect 107824 22822 107826 22874
rect 108006 22822 108008 22874
rect 107762 22820 107768 22822
rect 107824 22820 107848 22822
rect 107904 22820 107928 22822
rect 107984 22820 108008 22822
rect 108064 22820 108070 22822
rect 107762 22811 108070 22820
rect 107026 22332 107334 22341
rect 107026 22330 107032 22332
rect 107088 22330 107112 22332
rect 107168 22330 107192 22332
rect 107248 22330 107272 22332
rect 107328 22330 107334 22332
rect 107088 22278 107090 22330
rect 107270 22278 107272 22330
rect 107026 22276 107032 22278
rect 107088 22276 107112 22278
rect 107168 22276 107192 22278
rect 107248 22276 107272 22278
rect 107328 22276 107334 22278
rect 107026 22267 107334 22276
rect 107762 21788 108070 21797
rect 107762 21786 107768 21788
rect 107824 21786 107848 21788
rect 107904 21786 107928 21788
rect 107984 21786 108008 21788
rect 108064 21786 108070 21788
rect 107824 21734 107826 21786
rect 108006 21734 108008 21786
rect 107762 21732 107768 21734
rect 107824 21732 107848 21734
rect 107904 21732 107928 21734
rect 107984 21732 108008 21734
rect 108064 21732 108070 21734
rect 107762 21723 108070 21732
rect 107026 21244 107334 21253
rect 107026 21242 107032 21244
rect 107088 21242 107112 21244
rect 107168 21242 107192 21244
rect 107248 21242 107272 21244
rect 107328 21242 107334 21244
rect 107088 21190 107090 21242
rect 107270 21190 107272 21242
rect 107026 21188 107032 21190
rect 107088 21188 107112 21190
rect 107168 21188 107192 21190
rect 107248 21188 107272 21190
rect 107328 21188 107334 21190
rect 107026 21179 107334 21188
rect 106372 21004 106424 21010
rect 106372 20946 106424 20952
rect 104900 20868 104952 20874
rect 104900 20810 104952 20816
rect 106096 20800 106148 20806
rect 106096 20742 106148 20748
rect 106108 20398 106136 20742
rect 107762 20700 108070 20709
rect 107762 20698 107768 20700
rect 107824 20698 107848 20700
rect 107904 20698 107928 20700
rect 107984 20698 108008 20700
rect 108064 20698 108070 20700
rect 107824 20646 107826 20698
rect 108006 20646 108008 20698
rect 107762 20644 107768 20646
rect 107824 20644 107848 20646
rect 107904 20644 107928 20646
rect 107984 20644 108008 20646
rect 108064 20644 108070 20646
rect 107762 20635 108070 20644
rect 106096 20392 106148 20398
rect 106096 20334 106148 20340
rect 104716 20256 104768 20262
rect 104716 20198 104768 20204
rect 104728 19378 104756 20198
rect 107026 20156 107334 20165
rect 107026 20154 107032 20156
rect 107088 20154 107112 20156
rect 107168 20154 107192 20156
rect 107248 20154 107272 20156
rect 107328 20154 107334 20156
rect 107088 20102 107090 20154
rect 107270 20102 107272 20154
rect 107026 20100 107032 20102
rect 107088 20100 107112 20102
rect 107168 20100 107192 20102
rect 107248 20100 107272 20102
rect 107328 20100 107334 20102
rect 107026 20091 107334 20100
rect 107762 19612 108070 19621
rect 107762 19610 107768 19612
rect 107824 19610 107848 19612
rect 107904 19610 107928 19612
rect 107984 19610 108008 19612
rect 108064 19610 108070 19612
rect 107824 19558 107826 19610
rect 108006 19558 108008 19610
rect 107762 19556 107768 19558
rect 107824 19556 107848 19558
rect 107904 19556 107928 19558
rect 107984 19556 108008 19558
rect 108064 19556 108070 19558
rect 107762 19547 108070 19556
rect 104716 19372 104768 19378
rect 104716 19314 104768 19320
rect 104624 19304 104676 19310
rect 104624 19246 104676 19252
rect 107026 19068 107334 19077
rect 107026 19066 107032 19068
rect 107088 19066 107112 19068
rect 107168 19066 107192 19068
rect 107248 19066 107272 19068
rect 107328 19066 107334 19068
rect 107088 19014 107090 19066
rect 107270 19014 107272 19066
rect 107026 19012 107032 19014
rect 107088 19012 107112 19014
rect 107168 19012 107192 19014
rect 107248 19012 107272 19014
rect 107328 19012 107334 19014
rect 107026 19003 107334 19012
rect 107762 18524 108070 18533
rect 107762 18522 107768 18524
rect 107824 18522 107848 18524
rect 107904 18522 107928 18524
rect 107984 18522 108008 18524
rect 108064 18522 108070 18524
rect 107824 18470 107826 18522
rect 108006 18470 108008 18522
rect 107762 18468 107768 18470
rect 107824 18468 107848 18470
rect 107904 18468 107928 18470
rect 107984 18468 108008 18470
rect 108064 18468 108070 18470
rect 107762 18459 108070 18468
rect 107026 17980 107334 17989
rect 107026 17978 107032 17980
rect 107088 17978 107112 17980
rect 107168 17978 107192 17980
rect 107248 17978 107272 17980
rect 107328 17978 107334 17980
rect 107088 17926 107090 17978
rect 107270 17926 107272 17978
rect 107026 17924 107032 17926
rect 107088 17924 107112 17926
rect 107168 17924 107192 17926
rect 107248 17924 107272 17926
rect 107328 17924 107334 17926
rect 107026 17915 107334 17924
rect 107762 17436 108070 17445
rect 107762 17434 107768 17436
rect 107824 17434 107848 17436
rect 107904 17434 107928 17436
rect 107984 17434 108008 17436
rect 108064 17434 108070 17436
rect 107824 17382 107826 17434
rect 108006 17382 108008 17434
rect 107762 17380 107768 17382
rect 107824 17380 107848 17382
rect 107904 17380 107928 17382
rect 107984 17380 108008 17382
rect 108064 17380 108070 17382
rect 107762 17371 108070 17380
rect 107026 16892 107334 16901
rect 107026 16890 107032 16892
rect 107088 16890 107112 16892
rect 107168 16890 107192 16892
rect 107248 16890 107272 16892
rect 107328 16890 107334 16892
rect 107088 16838 107090 16890
rect 107270 16838 107272 16890
rect 107026 16836 107032 16838
rect 107088 16836 107112 16838
rect 107168 16836 107192 16838
rect 107248 16836 107272 16838
rect 107328 16836 107334 16838
rect 107026 16827 107334 16836
rect 107762 16348 108070 16357
rect 107762 16346 107768 16348
rect 107824 16346 107848 16348
rect 107904 16346 107928 16348
rect 107984 16346 108008 16348
rect 108064 16346 108070 16348
rect 107824 16294 107826 16346
rect 108006 16294 108008 16346
rect 107762 16292 107768 16294
rect 107824 16292 107848 16294
rect 107904 16292 107928 16294
rect 107984 16292 108008 16294
rect 108064 16292 108070 16294
rect 107762 16283 108070 16292
rect 107026 15804 107334 15813
rect 107026 15802 107032 15804
rect 107088 15802 107112 15804
rect 107168 15802 107192 15804
rect 107248 15802 107272 15804
rect 107328 15802 107334 15804
rect 107088 15750 107090 15802
rect 107270 15750 107272 15802
rect 107026 15748 107032 15750
rect 107088 15748 107112 15750
rect 107168 15748 107192 15750
rect 107248 15748 107272 15750
rect 107328 15748 107334 15750
rect 107026 15739 107334 15748
rect 107762 15260 108070 15269
rect 107762 15258 107768 15260
rect 107824 15258 107848 15260
rect 107904 15258 107928 15260
rect 107984 15258 108008 15260
rect 108064 15258 108070 15260
rect 107824 15206 107826 15258
rect 108006 15206 108008 15258
rect 107762 15204 107768 15206
rect 107824 15204 107848 15206
rect 107904 15204 107928 15206
rect 107984 15204 108008 15206
rect 108064 15204 108070 15206
rect 107762 15195 108070 15204
rect 107026 14716 107334 14725
rect 107026 14714 107032 14716
rect 107088 14714 107112 14716
rect 107168 14714 107192 14716
rect 107248 14714 107272 14716
rect 107328 14714 107334 14716
rect 107088 14662 107090 14714
rect 107270 14662 107272 14714
rect 107026 14660 107032 14662
rect 107088 14660 107112 14662
rect 107168 14660 107192 14662
rect 107248 14660 107272 14662
rect 107328 14660 107334 14662
rect 107026 14651 107334 14660
rect 107762 14172 108070 14181
rect 107762 14170 107768 14172
rect 107824 14170 107848 14172
rect 107904 14170 107928 14172
rect 107984 14170 108008 14172
rect 108064 14170 108070 14172
rect 107824 14118 107826 14170
rect 108006 14118 108008 14170
rect 107762 14116 107768 14118
rect 107824 14116 107848 14118
rect 107904 14116 107928 14118
rect 107984 14116 108008 14118
rect 108064 14116 108070 14118
rect 107762 14107 108070 14116
rect 107026 13628 107334 13637
rect 107026 13626 107032 13628
rect 107088 13626 107112 13628
rect 107168 13626 107192 13628
rect 107248 13626 107272 13628
rect 107328 13626 107334 13628
rect 107088 13574 107090 13626
rect 107270 13574 107272 13626
rect 107026 13572 107032 13574
rect 107088 13572 107112 13574
rect 107168 13572 107192 13574
rect 107248 13572 107272 13574
rect 107328 13572 107334 13574
rect 107026 13563 107334 13572
rect 107762 13084 108070 13093
rect 107762 13082 107768 13084
rect 107824 13082 107848 13084
rect 107904 13082 107928 13084
rect 107984 13082 108008 13084
rect 108064 13082 108070 13084
rect 107824 13030 107826 13082
rect 108006 13030 108008 13082
rect 107762 13028 107768 13030
rect 107824 13028 107848 13030
rect 107904 13028 107928 13030
rect 107984 13028 108008 13030
rect 108064 13028 108070 13030
rect 107762 13019 108070 13028
rect 107026 12540 107334 12549
rect 107026 12538 107032 12540
rect 107088 12538 107112 12540
rect 107168 12538 107192 12540
rect 107248 12538 107272 12540
rect 107328 12538 107334 12540
rect 107088 12486 107090 12538
rect 107270 12486 107272 12538
rect 107026 12484 107032 12486
rect 107088 12484 107112 12486
rect 107168 12484 107192 12486
rect 107248 12484 107272 12486
rect 107328 12484 107334 12486
rect 107026 12475 107334 12484
rect 107762 11996 108070 12005
rect 107762 11994 107768 11996
rect 107824 11994 107848 11996
rect 107904 11994 107928 11996
rect 107984 11994 108008 11996
rect 108064 11994 108070 11996
rect 107824 11942 107826 11994
rect 108006 11942 108008 11994
rect 107762 11940 107768 11942
rect 107824 11940 107848 11942
rect 107904 11940 107928 11942
rect 107984 11940 108008 11942
rect 108064 11940 108070 11942
rect 107762 11931 108070 11940
rect 110420 11756 110472 11762
rect 110420 11698 110472 11704
rect 107026 11452 107334 11461
rect 107026 11450 107032 11452
rect 107088 11450 107112 11452
rect 107168 11450 107192 11452
rect 107248 11450 107272 11452
rect 107328 11450 107334 11452
rect 107088 11398 107090 11450
rect 107270 11398 107272 11450
rect 107026 11396 107032 11398
rect 107088 11396 107112 11398
rect 107168 11396 107192 11398
rect 107248 11396 107272 11398
rect 107328 11396 107334 11398
rect 107026 11387 107334 11396
rect 107762 10908 108070 10917
rect 107762 10906 107768 10908
rect 107824 10906 107848 10908
rect 107904 10906 107928 10908
rect 107984 10906 108008 10908
rect 108064 10906 108070 10908
rect 107824 10854 107826 10906
rect 108006 10854 108008 10906
rect 107762 10852 107768 10854
rect 107824 10852 107848 10854
rect 107904 10852 107928 10854
rect 107984 10852 108008 10854
rect 108064 10852 108070 10854
rect 107762 10843 108070 10852
rect 107026 10364 107334 10373
rect 107026 10362 107032 10364
rect 107088 10362 107112 10364
rect 107168 10362 107192 10364
rect 107248 10362 107272 10364
rect 107328 10362 107334 10364
rect 107088 10310 107090 10362
rect 107270 10310 107272 10362
rect 107026 10308 107032 10310
rect 107088 10308 107112 10310
rect 107168 10308 107192 10310
rect 107248 10308 107272 10310
rect 107328 10308 107334 10310
rect 107026 10299 107334 10308
rect 110432 10305 110460 11698
rect 110418 10296 110474 10305
rect 110418 10231 110474 10240
rect 104440 10056 104492 10062
rect 104440 9998 104492 10004
rect 104254 9888 104310 9897
rect 104254 9823 104310 9832
rect 107762 9820 108070 9829
rect 107762 9818 107768 9820
rect 107824 9818 107848 9820
rect 107904 9818 107928 9820
rect 107984 9818 108008 9820
rect 108064 9818 108070 9820
rect 107824 9766 107826 9818
rect 108006 9766 108008 9818
rect 107762 9764 107768 9766
rect 107824 9764 107848 9766
rect 107904 9764 107928 9766
rect 107984 9764 108008 9766
rect 108064 9764 108070 9766
rect 107762 9755 108070 9764
rect 90730 9480 90786 9489
rect 90730 9415 90786 9424
rect 32862 8120 32918 8129
rect 32862 8055 32918 8064
rect 35254 8120 35310 8129
rect 35254 8055 35310 8064
rect 38658 8120 38714 8129
rect 38658 8055 38714 8064
rect 32876 7546 32904 8055
rect 33966 7576 34022 7585
rect 28262 7511 28264 7520
rect 26976 7482 27028 7488
rect 28316 7511 28318 7520
rect 29000 7540 29052 7546
rect 28264 7482 28316 7488
rect 29000 7482 29052 7488
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 31576 7540 31628 7546
rect 31576 7482 31628 7488
rect 32864 7540 32916 7546
rect 35268 7546 35296 8055
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 36358 7576 36414 7585
rect 33966 7511 33968 7520
rect 32864 7482 32916 7488
rect 34020 7511 34022 7520
rect 35256 7540 35308 7546
rect 33968 7482 34020 7488
rect 36084 7540 36136 7546
rect 35308 7500 35480 7528
rect 35256 7482 35308 7488
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 23216 800 23244 7482
rect 24688 6914 24716 7482
rect 24504 6886 24716 6914
rect 24504 800 24532 6886
rect 25792 800 25820 7482
rect 26988 6914 27016 7482
rect 28276 6914 28304 7482
rect 26988 6886 27108 6914
rect 28276 6886 28396 6914
rect 27080 800 27108 6886
rect 28368 800 28396 6886
rect 29012 800 29040 7482
rect 30484 6914 30512 7482
rect 30300 6886 30512 6914
rect 30300 800 30328 6886
rect 31588 800 31616 7482
rect 32876 800 32904 7482
rect 33980 6914 34008 7482
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 33980 6886 34192 6914
rect 34164 800 34192 6886
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35452 800 35480 7500
rect 36358 7511 36360 7520
rect 36084 7482 36136 7488
rect 36412 7511 36414 7520
rect 37462 7576 37518 7585
rect 38672 7546 38700 8055
rect 66314 7644 66622 7653
rect 66314 7642 66320 7644
rect 66376 7642 66400 7644
rect 66456 7642 66480 7644
rect 66536 7642 66560 7644
rect 66616 7642 66622 7644
rect 66376 7590 66378 7642
rect 66558 7590 66560 7642
rect 66314 7588 66320 7590
rect 66376 7588 66400 7590
rect 66456 7588 66480 7590
rect 66536 7588 66560 7590
rect 66616 7588 66622 7590
rect 39854 7576 39910 7585
rect 37462 7511 37464 7520
rect 36360 7482 36412 7488
rect 37516 7511 37518 7520
rect 38660 7540 38712 7546
rect 37464 7482 37516 7488
rect 39854 7511 39856 7520
rect 38660 7482 38712 7488
rect 39908 7511 39910 7520
rect 41050 7576 41106 7585
rect 42154 7576 42210 7585
rect 41050 7511 41052 7520
rect 39856 7482 39908 7488
rect 41104 7511 41106 7520
rect 41880 7540 41932 7546
rect 41052 7482 41104 7488
rect 42154 7511 42156 7520
rect 41880 7482 41932 7488
rect 42208 7511 42210 7520
rect 43350 7576 43406 7585
rect 66314 7579 66622 7588
rect 43350 7511 43352 7520
rect 42156 7482 42208 7488
rect 43404 7511 43406 7520
rect 90546 7576 90602 7585
rect 90744 7546 90772 9415
rect 107026 9276 107334 9285
rect 107026 9274 107032 9276
rect 107088 9274 107112 9276
rect 107168 9274 107192 9276
rect 107248 9274 107272 9276
rect 107328 9274 107334 9276
rect 107088 9222 107090 9274
rect 107270 9222 107272 9274
rect 107026 9220 107032 9222
rect 107088 9220 107112 9222
rect 107168 9220 107192 9222
rect 107248 9220 107272 9222
rect 107328 9220 107334 9222
rect 107026 9211 107334 9220
rect 107762 8732 108070 8741
rect 107762 8730 107768 8732
rect 107824 8730 107848 8732
rect 107904 8730 107928 8732
rect 107984 8730 108008 8732
rect 108064 8730 108070 8732
rect 107824 8678 107826 8730
rect 108006 8678 108008 8730
rect 107762 8676 107768 8678
rect 107824 8676 107848 8678
rect 107904 8676 107928 8678
rect 107984 8676 108008 8678
rect 108064 8676 108070 8678
rect 107762 8667 108070 8676
rect 107026 8188 107334 8197
rect 107026 8186 107032 8188
rect 107088 8186 107112 8188
rect 107168 8186 107192 8188
rect 107248 8186 107272 8188
rect 107328 8186 107334 8188
rect 107088 8134 107090 8186
rect 107270 8134 107272 8186
rect 107026 8132 107032 8134
rect 107088 8132 107112 8134
rect 107168 8132 107192 8134
rect 107248 8132 107272 8134
rect 107328 8132 107334 8134
rect 107026 8123 107334 8132
rect 97034 7644 97342 7653
rect 97034 7642 97040 7644
rect 97096 7642 97120 7644
rect 97176 7642 97200 7644
rect 97256 7642 97280 7644
rect 97336 7642 97342 7644
rect 97096 7590 97098 7642
rect 97278 7590 97280 7642
rect 97034 7588 97040 7590
rect 97096 7588 97120 7590
rect 97176 7588 97200 7590
rect 97256 7588 97280 7590
rect 97336 7588 97342 7590
rect 91006 7576 91062 7585
rect 97034 7579 97342 7588
rect 107762 7644 108070 7653
rect 107762 7642 107768 7644
rect 107824 7642 107848 7644
rect 107904 7642 107928 7644
rect 107984 7642 108008 7644
rect 108064 7642 108070 7644
rect 107824 7590 107826 7642
rect 108006 7590 108008 7642
rect 107762 7588 107768 7590
rect 107824 7588 107848 7590
rect 107904 7588 107928 7590
rect 107984 7588 108008 7590
rect 108064 7588 108070 7590
rect 107762 7579 108070 7588
rect 90546 7511 90548 7520
rect 43352 7482 43404 7488
rect 90600 7511 90602 7520
rect 90732 7540 90784 7546
rect 90548 7482 90600 7488
rect 91006 7511 91008 7520
rect 90732 7482 90784 7488
rect 91060 7511 91062 7520
rect 91008 7482 91060 7488
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36096 800 36124 7482
rect 37476 6914 37504 7482
rect 37384 6886 37504 6914
rect 37384 800 37412 6886
rect 38672 800 38700 7482
rect 39868 6914 39896 7482
rect 41064 6914 41092 7482
rect 39868 6886 39988 6914
rect 41064 6886 41276 6914
rect 39960 800 39988 6886
rect 41248 800 41276 6886
rect 41892 800 41920 7482
rect 43364 6914 43392 7482
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 96374 7100 96682 7109
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7035 96682 7044
rect 107026 7100 107334 7109
rect 107026 7098 107032 7100
rect 107088 7098 107112 7100
rect 107168 7098 107192 7100
rect 107248 7098 107272 7100
rect 107328 7098 107334 7100
rect 107088 7046 107090 7098
rect 107270 7046 107272 7098
rect 107026 7044 107032 7046
rect 107088 7044 107112 7046
rect 107168 7044 107192 7046
rect 107248 7044 107272 7046
rect 107328 7044 107334 7046
rect 107026 7035 107334 7044
rect 43180 6886 43392 6914
rect 43180 800 43208 6886
rect 66314 6556 66622 6565
rect 66314 6554 66320 6556
rect 66376 6554 66400 6556
rect 66456 6554 66480 6556
rect 66536 6554 66560 6556
rect 66616 6554 66622 6556
rect 66376 6502 66378 6554
rect 66558 6502 66560 6554
rect 66314 6500 66320 6502
rect 66376 6500 66400 6502
rect 66456 6500 66480 6502
rect 66536 6500 66560 6502
rect 66616 6500 66622 6502
rect 66314 6491 66622 6500
rect 97034 6556 97342 6565
rect 97034 6554 97040 6556
rect 97096 6554 97120 6556
rect 97176 6554 97200 6556
rect 97256 6554 97280 6556
rect 97336 6554 97342 6556
rect 97096 6502 97098 6554
rect 97278 6502 97280 6554
rect 97034 6500 97040 6502
rect 97096 6500 97120 6502
rect 97176 6500 97200 6502
rect 97256 6500 97280 6502
rect 97336 6500 97342 6502
rect 97034 6491 97342 6500
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 96374 6012 96682 6021
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5947 96682 5956
rect 66314 5468 66622 5477
rect 66314 5466 66320 5468
rect 66376 5466 66400 5468
rect 66456 5466 66480 5468
rect 66536 5466 66560 5468
rect 66616 5466 66622 5468
rect 66376 5414 66378 5466
rect 66558 5414 66560 5466
rect 66314 5412 66320 5414
rect 66376 5412 66400 5414
rect 66456 5412 66480 5414
rect 66536 5412 66560 5414
rect 66616 5412 66622 5414
rect 66314 5403 66622 5412
rect 97034 5468 97342 5477
rect 97034 5466 97040 5468
rect 97096 5466 97120 5468
rect 97176 5466 97200 5468
rect 97256 5466 97280 5468
rect 97336 5466 97342 5468
rect 97096 5414 97098 5466
rect 97278 5414 97280 5466
rect 97034 5412 97040 5414
rect 97096 5412 97120 5414
rect 97176 5412 97200 5414
rect 97256 5412 97280 5414
rect 97336 5412 97342 5414
rect 97034 5403 97342 5412
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 96374 4924 96682 4933
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4859 96682 4868
rect 66314 4380 66622 4389
rect 66314 4378 66320 4380
rect 66376 4378 66400 4380
rect 66456 4378 66480 4380
rect 66536 4378 66560 4380
rect 66616 4378 66622 4380
rect 66376 4326 66378 4378
rect 66558 4326 66560 4378
rect 66314 4324 66320 4326
rect 66376 4324 66400 4326
rect 66456 4324 66480 4326
rect 66536 4324 66560 4326
rect 66616 4324 66622 4326
rect 66314 4315 66622 4324
rect 97034 4380 97342 4389
rect 97034 4378 97040 4380
rect 97096 4378 97120 4380
rect 97176 4378 97200 4380
rect 97256 4378 97280 4380
rect 97336 4378 97342 4380
rect 97096 4326 97098 4378
rect 97278 4326 97280 4378
rect 97034 4324 97040 4326
rect 97096 4324 97120 4326
rect 97176 4324 97200 4326
rect 97256 4324 97280 4326
rect 97336 4324 97342 4326
rect 97034 4315 97342 4324
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 96374 3836 96682 3845
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3771 96682 3780
rect 66314 3292 66622 3301
rect 66314 3290 66320 3292
rect 66376 3290 66400 3292
rect 66456 3290 66480 3292
rect 66536 3290 66560 3292
rect 66616 3290 66622 3292
rect 66376 3238 66378 3290
rect 66558 3238 66560 3290
rect 66314 3236 66320 3238
rect 66376 3236 66400 3238
rect 66456 3236 66480 3238
rect 66536 3236 66560 3238
rect 66616 3236 66622 3238
rect 66314 3227 66622 3236
rect 97034 3292 97342 3301
rect 97034 3290 97040 3292
rect 97096 3290 97120 3292
rect 97176 3290 97200 3292
rect 97256 3290 97280 3292
rect 97336 3290 97342 3292
rect 97096 3238 97098 3290
rect 97278 3238 97280 3290
rect 97034 3236 97040 3238
rect 97096 3236 97120 3238
rect 97176 3236 97200 3238
rect 97256 3236 97280 3238
rect 97336 3236 97342 3238
rect 97034 3227 97342 3236
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 96374 2748 96682 2757
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2683 96682 2692
rect 66314 2204 66622 2213
rect 66314 2202 66320 2204
rect 66376 2202 66400 2204
rect 66456 2202 66480 2204
rect 66536 2202 66560 2204
rect 66616 2202 66622 2204
rect 66376 2150 66378 2202
rect 66558 2150 66560 2202
rect 66314 2148 66320 2150
rect 66376 2148 66400 2150
rect 66456 2148 66480 2150
rect 66536 2148 66560 2150
rect 66616 2148 66622 2150
rect 66314 2139 66622 2148
rect 97034 2204 97342 2213
rect 97034 2202 97040 2204
rect 97096 2202 97120 2204
rect 97176 2202 97200 2204
rect 97256 2202 97280 2204
rect 97336 2202 97342 2204
rect 97096 2150 97098 2202
rect 97278 2150 97280 2202
rect 97034 2148 97040 2150
rect 97096 2148 97120 2150
rect 97176 2148 97200 2150
rect 97256 2148 97280 2150
rect 97336 2148 97342 2150
rect 97034 2139 97342 2148
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 43166 0 43222 800
<< via2 >>
rect 4880 71834 4936 71836
rect 4960 71834 5016 71836
rect 5040 71834 5096 71836
rect 5120 71834 5176 71836
rect 4880 71782 4926 71834
rect 4926 71782 4936 71834
rect 4960 71782 4990 71834
rect 4990 71782 5002 71834
rect 5002 71782 5016 71834
rect 5040 71782 5054 71834
rect 5054 71782 5066 71834
rect 5066 71782 5096 71834
rect 5120 71782 5130 71834
rect 5130 71782 5176 71834
rect 4880 71780 4936 71782
rect 4960 71780 5016 71782
rect 5040 71780 5096 71782
rect 5120 71780 5176 71782
rect 35600 71834 35656 71836
rect 35680 71834 35736 71836
rect 35760 71834 35816 71836
rect 35840 71834 35896 71836
rect 35600 71782 35646 71834
rect 35646 71782 35656 71834
rect 35680 71782 35710 71834
rect 35710 71782 35722 71834
rect 35722 71782 35736 71834
rect 35760 71782 35774 71834
rect 35774 71782 35786 71834
rect 35786 71782 35816 71834
rect 35840 71782 35850 71834
rect 35850 71782 35896 71834
rect 35600 71780 35656 71782
rect 35680 71780 35736 71782
rect 35760 71780 35816 71782
rect 35840 71780 35896 71782
rect 66320 71834 66376 71836
rect 66400 71834 66456 71836
rect 66480 71834 66536 71836
rect 66560 71834 66616 71836
rect 66320 71782 66366 71834
rect 66366 71782 66376 71834
rect 66400 71782 66430 71834
rect 66430 71782 66442 71834
rect 66442 71782 66456 71834
rect 66480 71782 66494 71834
rect 66494 71782 66506 71834
rect 66506 71782 66536 71834
rect 66560 71782 66570 71834
rect 66570 71782 66616 71834
rect 66320 71780 66376 71782
rect 66400 71780 66456 71782
rect 66480 71780 66536 71782
rect 66560 71780 66616 71782
rect 97040 71834 97096 71836
rect 97120 71834 97176 71836
rect 97200 71834 97256 71836
rect 97280 71834 97336 71836
rect 97040 71782 97086 71834
rect 97086 71782 97096 71834
rect 97120 71782 97150 71834
rect 97150 71782 97162 71834
rect 97162 71782 97176 71834
rect 97200 71782 97214 71834
rect 97214 71782 97226 71834
rect 97226 71782 97256 71834
rect 97280 71782 97290 71834
rect 97290 71782 97336 71834
rect 97040 71780 97096 71782
rect 97120 71780 97176 71782
rect 97200 71780 97256 71782
rect 97280 71780 97336 71782
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 34940 71290 34996 71292
rect 35020 71290 35076 71292
rect 35100 71290 35156 71292
rect 35180 71290 35236 71292
rect 34940 71238 34986 71290
rect 34986 71238 34996 71290
rect 35020 71238 35050 71290
rect 35050 71238 35062 71290
rect 35062 71238 35076 71290
rect 35100 71238 35114 71290
rect 35114 71238 35126 71290
rect 35126 71238 35156 71290
rect 35180 71238 35190 71290
rect 35190 71238 35236 71290
rect 34940 71236 34996 71238
rect 35020 71236 35076 71238
rect 35100 71236 35156 71238
rect 35180 71236 35236 71238
rect 4880 70746 4936 70748
rect 4960 70746 5016 70748
rect 5040 70746 5096 70748
rect 5120 70746 5176 70748
rect 4880 70694 4926 70746
rect 4926 70694 4936 70746
rect 4960 70694 4990 70746
rect 4990 70694 5002 70746
rect 5002 70694 5016 70746
rect 5040 70694 5054 70746
rect 5054 70694 5066 70746
rect 5066 70694 5096 70746
rect 5120 70694 5130 70746
rect 5130 70694 5176 70746
rect 4880 70692 4936 70694
rect 4960 70692 5016 70694
rect 5040 70692 5096 70694
rect 5120 70692 5176 70694
rect 35600 70746 35656 70748
rect 35680 70746 35736 70748
rect 35760 70746 35816 70748
rect 35840 70746 35896 70748
rect 35600 70694 35646 70746
rect 35646 70694 35656 70746
rect 35680 70694 35710 70746
rect 35710 70694 35722 70746
rect 35722 70694 35736 70746
rect 35760 70694 35774 70746
rect 35774 70694 35786 70746
rect 35786 70694 35816 70746
rect 35840 70694 35850 70746
rect 35850 70694 35896 70746
rect 35600 70692 35656 70694
rect 35680 70692 35736 70694
rect 35760 70692 35816 70694
rect 35840 70692 35896 70694
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 34940 70202 34996 70204
rect 35020 70202 35076 70204
rect 35100 70202 35156 70204
rect 35180 70202 35236 70204
rect 34940 70150 34986 70202
rect 34986 70150 34996 70202
rect 35020 70150 35050 70202
rect 35050 70150 35062 70202
rect 35062 70150 35076 70202
rect 35100 70150 35114 70202
rect 35114 70150 35126 70202
rect 35126 70150 35156 70202
rect 35180 70150 35190 70202
rect 35190 70150 35236 70202
rect 34940 70148 34996 70150
rect 35020 70148 35076 70150
rect 35100 70148 35156 70150
rect 35180 70148 35236 70150
rect 4880 69658 4936 69660
rect 4960 69658 5016 69660
rect 5040 69658 5096 69660
rect 5120 69658 5176 69660
rect 4880 69606 4926 69658
rect 4926 69606 4936 69658
rect 4960 69606 4990 69658
rect 4990 69606 5002 69658
rect 5002 69606 5016 69658
rect 5040 69606 5054 69658
rect 5054 69606 5066 69658
rect 5066 69606 5096 69658
rect 5120 69606 5130 69658
rect 5130 69606 5176 69658
rect 4880 69604 4936 69606
rect 4960 69604 5016 69606
rect 5040 69604 5096 69606
rect 5120 69604 5176 69606
rect 35600 69658 35656 69660
rect 35680 69658 35736 69660
rect 35760 69658 35816 69660
rect 35840 69658 35896 69660
rect 35600 69606 35646 69658
rect 35646 69606 35656 69658
rect 35680 69606 35710 69658
rect 35710 69606 35722 69658
rect 35722 69606 35736 69658
rect 35760 69606 35774 69658
rect 35774 69606 35786 69658
rect 35786 69606 35816 69658
rect 35840 69606 35850 69658
rect 35850 69606 35896 69658
rect 35600 69604 35656 69606
rect 35680 69604 35736 69606
rect 35760 69604 35816 69606
rect 35840 69604 35896 69606
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 4880 68570 4936 68572
rect 4960 68570 5016 68572
rect 5040 68570 5096 68572
rect 5120 68570 5176 68572
rect 4880 68518 4926 68570
rect 4926 68518 4936 68570
rect 4960 68518 4990 68570
rect 4990 68518 5002 68570
rect 5002 68518 5016 68570
rect 5040 68518 5054 68570
rect 5054 68518 5066 68570
rect 5066 68518 5096 68570
rect 5120 68518 5130 68570
rect 5130 68518 5176 68570
rect 4880 68516 4936 68518
rect 4960 68516 5016 68518
rect 5040 68516 5096 68518
rect 5120 68516 5176 68518
rect 35600 68570 35656 68572
rect 35680 68570 35736 68572
rect 35760 68570 35816 68572
rect 35840 68570 35896 68572
rect 35600 68518 35646 68570
rect 35646 68518 35656 68570
rect 35680 68518 35710 68570
rect 35710 68518 35722 68570
rect 35722 68518 35736 68570
rect 35760 68518 35774 68570
rect 35774 68518 35786 68570
rect 35786 68518 35816 68570
rect 35840 68518 35850 68570
rect 35850 68518 35896 68570
rect 35600 68516 35656 68518
rect 35680 68516 35736 68518
rect 35760 68516 35816 68518
rect 35840 68516 35896 68518
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 4880 67482 4936 67484
rect 4960 67482 5016 67484
rect 5040 67482 5096 67484
rect 5120 67482 5176 67484
rect 4880 67430 4926 67482
rect 4926 67430 4936 67482
rect 4960 67430 4990 67482
rect 4990 67430 5002 67482
rect 5002 67430 5016 67482
rect 5040 67430 5054 67482
rect 5054 67430 5066 67482
rect 5066 67430 5096 67482
rect 5120 67430 5130 67482
rect 5130 67430 5176 67482
rect 4880 67428 4936 67430
rect 4960 67428 5016 67430
rect 5040 67428 5096 67430
rect 5120 67428 5176 67430
rect 35600 67482 35656 67484
rect 35680 67482 35736 67484
rect 35760 67482 35816 67484
rect 35840 67482 35896 67484
rect 35600 67430 35646 67482
rect 35646 67430 35656 67482
rect 35680 67430 35710 67482
rect 35710 67430 35722 67482
rect 35722 67430 35736 67482
rect 35760 67430 35774 67482
rect 35774 67430 35786 67482
rect 35786 67430 35816 67482
rect 35840 67430 35850 67482
rect 35850 67430 35896 67482
rect 35600 67428 35656 67430
rect 35680 67428 35736 67430
rect 35760 67428 35816 67430
rect 35840 67428 35896 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 4880 66394 4936 66396
rect 4960 66394 5016 66396
rect 5040 66394 5096 66396
rect 5120 66394 5176 66396
rect 4880 66342 4926 66394
rect 4926 66342 4936 66394
rect 4960 66342 4990 66394
rect 4990 66342 5002 66394
rect 5002 66342 5016 66394
rect 5040 66342 5054 66394
rect 5054 66342 5066 66394
rect 5066 66342 5096 66394
rect 5120 66342 5130 66394
rect 5130 66342 5176 66394
rect 4880 66340 4936 66342
rect 4960 66340 5016 66342
rect 5040 66340 5096 66342
rect 5120 66340 5176 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 4880 65306 4936 65308
rect 4960 65306 5016 65308
rect 5040 65306 5096 65308
rect 5120 65306 5176 65308
rect 4880 65254 4926 65306
rect 4926 65254 4936 65306
rect 4960 65254 4990 65306
rect 4990 65254 5002 65306
rect 5002 65254 5016 65306
rect 5040 65254 5054 65306
rect 5054 65254 5066 65306
rect 5066 65254 5096 65306
rect 5120 65254 5130 65306
rect 5130 65254 5176 65306
rect 4880 65252 4936 65254
rect 4960 65252 5016 65254
rect 5040 65252 5096 65254
rect 5120 65252 5176 65254
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 4880 64218 4936 64220
rect 4960 64218 5016 64220
rect 5040 64218 5096 64220
rect 5120 64218 5176 64220
rect 4880 64166 4926 64218
rect 4926 64166 4936 64218
rect 4960 64166 4990 64218
rect 4990 64166 5002 64218
rect 5002 64166 5016 64218
rect 5040 64166 5054 64218
rect 5054 64166 5066 64218
rect 5066 64166 5096 64218
rect 5120 64166 5130 64218
rect 5130 64166 5176 64218
rect 4880 64164 4936 64166
rect 4960 64164 5016 64166
rect 5040 64164 5096 64166
rect 5120 64164 5176 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 4880 63130 4936 63132
rect 4960 63130 5016 63132
rect 5040 63130 5096 63132
rect 5120 63130 5176 63132
rect 4880 63078 4926 63130
rect 4926 63078 4936 63130
rect 4960 63078 4990 63130
rect 4990 63078 5002 63130
rect 5002 63078 5016 63130
rect 5040 63078 5054 63130
rect 5054 63078 5066 63130
rect 5066 63078 5096 63130
rect 5120 63078 5130 63130
rect 5130 63078 5176 63130
rect 4880 63076 4936 63078
rect 4960 63076 5016 63078
rect 5040 63076 5096 63078
rect 5120 63076 5176 63078
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 4880 62042 4936 62044
rect 4960 62042 5016 62044
rect 5040 62042 5096 62044
rect 5120 62042 5176 62044
rect 4880 61990 4926 62042
rect 4926 61990 4936 62042
rect 4960 61990 4990 62042
rect 4990 61990 5002 62042
rect 5002 61990 5016 62042
rect 5040 61990 5054 62042
rect 5054 61990 5066 62042
rect 5066 61990 5096 62042
rect 5120 61990 5130 62042
rect 5130 61990 5176 62042
rect 4880 61988 4936 61990
rect 4960 61988 5016 61990
rect 5040 61988 5096 61990
rect 5120 61988 5176 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4880 60954 4936 60956
rect 4960 60954 5016 60956
rect 5040 60954 5096 60956
rect 5120 60954 5176 60956
rect 4880 60902 4926 60954
rect 4926 60902 4936 60954
rect 4960 60902 4990 60954
rect 4990 60902 5002 60954
rect 5002 60902 5016 60954
rect 5040 60902 5054 60954
rect 5054 60902 5066 60954
rect 5066 60902 5096 60954
rect 5120 60902 5130 60954
rect 5130 60902 5176 60954
rect 4880 60900 4936 60902
rect 4960 60900 5016 60902
rect 5040 60900 5096 60902
rect 5120 60900 5176 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4880 59866 4936 59868
rect 4960 59866 5016 59868
rect 5040 59866 5096 59868
rect 5120 59866 5176 59868
rect 4880 59814 4926 59866
rect 4926 59814 4936 59866
rect 4960 59814 4990 59866
rect 4990 59814 5002 59866
rect 5002 59814 5016 59866
rect 5040 59814 5054 59866
rect 5054 59814 5066 59866
rect 5066 59814 5096 59866
rect 5120 59814 5130 59866
rect 5130 59814 5176 59866
rect 4880 59812 4936 59814
rect 4960 59812 5016 59814
rect 5040 59812 5096 59814
rect 5120 59812 5176 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4880 58778 4936 58780
rect 4960 58778 5016 58780
rect 5040 58778 5096 58780
rect 5120 58778 5176 58780
rect 4880 58726 4926 58778
rect 4926 58726 4936 58778
rect 4960 58726 4990 58778
rect 4990 58726 5002 58778
rect 5002 58726 5016 58778
rect 5040 58726 5054 58778
rect 5054 58726 5066 58778
rect 5066 58726 5096 58778
rect 5120 58726 5130 58778
rect 5130 58726 5176 58778
rect 4880 58724 4936 58726
rect 4960 58724 5016 58726
rect 5040 58724 5096 58726
rect 5120 58724 5176 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4880 57690 4936 57692
rect 4960 57690 5016 57692
rect 5040 57690 5096 57692
rect 5120 57690 5176 57692
rect 4880 57638 4926 57690
rect 4926 57638 4936 57690
rect 4960 57638 4990 57690
rect 4990 57638 5002 57690
rect 5002 57638 5016 57690
rect 5040 57638 5054 57690
rect 5054 57638 5066 57690
rect 5066 57638 5096 57690
rect 5120 57638 5130 57690
rect 5130 57638 5176 57690
rect 4880 57636 4936 57638
rect 4960 57636 5016 57638
rect 5040 57636 5096 57638
rect 5120 57636 5176 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4880 56602 4936 56604
rect 4960 56602 5016 56604
rect 5040 56602 5096 56604
rect 5120 56602 5176 56604
rect 4880 56550 4926 56602
rect 4926 56550 4936 56602
rect 4960 56550 4990 56602
rect 4990 56550 5002 56602
rect 5002 56550 5016 56602
rect 5040 56550 5054 56602
rect 5054 56550 5066 56602
rect 5066 56550 5096 56602
rect 5120 56550 5130 56602
rect 5130 56550 5176 56602
rect 4880 56548 4936 56550
rect 4960 56548 5016 56550
rect 5040 56548 5096 56550
rect 5120 56548 5176 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4880 55514 4936 55516
rect 4960 55514 5016 55516
rect 5040 55514 5096 55516
rect 5120 55514 5176 55516
rect 4880 55462 4926 55514
rect 4926 55462 4936 55514
rect 4960 55462 4990 55514
rect 4990 55462 5002 55514
rect 5002 55462 5016 55514
rect 5040 55462 5054 55514
rect 5054 55462 5066 55514
rect 5066 55462 5096 55514
rect 5120 55462 5130 55514
rect 5130 55462 5176 55514
rect 4880 55460 4936 55462
rect 4960 55460 5016 55462
rect 5040 55460 5096 55462
rect 5120 55460 5176 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4880 54426 4936 54428
rect 4960 54426 5016 54428
rect 5040 54426 5096 54428
rect 5120 54426 5176 54428
rect 4880 54374 4926 54426
rect 4926 54374 4936 54426
rect 4960 54374 4990 54426
rect 4990 54374 5002 54426
rect 5002 54374 5016 54426
rect 5040 54374 5054 54426
rect 5054 54374 5066 54426
rect 5066 54374 5096 54426
rect 5120 54374 5130 54426
rect 5130 54374 5176 54426
rect 4880 54372 4936 54374
rect 4960 54372 5016 54374
rect 5040 54372 5096 54374
rect 5120 54372 5176 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4880 53338 4936 53340
rect 4960 53338 5016 53340
rect 5040 53338 5096 53340
rect 5120 53338 5176 53340
rect 4880 53286 4926 53338
rect 4926 53286 4936 53338
rect 4960 53286 4990 53338
rect 4990 53286 5002 53338
rect 5002 53286 5016 53338
rect 5040 53286 5054 53338
rect 5054 53286 5066 53338
rect 5066 53286 5096 53338
rect 5120 53286 5130 53338
rect 5130 53286 5176 53338
rect 4880 53284 4936 53286
rect 4960 53284 5016 53286
rect 5040 53284 5096 53286
rect 5120 53284 5176 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4880 52250 4936 52252
rect 4960 52250 5016 52252
rect 5040 52250 5096 52252
rect 5120 52250 5176 52252
rect 4880 52198 4926 52250
rect 4926 52198 4936 52250
rect 4960 52198 4990 52250
rect 4990 52198 5002 52250
rect 5002 52198 5016 52250
rect 5040 52198 5054 52250
rect 5054 52198 5066 52250
rect 5066 52198 5096 52250
rect 5120 52198 5130 52250
rect 5130 52198 5176 52250
rect 4880 52196 4936 52198
rect 4960 52196 5016 52198
rect 5040 52196 5096 52198
rect 5120 52196 5176 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4880 51162 4936 51164
rect 4960 51162 5016 51164
rect 5040 51162 5096 51164
rect 5120 51162 5176 51164
rect 4880 51110 4926 51162
rect 4926 51110 4936 51162
rect 4960 51110 4990 51162
rect 4990 51110 5002 51162
rect 5002 51110 5016 51162
rect 5040 51110 5054 51162
rect 5054 51110 5066 51162
rect 5066 51110 5096 51162
rect 5120 51110 5130 51162
rect 5130 51110 5176 51162
rect 4880 51108 4936 51110
rect 4960 51108 5016 51110
rect 5040 51108 5096 51110
rect 5120 51108 5176 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4880 50074 4936 50076
rect 4960 50074 5016 50076
rect 5040 50074 5096 50076
rect 5120 50074 5176 50076
rect 4880 50022 4926 50074
rect 4926 50022 4936 50074
rect 4960 50022 4990 50074
rect 4990 50022 5002 50074
rect 5002 50022 5016 50074
rect 5040 50022 5054 50074
rect 5054 50022 5066 50074
rect 5066 50022 5096 50074
rect 5120 50022 5130 50074
rect 5130 50022 5176 50074
rect 4880 50020 4936 50022
rect 4960 50020 5016 50022
rect 5040 50020 5096 50022
rect 5120 50020 5176 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4880 48986 4936 48988
rect 4960 48986 5016 48988
rect 5040 48986 5096 48988
rect 5120 48986 5176 48988
rect 4880 48934 4926 48986
rect 4926 48934 4936 48986
rect 4960 48934 4990 48986
rect 4990 48934 5002 48986
rect 5002 48934 5016 48986
rect 5040 48934 5054 48986
rect 5054 48934 5066 48986
rect 5066 48934 5096 48986
rect 5120 48934 5130 48986
rect 5130 48934 5176 48986
rect 4880 48932 4936 48934
rect 4960 48932 5016 48934
rect 5040 48932 5096 48934
rect 5120 48932 5176 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4880 47898 4936 47900
rect 4960 47898 5016 47900
rect 5040 47898 5096 47900
rect 5120 47898 5176 47900
rect 4880 47846 4926 47898
rect 4926 47846 4936 47898
rect 4960 47846 4990 47898
rect 4990 47846 5002 47898
rect 5002 47846 5016 47898
rect 5040 47846 5054 47898
rect 5054 47846 5066 47898
rect 5066 47846 5096 47898
rect 5120 47846 5130 47898
rect 5130 47846 5176 47898
rect 4880 47844 4936 47846
rect 4960 47844 5016 47846
rect 5040 47844 5096 47846
rect 5120 47844 5176 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4880 46810 4936 46812
rect 4960 46810 5016 46812
rect 5040 46810 5096 46812
rect 5120 46810 5176 46812
rect 4880 46758 4926 46810
rect 4926 46758 4936 46810
rect 4960 46758 4990 46810
rect 4990 46758 5002 46810
rect 5002 46758 5016 46810
rect 5040 46758 5054 46810
rect 5054 46758 5066 46810
rect 5066 46758 5096 46810
rect 5120 46758 5130 46810
rect 5130 46758 5176 46810
rect 4880 46756 4936 46758
rect 4960 46756 5016 46758
rect 5040 46756 5096 46758
rect 5120 46756 5176 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4880 45722 4936 45724
rect 4960 45722 5016 45724
rect 5040 45722 5096 45724
rect 5120 45722 5176 45724
rect 4880 45670 4926 45722
rect 4926 45670 4936 45722
rect 4960 45670 4990 45722
rect 4990 45670 5002 45722
rect 5002 45670 5016 45722
rect 5040 45670 5054 45722
rect 5054 45670 5066 45722
rect 5066 45670 5096 45722
rect 5120 45670 5130 45722
rect 5130 45670 5176 45722
rect 4880 45668 4936 45670
rect 4960 45668 5016 45670
rect 5040 45668 5096 45670
rect 5120 45668 5176 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4880 44634 4936 44636
rect 4960 44634 5016 44636
rect 5040 44634 5096 44636
rect 5120 44634 5176 44636
rect 4880 44582 4926 44634
rect 4926 44582 4936 44634
rect 4960 44582 4990 44634
rect 4990 44582 5002 44634
rect 5002 44582 5016 44634
rect 5040 44582 5054 44634
rect 5054 44582 5066 44634
rect 5066 44582 5096 44634
rect 5120 44582 5130 44634
rect 5130 44582 5176 44634
rect 4880 44580 4936 44582
rect 4960 44580 5016 44582
rect 5040 44580 5096 44582
rect 5120 44580 5176 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 7562 41248 7618 41304
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 7562 39480 7618 39536
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 7562 38256 7618 38312
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 7562 36780 7618 36816
rect 7562 36760 7564 36780
rect 7564 36760 7616 36780
rect 7616 36760 7618 36780
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 7562 35556 7618 35592
rect 7562 35536 7564 35556
rect 7564 35536 7616 35556
rect 7616 35536 7618 35556
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 7562 34060 7618 34096
rect 7562 34040 7564 34060
rect 7564 34040 7616 34060
rect 7616 34040 7618 34060
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 7562 15564 7618 15600
rect 7562 15544 7564 15564
rect 7564 15544 7616 15564
rect 7616 15544 7618 15564
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 35600 66394 35656 66396
rect 35680 66394 35736 66396
rect 35760 66394 35816 66396
rect 35840 66394 35896 66396
rect 35600 66342 35646 66394
rect 35646 66342 35656 66394
rect 35680 66342 35710 66394
rect 35710 66342 35722 66394
rect 35722 66342 35736 66394
rect 35760 66342 35774 66394
rect 35774 66342 35786 66394
rect 35786 66342 35816 66394
rect 35840 66342 35850 66394
rect 35850 66342 35896 66394
rect 35600 66340 35656 66342
rect 35680 66340 35736 66342
rect 35760 66340 35816 66342
rect 35840 66340 35896 66342
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 43166 64096 43222 64152
rect 49698 66272 49754 66328
rect 53654 66408 53710 66464
rect 55678 66680 55734 66736
rect 49974 64096 50030 64152
rect 47582 63960 47638 64016
rect 60002 66408 60058 66464
rect 61658 66272 61714 66328
rect 65660 71290 65716 71292
rect 65740 71290 65796 71292
rect 65820 71290 65876 71292
rect 65900 71290 65956 71292
rect 65660 71238 65706 71290
rect 65706 71238 65716 71290
rect 65740 71238 65770 71290
rect 65770 71238 65782 71290
rect 65782 71238 65796 71290
rect 65820 71238 65834 71290
rect 65834 71238 65846 71290
rect 65846 71238 65876 71290
rect 65900 71238 65910 71290
rect 65910 71238 65956 71290
rect 65660 71236 65716 71238
rect 65740 71236 65796 71238
rect 65820 71236 65876 71238
rect 65900 71236 65956 71238
rect 66320 70746 66376 70748
rect 66400 70746 66456 70748
rect 66480 70746 66536 70748
rect 66560 70746 66616 70748
rect 66320 70694 66366 70746
rect 66366 70694 66376 70746
rect 66400 70694 66430 70746
rect 66430 70694 66442 70746
rect 66442 70694 66456 70746
rect 66480 70694 66494 70746
rect 66494 70694 66506 70746
rect 66506 70694 66536 70746
rect 66560 70694 66570 70746
rect 66570 70694 66616 70746
rect 66320 70692 66376 70694
rect 66400 70692 66456 70694
rect 66480 70692 66536 70694
rect 66560 70692 66616 70694
rect 65660 70202 65716 70204
rect 65740 70202 65796 70204
rect 65820 70202 65876 70204
rect 65900 70202 65956 70204
rect 65660 70150 65706 70202
rect 65706 70150 65716 70202
rect 65740 70150 65770 70202
rect 65770 70150 65782 70202
rect 65782 70150 65796 70202
rect 65820 70150 65834 70202
rect 65834 70150 65846 70202
rect 65846 70150 65876 70202
rect 65900 70150 65910 70202
rect 65910 70150 65956 70202
rect 65660 70148 65716 70150
rect 65740 70148 65796 70150
rect 65820 70148 65876 70150
rect 65900 70148 65956 70150
rect 66320 69658 66376 69660
rect 66400 69658 66456 69660
rect 66480 69658 66536 69660
rect 66560 69658 66616 69660
rect 66320 69606 66366 69658
rect 66366 69606 66376 69658
rect 66400 69606 66430 69658
rect 66430 69606 66442 69658
rect 66442 69606 66456 69658
rect 66480 69606 66494 69658
rect 66494 69606 66506 69658
rect 66506 69606 66536 69658
rect 66560 69606 66570 69658
rect 66570 69606 66616 69658
rect 66320 69604 66376 69606
rect 66400 69604 66456 69606
rect 66480 69604 66536 69606
rect 66560 69604 66616 69606
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 66320 68570 66376 68572
rect 66400 68570 66456 68572
rect 66480 68570 66536 68572
rect 66560 68570 66616 68572
rect 66320 68518 66366 68570
rect 66366 68518 66376 68570
rect 66400 68518 66430 68570
rect 66430 68518 66442 68570
rect 66442 68518 66456 68570
rect 66480 68518 66494 68570
rect 66494 68518 66506 68570
rect 66506 68518 66536 68570
rect 66560 68518 66570 68570
rect 66570 68518 66616 68570
rect 66320 68516 66376 68518
rect 66400 68516 66456 68518
rect 66480 68516 66536 68518
rect 66560 68516 66616 68518
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 66320 67482 66376 67484
rect 66400 67482 66456 67484
rect 66480 67482 66536 67484
rect 66560 67482 66616 67484
rect 66320 67430 66366 67482
rect 66366 67430 66376 67482
rect 66400 67430 66430 67482
rect 66430 67430 66442 67482
rect 66442 67430 66456 67482
rect 66480 67430 66494 67482
rect 66494 67430 66506 67482
rect 66506 67430 66536 67482
rect 66560 67430 66570 67482
rect 66570 67430 66616 67482
rect 66320 67428 66376 67430
rect 66400 67428 66456 67430
rect 66480 67428 66536 67430
rect 66560 67428 66616 67430
rect 63958 66408 64014 66464
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 66320 66394 66376 66396
rect 66400 66394 66456 66396
rect 66480 66394 66536 66396
rect 66560 66394 66616 66396
rect 66320 66342 66366 66394
rect 66366 66342 66376 66394
rect 66400 66342 66430 66394
rect 66430 66342 66442 66394
rect 66442 66342 66456 66394
rect 66480 66342 66494 66394
rect 66494 66342 66506 66394
rect 66506 66342 66536 66394
rect 66560 66342 66570 66394
rect 66570 66342 66616 66394
rect 66320 66340 66376 66342
rect 66400 66340 66456 66342
rect 66480 66340 66536 66342
rect 66560 66340 66616 66342
rect 68466 66544 68522 66600
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 64694 65456 64750 65512
rect 68742 65320 68798 65376
rect 96380 71290 96436 71292
rect 96460 71290 96516 71292
rect 96540 71290 96596 71292
rect 96620 71290 96676 71292
rect 96380 71238 96426 71290
rect 96426 71238 96436 71290
rect 96460 71238 96490 71290
rect 96490 71238 96502 71290
rect 96502 71238 96516 71290
rect 96540 71238 96554 71290
rect 96554 71238 96566 71290
rect 96566 71238 96596 71290
rect 96620 71238 96630 71290
rect 96630 71238 96676 71290
rect 96380 71236 96436 71238
rect 96460 71236 96516 71238
rect 96540 71236 96596 71238
rect 96620 71236 96676 71238
rect 97040 70746 97096 70748
rect 97120 70746 97176 70748
rect 97200 70746 97256 70748
rect 97280 70746 97336 70748
rect 97040 70694 97086 70746
rect 97086 70694 97096 70746
rect 97120 70694 97150 70746
rect 97150 70694 97162 70746
rect 97162 70694 97176 70746
rect 97200 70694 97214 70746
rect 97214 70694 97226 70746
rect 97226 70694 97256 70746
rect 97280 70694 97290 70746
rect 97290 70694 97336 70746
rect 97040 70692 97096 70694
rect 97120 70692 97176 70694
rect 97200 70692 97256 70694
rect 97280 70692 97336 70694
rect 96380 70202 96436 70204
rect 96460 70202 96516 70204
rect 96540 70202 96596 70204
rect 96620 70202 96676 70204
rect 96380 70150 96426 70202
rect 96426 70150 96436 70202
rect 96460 70150 96490 70202
rect 96490 70150 96502 70202
rect 96502 70150 96516 70202
rect 96540 70150 96554 70202
rect 96554 70150 96566 70202
rect 96566 70150 96596 70202
rect 96620 70150 96630 70202
rect 96630 70150 96676 70202
rect 96380 70148 96436 70150
rect 96460 70148 96516 70150
rect 96540 70148 96596 70150
rect 96620 70148 96676 70150
rect 97040 69658 97096 69660
rect 97120 69658 97176 69660
rect 97200 69658 97256 69660
rect 97280 69658 97336 69660
rect 97040 69606 97086 69658
rect 97086 69606 97096 69658
rect 97120 69606 97150 69658
rect 97150 69606 97162 69658
rect 97162 69606 97176 69658
rect 97200 69606 97214 69658
rect 97214 69606 97226 69658
rect 97226 69606 97256 69658
rect 97280 69606 97290 69658
rect 97290 69606 97336 69658
rect 97040 69604 97096 69606
rect 97120 69604 97176 69606
rect 97200 69604 97256 69606
rect 97280 69604 97336 69606
rect 96380 69114 96436 69116
rect 96460 69114 96516 69116
rect 96540 69114 96596 69116
rect 96620 69114 96676 69116
rect 96380 69062 96426 69114
rect 96426 69062 96436 69114
rect 96460 69062 96490 69114
rect 96490 69062 96502 69114
rect 96502 69062 96516 69114
rect 96540 69062 96554 69114
rect 96554 69062 96566 69114
rect 96566 69062 96596 69114
rect 96620 69062 96630 69114
rect 96630 69062 96676 69114
rect 96380 69060 96436 69062
rect 96460 69060 96516 69062
rect 96540 69060 96596 69062
rect 96620 69060 96676 69062
rect 97040 68570 97096 68572
rect 97120 68570 97176 68572
rect 97200 68570 97256 68572
rect 97280 68570 97336 68572
rect 97040 68518 97086 68570
rect 97086 68518 97096 68570
rect 97120 68518 97150 68570
rect 97150 68518 97162 68570
rect 97162 68518 97176 68570
rect 97200 68518 97214 68570
rect 97214 68518 97226 68570
rect 97226 68518 97256 68570
rect 97280 68518 97290 68570
rect 97290 68518 97336 68570
rect 97040 68516 97096 68518
rect 97120 68516 97176 68518
rect 97200 68516 97256 68518
rect 97280 68516 97336 68518
rect 96380 68026 96436 68028
rect 96460 68026 96516 68028
rect 96540 68026 96596 68028
rect 96620 68026 96676 68028
rect 96380 67974 96426 68026
rect 96426 67974 96436 68026
rect 96460 67974 96490 68026
rect 96490 67974 96502 68026
rect 96502 67974 96516 68026
rect 96540 67974 96554 68026
rect 96554 67974 96566 68026
rect 96566 67974 96596 68026
rect 96620 67974 96630 68026
rect 96630 67974 96676 68026
rect 96380 67972 96436 67974
rect 96460 67972 96516 67974
rect 96540 67972 96596 67974
rect 96620 67972 96676 67974
rect 97040 67482 97096 67484
rect 97120 67482 97176 67484
rect 97200 67482 97256 67484
rect 97280 67482 97336 67484
rect 97040 67430 97086 67482
rect 97086 67430 97096 67482
rect 97120 67430 97150 67482
rect 97150 67430 97162 67482
rect 97162 67430 97176 67482
rect 97200 67430 97214 67482
rect 97214 67430 97226 67482
rect 97226 67430 97256 67482
rect 97280 67430 97290 67482
rect 97290 67430 97336 67482
rect 97040 67428 97096 67430
rect 97120 67428 97176 67430
rect 97200 67428 97256 67430
rect 97280 67428 97336 67430
rect 96380 66938 96436 66940
rect 96460 66938 96516 66940
rect 96540 66938 96596 66940
rect 96620 66938 96676 66940
rect 96380 66886 96426 66938
rect 96426 66886 96436 66938
rect 96460 66886 96490 66938
rect 96490 66886 96502 66938
rect 96502 66886 96516 66938
rect 96540 66886 96554 66938
rect 96554 66886 96566 66938
rect 96566 66886 96596 66938
rect 96620 66886 96630 66938
rect 96630 66886 96676 66938
rect 96380 66884 96436 66886
rect 96460 66884 96516 66886
rect 96540 66884 96596 66886
rect 96620 66884 96676 66886
rect 97040 66394 97096 66396
rect 97120 66394 97176 66396
rect 97200 66394 97256 66396
rect 97280 66394 97336 66396
rect 97040 66342 97086 66394
rect 97086 66342 97096 66394
rect 97120 66342 97150 66394
rect 97150 66342 97162 66394
rect 97162 66342 97176 66394
rect 97200 66342 97214 66394
rect 97214 66342 97226 66394
rect 97226 66342 97256 66394
rect 97280 66342 97290 66394
rect 97290 66342 97336 66394
rect 97040 66340 97096 66342
rect 97120 66340 97176 66342
rect 97200 66340 97256 66342
rect 97280 66340 97336 66342
rect 107768 66394 107824 66396
rect 107848 66394 107904 66396
rect 107928 66394 107984 66396
rect 108008 66394 108064 66396
rect 107768 66342 107814 66394
rect 107814 66342 107824 66394
rect 107848 66342 107878 66394
rect 107878 66342 107890 66394
rect 107890 66342 107904 66394
rect 107928 66342 107942 66394
rect 107942 66342 107954 66394
rect 107954 66342 107984 66394
rect 108008 66342 108018 66394
rect 108018 66342 108064 66394
rect 107768 66340 107824 66342
rect 107848 66340 107904 66342
rect 107928 66340 107984 66342
rect 108008 66340 108064 66342
rect 74078 65320 74134 65376
rect 71226 65048 71282 65104
rect 87326 65320 87382 65376
rect 86314 63960 86370 64016
rect 96380 65850 96436 65852
rect 96460 65850 96516 65852
rect 96540 65850 96596 65852
rect 96620 65850 96676 65852
rect 96380 65798 96426 65850
rect 96426 65798 96436 65850
rect 96460 65798 96490 65850
rect 96490 65798 96502 65850
rect 96502 65798 96516 65850
rect 96540 65798 96554 65850
rect 96554 65798 96566 65850
rect 96566 65798 96596 65850
rect 96620 65798 96630 65850
rect 96630 65798 96676 65850
rect 96380 65796 96436 65798
rect 96460 65796 96516 65798
rect 96540 65796 96596 65798
rect 96620 65796 96676 65798
rect 45374 63824 45430 63880
rect 58162 63824 58218 63880
rect 95882 63824 95938 63880
rect 107032 65850 107088 65852
rect 107112 65850 107168 65852
rect 107192 65850 107248 65852
rect 107272 65850 107328 65852
rect 107032 65798 107078 65850
rect 107078 65798 107088 65850
rect 107112 65798 107142 65850
rect 107142 65798 107154 65850
rect 107154 65798 107168 65850
rect 107192 65798 107206 65850
rect 107206 65798 107218 65850
rect 107218 65798 107248 65850
rect 107272 65798 107282 65850
rect 107282 65798 107328 65850
rect 107032 65796 107088 65798
rect 107112 65796 107168 65798
rect 107192 65796 107248 65798
rect 107272 65796 107328 65798
rect 107768 65306 107824 65308
rect 107848 65306 107904 65308
rect 107928 65306 107984 65308
rect 108008 65306 108064 65308
rect 107768 65254 107814 65306
rect 107814 65254 107824 65306
rect 107848 65254 107878 65306
rect 107878 65254 107890 65306
rect 107890 65254 107904 65306
rect 107928 65254 107942 65306
rect 107942 65254 107954 65306
rect 107954 65254 107984 65306
rect 108008 65254 108018 65306
rect 108018 65254 108064 65306
rect 107768 65252 107824 65254
rect 107848 65252 107904 65254
rect 107928 65252 107984 65254
rect 108008 65252 108064 65254
rect 107032 64762 107088 64764
rect 107112 64762 107168 64764
rect 107192 64762 107248 64764
rect 107272 64762 107328 64764
rect 107032 64710 107078 64762
rect 107078 64710 107088 64762
rect 107112 64710 107142 64762
rect 107142 64710 107154 64762
rect 107154 64710 107168 64762
rect 107192 64710 107206 64762
rect 107206 64710 107218 64762
rect 107218 64710 107248 64762
rect 107272 64710 107282 64762
rect 107282 64710 107328 64762
rect 107032 64708 107088 64710
rect 107112 64708 107168 64710
rect 107192 64708 107248 64710
rect 107272 64708 107328 64710
rect 104346 63824 104402 63880
rect 103702 59744 103758 59800
rect 107768 64218 107824 64220
rect 107848 64218 107904 64220
rect 107928 64218 107984 64220
rect 108008 64218 108064 64220
rect 107768 64166 107814 64218
rect 107814 64166 107824 64218
rect 107848 64166 107878 64218
rect 107878 64166 107890 64218
rect 107890 64166 107904 64218
rect 107928 64166 107942 64218
rect 107942 64166 107954 64218
rect 107954 64166 107984 64218
rect 108008 64166 108018 64218
rect 108018 64166 108064 64218
rect 107768 64164 107824 64166
rect 107848 64164 107904 64166
rect 107928 64164 107984 64166
rect 108008 64164 108064 64166
rect 104990 64096 105046 64152
rect 106186 63960 106242 64016
rect 107032 63674 107088 63676
rect 107112 63674 107168 63676
rect 107192 63674 107248 63676
rect 107272 63674 107328 63676
rect 107032 63622 107078 63674
rect 107078 63622 107088 63674
rect 107112 63622 107142 63674
rect 107142 63622 107154 63674
rect 107154 63622 107168 63674
rect 107192 63622 107206 63674
rect 107206 63622 107218 63674
rect 107218 63622 107248 63674
rect 107272 63622 107282 63674
rect 107282 63622 107328 63674
rect 107032 63620 107088 63622
rect 107112 63620 107168 63622
rect 107192 63620 107248 63622
rect 107272 63620 107328 63622
rect 107768 63130 107824 63132
rect 107848 63130 107904 63132
rect 107928 63130 107984 63132
rect 108008 63130 108064 63132
rect 107768 63078 107814 63130
rect 107814 63078 107824 63130
rect 107848 63078 107878 63130
rect 107878 63078 107890 63130
rect 107890 63078 107904 63130
rect 107928 63078 107942 63130
rect 107942 63078 107954 63130
rect 107954 63078 107984 63130
rect 108008 63078 108018 63130
rect 108018 63078 108064 63130
rect 107768 63076 107824 63078
rect 107848 63076 107904 63078
rect 107928 63076 107984 63078
rect 108008 63076 108064 63078
rect 107032 62586 107088 62588
rect 107112 62586 107168 62588
rect 107192 62586 107248 62588
rect 107272 62586 107328 62588
rect 107032 62534 107078 62586
rect 107078 62534 107088 62586
rect 107112 62534 107142 62586
rect 107142 62534 107154 62586
rect 107154 62534 107168 62586
rect 107192 62534 107206 62586
rect 107206 62534 107218 62586
rect 107218 62534 107248 62586
rect 107272 62534 107282 62586
rect 107282 62534 107328 62586
rect 107032 62532 107088 62534
rect 107112 62532 107168 62534
rect 107192 62532 107248 62534
rect 107272 62532 107328 62534
rect 107768 62042 107824 62044
rect 107848 62042 107904 62044
rect 107928 62042 107984 62044
rect 108008 62042 108064 62044
rect 107768 61990 107814 62042
rect 107814 61990 107824 62042
rect 107848 61990 107878 62042
rect 107878 61990 107890 62042
rect 107890 61990 107904 62042
rect 107928 61990 107942 62042
rect 107942 61990 107954 62042
rect 107954 61990 107984 62042
rect 108008 61990 108018 62042
rect 108018 61990 108064 62042
rect 107768 61988 107824 61990
rect 107848 61988 107904 61990
rect 107928 61988 107984 61990
rect 108008 61988 108064 61990
rect 107032 61498 107088 61500
rect 107112 61498 107168 61500
rect 107192 61498 107248 61500
rect 107272 61498 107328 61500
rect 107032 61446 107078 61498
rect 107078 61446 107088 61498
rect 107112 61446 107142 61498
rect 107142 61446 107154 61498
rect 107154 61446 107168 61498
rect 107192 61446 107206 61498
rect 107206 61446 107218 61498
rect 107218 61446 107248 61498
rect 107272 61446 107282 61498
rect 107282 61446 107328 61498
rect 107032 61444 107088 61446
rect 107112 61444 107168 61446
rect 107192 61444 107248 61446
rect 107272 61444 107328 61446
rect 107768 60954 107824 60956
rect 107848 60954 107904 60956
rect 107928 60954 107984 60956
rect 108008 60954 108064 60956
rect 107768 60902 107814 60954
rect 107814 60902 107824 60954
rect 107848 60902 107878 60954
rect 107878 60902 107890 60954
rect 107890 60902 107904 60954
rect 107928 60902 107942 60954
rect 107942 60902 107954 60954
rect 107954 60902 107984 60954
rect 108008 60902 108018 60954
rect 108018 60902 108064 60954
rect 107768 60900 107824 60902
rect 107848 60900 107904 60902
rect 107928 60900 107984 60902
rect 108008 60900 108064 60902
rect 107032 60410 107088 60412
rect 107112 60410 107168 60412
rect 107192 60410 107248 60412
rect 107272 60410 107328 60412
rect 107032 60358 107078 60410
rect 107078 60358 107088 60410
rect 107112 60358 107142 60410
rect 107142 60358 107154 60410
rect 107154 60358 107168 60410
rect 107192 60358 107206 60410
rect 107206 60358 107218 60410
rect 107218 60358 107248 60410
rect 107272 60358 107282 60410
rect 107282 60358 107328 60410
rect 107032 60356 107088 60358
rect 107112 60356 107168 60358
rect 107192 60356 107248 60358
rect 107272 60356 107328 60358
rect 107768 59866 107824 59868
rect 107848 59866 107904 59868
rect 107928 59866 107984 59868
rect 108008 59866 108064 59868
rect 107768 59814 107814 59866
rect 107814 59814 107824 59866
rect 107848 59814 107878 59866
rect 107878 59814 107890 59866
rect 107890 59814 107904 59866
rect 107928 59814 107942 59866
rect 107942 59814 107954 59866
rect 107954 59814 107984 59866
rect 108008 59814 108018 59866
rect 108018 59814 108064 59866
rect 107768 59812 107824 59814
rect 107848 59812 107904 59814
rect 107928 59812 107984 59814
rect 108008 59812 108064 59814
rect 107032 59322 107088 59324
rect 107112 59322 107168 59324
rect 107192 59322 107248 59324
rect 107272 59322 107328 59324
rect 107032 59270 107078 59322
rect 107078 59270 107088 59322
rect 107112 59270 107142 59322
rect 107142 59270 107154 59322
rect 107154 59270 107168 59322
rect 107192 59270 107206 59322
rect 107206 59270 107218 59322
rect 107218 59270 107248 59322
rect 107272 59270 107282 59322
rect 107282 59270 107328 59322
rect 107032 59268 107088 59270
rect 107112 59268 107168 59270
rect 107192 59268 107248 59270
rect 107272 59268 107328 59270
rect 107768 58778 107824 58780
rect 107848 58778 107904 58780
rect 107928 58778 107984 58780
rect 108008 58778 108064 58780
rect 107768 58726 107814 58778
rect 107814 58726 107824 58778
rect 107848 58726 107878 58778
rect 107878 58726 107890 58778
rect 107890 58726 107904 58778
rect 107928 58726 107942 58778
rect 107942 58726 107954 58778
rect 107954 58726 107984 58778
rect 108008 58726 108018 58778
rect 108018 58726 108064 58778
rect 107768 58724 107824 58726
rect 107848 58724 107904 58726
rect 107928 58724 107984 58726
rect 108008 58724 108064 58726
rect 107032 58234 107088 58236
rect 107112 58234 107168 58236
rect 107192 58234 107248 58236
rect 107272 58234 107328 58236
rect 107032 58182 107078 58234
rect 107078 58182 107088 58234
rect 107112 58182 107142 58234
rect 107142 58182 107154 58234
rect 107154 58182 107168 58234
rect 107192 58182 107206 58234
rect 107206 58182 107218 58234
rect 107218 58182 107248 58234
rect 107272 58182 107282 58234
rect 107282 58182 107328 58234
rect 107032 58180 107088 58182
rect 107112 58180 107168 58182
rect 107192 58180 107248 58182
rect 107272 58180 107328 58182
rect 107768 57690 107824 57692
rect 107848 57690 107904 57692
rect 107928 57690 107984 57692
rect 108008 57690 108064 57692
rect 107768 57638 107814 57690
rect 107814 57638 107824 57690
rect 107848 57638 107878 57690
rect 107878 57638 107890 57690
rect 107890 57638 107904 57690
rect 107928 57638 107942 57690
rect 107942 57638 107954 57690
rect 107954 57638 107984 57690
rect 108008 57638 108018 57690
rect 108018 57638 108064 57690
rect 107768 57636 107824 57638
rect 107848 57636 107904 57638
rect 107928 57636 107984 57638
rect 108008 57636 108064 57638
rect 107032 57146 107088 57148
rect 107112 57146 107168 57148
rect 107192 57146 107248 57148
rect 107272 57146 107328 57148
rect 107032 57094 107078 57146
rect 107078 57094 107088 57146
rect 107112 57094 107142 57146
rect 107142 57094 107154 57146
rect 107154 57094 107168 57146
rect 107192 57094 107206 57146
rect 107206 57094 107218 57146
rect 107218 57094 107248 57146
rect 107272 57094 107282 57146
rect 107282 57094 107328 57146
rect 107032 57092 107088 57094
rect 107112 57092 107168 57094
rect 107192 57092 107248 57094
rect 107272 57092 107328 57094
rect 107768 56602 107824 56604
rect 107848 56602 107904 56604
rect 107928 56602 107984 56604
rect 108008 56602 108064 56604
rect 107768 56550 107814 56602
rect 107814 56550 107824 56602
rect 107848 56550 107878 56602
rect 107878 56550 107890 56602
rect 107890 56550 107904 56602
rect 107928 56550 107942 56602
rect 107942 56550 107954 56602
rect 107954 56550 107984 56602
rect 108008 56550 108018 56602
rect 108018 56550 108064 56602
rect 107768 56548 107824 56550
rect 107848 56548 107904 56550
rect 107928 56548 107984 56550
rect 108008 56548 108064 56550
rect 107032 56058 107088 56060
rect 107112 56058 107168 56060
rect 107192 56058 107248 56060
rect 107272 56058 107328 56060
rect 107032 56006 107078 56058
rect 107078 56006 107088 56058
rect 107112 56006 107142 56058
rect 107142 56006 107154 56058
rect 107154 56006 107168 56058
rect 107192 56006 107206 56058
rect 107206 56006 107218 56058
rect 107218 56006 107248 56058
rect 107272 56006 107282 56058
rect 107282 56006 107328 56058
rect 107032 56004 107088 56006
rect 107112 56004 107168 56006
rect 107192 56004 107248 56006
rect 107272 56004 107328 56006
rect 107768 55514 107824 55516
rect 107848 55514 107904 55516
rect 107928 55514 107984 55516
rect 108008 55514 108064 55516
rect 107768 55462 107814 55514
rect 107814 55462 107824 55514
rect 107848 55462 107878 55514
rect 107878 55462 107890 55514
rect 107890 55462 107904 55514
rect 107928 55462 107942 55514
rect 107942 55462 107954 55514
rect 107954 55462 107984 55514
rect 108008 55462 108018 55514
rect 108018 55462 108064 55514
rect 107768 55460 107824 55462
rect 107848 55460 107904 55462
rect 107928 55460 107984 55462
rect 108008 55460 108064 55462
rect 107032 54970 107088 54972
rect 107112 54970 107168 54972
rect 107192 54970 107248 54972
rect 107272 54970 107328 54972
rect 107032 54918 107078 54970
rect 107078 54918 107088 54970
rect 107112 54918 107142 54970
rect 107142 54918 107154 54970
rect 107154 54918 107168 54970
rect 107192 54918 107206 54970
rect 107206 54918 107218 54970
rect 107218 54918 107248 54970
rect 107272 54918 107282 54970
rect 107282 54918 107328 54970
rect 107032 54916 107088 54918
rect 107112 54916 107168 54918
rect 107192 54916 107248 54918
rect 107272 54916 107328 54918
rect 107768 54426 107824 54428
rect 107848 54426 107904 54428
rect 107928 54426 107984 54428
rect 108008 54426 108064 54428
rect 107768 54374 107814 54426
rect 107814 54374 107824 54426
rect 107848 54374 107878 54426
rect 107878 54374 107890 54426
rect 107890 54374 107904 54426
rect 107928 54374 107942 54426
rect 107942 54374 107954 54426
rect 107954 54374 107984 54426
rect 108008 54374 108018 54426
rect 108018 54374 108064 54426
rect 107768 54372 107824 54374
rect 107848 54372 107904 54374
rect 107928 54372 107984 54374
rect 108008 54372 108064 54374
rect 107032 53882 107088 53884
rect 107112 53882 107168 53884
rect 107192 53882 107248 53884
rect 107272 53882 107328 53884
rect 107032 53830 107078 53882
rect 107078 53830 107088 53882
rect 107112 53830 107142 53882
rect 107142 53830 107154 53882
rect 107154 53830 107168 53882
rect 107192 53830 107206 53882
rect 107206 53830 107218 53882
rect 107218 53830 107248 53882
rect 107272 53830 107282 53882
rect 107282 53830 107328 53882
rect 107032 53828 107088 53830
rect 107112 53828 107168 53830
rect 107192 53828 107248 53830
rect 107272 53828 107328 53830
rect 107768 53338 107824 53340
rect 107848 53338 107904 53340
rect 107928 53338 107984 53340
rect 108008 53338 108064 53340
rect 107768 53286 107814 53338
rect 107814 53286 107824 53338
rect 107848 53286 107878 53338
rect 107878 53286 107890 53338
rect 107890 53286 107904 53338
rect 107928 53286 107942 53338
rect 107942 53286 107954 53338
rect 107954 53286 107984 53338
rect 108008 53286 108018 53338
rect 108018 53286 108064 53338
rect 107768 53284 107824 53286
rect 107848 53284 107904 53286
rect 107928 53284 107984 53286
rect 108008 53284 108064 53286
rect 107032 52794 107088 52796
rect 107112 52794 107168 52796
rect 107192 52794 107248 52796
rect 107272 52794 107328 52796
rect 107032 52742 107078 52794
rect 107078 52742 107088 52794
rect 107112 52742 107142 52794
rect 107142 52742 107154 52794
rect 107154 52742 107168 52794
rect 107192 52742 107206 52794
rect 107206 52742 107218 52794
rect 107218 52742 107248 52794
rect 107272 52742 107282 52794
rect 107282 52742 107328 52794
rect 107032 52740 107088 52742
rect 107112 52740 107168 52742
rect 107192 52740 107248 52742
rect 107272 52740 107328 52742
rect 107768 52250 107824 52252
rect 107848 52250 107904 52252
rect 107928 52250 107984 52252
rect 108008 52250 108064 52252
rect 107768 52198 107814 52250
rect 107814 52198 107824 52250
rect 107848 52198 107878 52250
rect 107878 52198 107890 52250
rect 107890 52198 107904 52250
rect 107928 52198 107942 52250
rect 107942 52198 107954 52250
rect 107954 52198 107984 52250
rect 108008 52198 108018 52250
rect 108018 52198 108064 52250
rect 107768 52196 107824 52198
rect 107848 52196 107904 52198
rect 107928 52196 107984 52198
rect 108008 52196 108064 52198
rect 107032 51706 107088 51708
rect 107112 51706 107168 51708
rect 107192 51706 107248 51708
rect 107272 51706 107328 51708
rect 107032 51654 107078 51706
rect 107078 51654 107088 51706
rect 107112 51654 107142 51706
rect 107142 51654 107154 51706
rect 107154 51654 107168 51706
rect 107192 51654 107206 51706
rect 107206 51654 107218 51706
rect 107218 51654 107248 51706
rect 107272 51654 107282 51706
rect 107282 51654 107328 51706
rect 107032 51652 107088 51654
rect 107112 51652 107168 51654
rect 107192 51652 107248 51654
rect 107272 51652 107328 51654
rect 107768 51162 107824 51164
rect 107848 51162 107904 51164
rect 107928 51162 107984 51164
rect 108008 51162 108064 51164
rect 107768 51110 107814 51162
rect 107814 51110 107824 51162
rect 107848 51110 107878 51162
rect 107878 51110 107890 51162
rect 107890 51110 107904 51162
rect 107928 51110 107942 51162
rect 107942 51110 107954 51162
rect 107954 51110 107984 51162
rect 108008 51110 108018 51162
rect 108018 51110 108064 51162
rect 107768 51108 107824 51110
rect 107848 51108 107904 51110
rect 107928 51108 107984 51110
rect 108008 51108 108064 51110
rect 107032 50618 107088 50620
rect 107112 50618 107168 50620
rect 107192 50618 107248 50620
rect 107272 50618 107328 50620
rect 107032 50566 107078 50618
rect 107078 50566 107088 50618
rect 107112 50566 107142 50618
rect 107142 50566 107154 50618
rect 107154 50566 107168 50618
rect 107192 50566 107206 50618
rect 107206 50566 107218 50618
rect 107218 50566 107248 50618
rect 107272 50566 107282 50618
rect 107282 50566 107328 50618
rect 107032 50564 107088 50566
rect 107112 50564 107168 50566
rect 107192 50564 107248 50566
rect 107272 50564 107328 50566
rect 107768 50074 107824 50076
rect 107848 50074 107904 50076
rect 107928 50074 107984 50076
rect 108008 50074 108064 50076
rect 107768 50022 107814 50074
rect 107814 50022 107824 50074
rect 107848 50022 107878 50074
rect 107878 50022 107890 50074
rect 107890 50022 107904 50074
rect 107928 50022 107942 50074
rect 107942 50022 107954 50074
rect 107954 50022 107984 50074
rect 108008 50022 108018 50074
rect 108018 50022 108064 50074
rect 107768 50020 107824 50022
rect 107848 50020 107904 50022
rect 107928 50020 107984 50022
rect 108008 50020 108064 50022
rect 107032 49530 107088 49532
rect 107112 49530 107168 49532
rect 107192 49530 107248 49532
rect 107272 49530 107328 49532
rect 107032 49478 107078 49530
rect 107078 49478 107088 49530
rect 107112 49478 107142 49530
rect 107142 49478 107154 49530
rect 107154 49478 107168 49530
rect 107192 49478 107206 49530
rect 107206 49478 107218 49530
rect 107218 49478 107248 49530
rect 107272 49478 107282 49530
rect 107282 49478 107328 49530
rect 107032 49476 107088 49478
rect 107112 49476 107168 49478
rect 107192 49476 107248 49478
rect 107272 49476 107328 49478
rect 107768 48986 107824 48988
rect 107848 48986 107904 48988
rect 107928 48986 107984 48988
rect 108008 48986 108064 48988
rect 107768 48934 107814 48986
rect 107814 48934 107824 48986
rect 107848 48934 107878 48986
rect 107878 48934 107890 48986
rect 107890 48934 107904 48986
rect 107928 48934 107942 48986
rect 107942 48934 107954 48986
rect 107954 48934 107984 48986
rect 108008 48934 108018 48986
rect 108018 48934 108064 48986
rect 107768 48932 107824 48934
rect 107848 48932 107904 48934
rect 107928 48932 107984 48934
rect 108008 48932 108064 48934
rect 107032 48442 107088 48444
rect 107112 48442 107168 48444
rect 107192 48442 107248 48444
rect 107272 48442 107328 48444
rect 107032 48390 107078 48442
rect 107078 48390 107088 48442
rect 107112 48390 107142 48442
rect 107142 48390 107154 48442
rect 107154 48390 107168 48442
rect 107192 48390 107206 48442
rect 107206 48390 107218 48442
rect 107218 48390 107248 48442
rect 107272 48390 107282 48442
rect 107282 48390 107328 48442
rect 107032 48388 107088 48390
rect 107112 48388 107168 48390
rect 107192 48388 107248 48390
rect 107272 48388 107328 48390
rect 107768 47898 107824 47900
rect 107848 47898 107904 47900
rect 107928 47898 107984 47900
rect 108008 47898 108064 47900
rect 107768 47846 107814 47898
rect 107814 47846 107824 47898
rect 107848 47846 107878 47898
rect 107878 47846 107890 47898
rect 107890 47846 107904 47898
rect 107928 47846 107942 47898
rect 107942 47846 107954 47898
rect 107954 47846 107984 47898
rect 108008 47846 108018 47898
rect 108018 47846 108064 47898
rect 107768 47844 107824 47846
rect 107848 47844 107904 47846
rect 107928 47844 107984 47846
rect 108008 47844 108064 47846
rect 107032 47354 107088 47356
rect 107112 47354 107168 47356
rect 107192 47354 107248 47356
rect 107272 47354 107328 47356
rect 107032 47302 107078 47354
rect 107078 47302 107088 47354
rect 107112 47302 107142 47354
rect 107142 47302 107154 47354
rect 107154 47302 107168 47354
rect 107192 47302 107206 47354
rect 107206 47302 107218 47354
rect 107218 47302 107248 47354
rect 107272 47302 107282 47354
rect 107282 47302 107328 47354
rect 107032 47300 107088 47302
rect 107112 47300 107168 47302
rect 107192 47300 107248 47302
rect 107272 47300 107328 47302
rect 107768 46810 107824 46812
rect 107848 46810 107904 46812
rect 107928 46810 107984 46812
rect 108008 46810 108064 46812
rect 107768 46758 107814 46810
rect 107814 46758 107824 46810
rect 107848 46758 107878 46810
rect 107878 46758 107890 46810
rect 107890 46758 107904 46810
rect 107928 46758 107942 46810
rect 107942 46758 107954 46810
rect 107954 46758 107984 46810
rect 108008 46758 108018 46810
rect 108018 46758 108064 46810
rect 107768 46756 107824 46758
rect 107848 46756 107904 46758
rect 107928 46756 107984 46758
rect 108008 46756 108064 46758
rect 107032 46266 107088 46268
rect 107112 46266 107168 46268
rect 107192 46266 107248 46268
rect 107272 46266 107328 46268
rect 107032 46214 107078 46266
rect 107078 46214 107088 46266
rect 107112 46214 107142 46266
rect 107142 46214 107154 46266
rect 107154 46214 107168 46266
rect 107192 46214 107206 46266
rect 107206 46214 107218 46266
rect 107218 46214 107248 46266
rect 107272 46214 107282 46266
rect 107282 46214 107328 46266
rect 107032 46212 107088 46214
rect 107112 46212 107168 46214
rect 107192 46212 107248 46214
rect 107272 46212 107328 46214
rect 107768 45722 107824 45724
rect 107848 45722 107904 45724
rect 107928 45722 107984 45724
rect 108008 45722 108064 45724
rect 107768 45670 107814 45722
rect 107814 45670 107824 45722
rect 107848 45670 107878 45722
rect 107878 45670 107890 45722
rect 107890 45670 107904 45722
rect 107928 45670 107942 45722
rect 107942 45670 107954 45722
rect 107954 45670 107984 45722
rect 108008 45670 108018 45722
rect 108018 45670 108064 45722
rect 107768 45668 107824 45670
rect 107848 45668 107904 45670
rect 107928 45668 107984 45670
rect 108008 45668 108064 45670
rect 107032 45178 107088 45180
rect 107112 45178 107168 45180
rect 107192 45178 107248 45180
rect 107272 45178 107328 45180
rect 107032 45126 107078 45178
rect 107078 45126 107088 45178
rect 107112 45126 107142 45178
rect 107142 45126 107154 45178
rect 107154 45126 107168 45178
rect 107192 45126 107206 45178
rect 107206 45126 107218 45178
rect 107218 45126 107248 45178
rect 107272 45126 107282 45178
rect 107282 45126 107328 45178
rect 107032 45124 107088 45126
rect 107112 45124 107168 45126
rect 107192 45124 107248 45126
rect 107272 45124 107328 45126
rect 107768 44634 107824 44636
rect 107848 44634 107904 44636
rect 107928 44634 107984 44636
rect 108008 44634 108064 44636
rect 107768 44582 107814 44634
rect 107814 44582 107824 44634
rect 107848 44582 107878 44634
rect 107878 44582 107890 44634
rect 107890 44582 107904 44634
rect 107928 44582 107942 44634
rect 107942 44582 107954 44634
rect 107954 44582 107984 44634
rect 108008 44582 108018 44634
rect 108018 44582 108064 44634
rect 107768 44580 107824 44582
rect 107848 44580 107904 44582
rect 107928 44580 107984 44582
rect 108008 44580 108064 44582
rect 107032 44090 107088 44092
rect 107112 44090 107168 44092
rect 107192 44090 107248 44092
rect 107272 44090 107328 44092
rect 107032 44038 107078 44090
rect 107078 44038 107088 44090
rect 107112 44038 107142 44090
rect 107142 44038 107154 44090
rect 107154 44038 107168 44090
rect 107192 44038 107206 44090
rect 107206 44038 107218 44090
rect 107218 44038 107248 44090
rect 107272 44038 107282 44090
rect 107282 44038 107328 44090
rect 107032 44036 107088 44038
rect 107112 44036 107168 44038
rect 107192 44036 107248 44038
rect 107272 44036 107328 44038
rect 107768 43546 107824 43548
rect 107848 43546 107904 43548
rect 107928 43546 107984 43548
rect 108008 43546 108064 43548
rect 107768 43494 107814 43546
rect 107814 43494 107824 43546
rect 107848 43494 107878 43546
rect 107878 43494 107890 43546
rect 107890 43494 107904 43546
rect 107928 43494 107942 43546
rect 107942 43494 107954 43546
rect 107954 43494 107984 43546
rect 108008 43494 108018 43546
rect 108018 43494 108064 43546
rect 107768 43492 107824 43494
rect 107848 43492 107904 43494
rect 107928 43492 107984 43494
rect 108008 43492 108064 43494
rect 107032 43002 107088 43004
rect 107112 43002 107168 43004
rect 107192 43002 107248 43004
rect 107272 43002 107328 43004
rect 107032 42950 107078 43002
rect 107078 42950 107088 43002
rect 107112 42950 107142 43002
rect 107142 42950 107154 43002
rect 107154 42950 107168 43002
rect 107192 42950 107206 43002
rect 107206 42950 107218 43002
rect 107218 42950 107248 43002
rect 107272 42950 107282 43002
rect 107282 42950 107328 43002
rect 107032 42948 107088 42950
rect 107112 42948 107168 42950
rect 107192 42948 107248 42950
rect 107272 42948 107328 42950
rect 107768 42458 107824 42460
rect 107848 42458 107904 42460
rect 107928 42458 107984 42460
rect 108008 42458 108064 42460
rect 107768 42406 107814 42458
rect 107814 42406 107824 42458
rect 107848 42406 107878 42458
rect 107878 42406 107890 42458
rect 107890 42406 107904 42458
rect 107928 42406 107942 42458
rect 107942 42406 107954 42458
rect 107954 42406 107984 42458
rect 108008 42406 108018 42458
rect 108018 42406 108064 42458
rect 107768 42404 107824 42406
rect 107848 42404 107904 42406
rect 107928 42404 107984 42406
rect 108008 42404 108064 42406
rect 107032 41914 107088 41916
rect 107112 41914 107168 41916
rect 107192 41914 107248 41916
rect 107272 41914 107328 41916
rect 107032 41862 107078 41914
rect 107078 41862 107088 41914
rect 107112 41862 107142 41914
rect 107142 41862 107154 41914
rect 107154 41862 107168 41914
rect 107192 41862 107206 41914
rect 107206 41862 107218 41914
rect 107218 41862 107248 41914
rect 107272 41862 107282 41914
rect 107282 41862 107328 41914
rect 107032 41860 107088 41862
rect 107112 41860 107168 41862
rect 107192 41860 107248 41862
rect 107272 41860 107328 41862
rect 107768 41370 107824 41372
rect 107848 41370 107904 41372
rect 107928 41370 107984 41372
rect 108008 41370 108064 41372
rect 107768 41318 107814 41370
rect 107814 41318 107824 41370
rect 107848 41318 107878 41370
rect 107878 41318 107890 41370
rect 107890 41318 107904 41370
rect 107928 41318 107942 41370
rect 107942 41318 107954 41370
rect 107954 41318 107984 41370
rect 108008 41318 108018 41370
rect 108018 41318 108064 41370
rect 107768 41316 107824 41318
rect 107848 41316 107904 41318
rect 107928 41316 107984 41318
rect 108008 41316 108064 41318
rect 107032 40826 107088 40828
rect 107112 40826 107168 40828
rect 107192 40826 107248 40828
rect 107272 40826 107328 40828
rect 107032 40774 107078 40826
rect 107078 40774 107088 40826
rect 107112 40774 107142 40826
rect 107142 40774 107154 40826
rect 107154 40774 107168 40826
rect 107192 40774 107206 40826
rect 107206 40774 107218 40826
rect 107218 40774 107248 40826
rect 107272 40774 107282 40826
rect 107282 40774 107328 40826
rect 107032 40772 107088 40774
rect 107112 40772 107168 40774
rect 107192 40772 107248 40774
rect 107272 40772 107328 40774
rect 107768 40282 107824 40284
rect 107848 40282 107904 40284
rect 107928 40282 107984 40284
rect 108008 40282 108064 40284
rect 107768 40230 107814 40282
rect 107814 40230 107824 40282
rect 107848 40230 107878 40282
rect 107878 40230 107890 40282
rect 107890 40230 107904 40282
rect 107928 40230 107942 40282
rect 107942 40230 107954 40282
rect 107954 40230 107984 40282
rect 108008 40230 108018 40282
rect 108018 40230 108064 40282
rect 107768 40228 107824 40230
rect 107848 40228 107904 40230
rect 107928 40228 107984 40230
rect 108008 40228 108064 40230
rect 107032 39738 107088 39740
rect 107112 39738 107168 39740
rect 107192 39738 107248 39740
rect 107272 39738 107328 39740
rect 107032 39686 107078 39738
rect 107078 39686 107088 39738
rect 107112 39686 107142 39738
rect 107142 39686 107154 39738
rect 107154 39686 107168 39738
rect 107192 39686 107206 39738
rect 107206 39686 107218 39738
rect 107218 39686 107248 39738
rect 107272 39686 107282 39738
rect 107282 39686 107328 39738
rect 107032 39684 107088 39686
rect 107112 39684 107168 39686
rect 107192 39684 107248 39686
rect 107272 39684 107328 39686
rect 107768 39194 107824 39196
rect 107848 39194 107904 39196
rect 107928 39194 107984 39196
rect 108008 39194 108064 39196
rect 107768 39142 107814 39194
rect 107814 39142 107824 39194
rect 107848 39142 107878 39194
rect 107878 39142 107890 39194
rect 107890 39142 107904 39194
rect 107928 39142 107942 39194
rect 107942 39142 107954 39194
rect 107954 39142 107984 39194
rect 108008 39142 108018 39194
rect 108018 39142 108064 39194
rect 107768 39140 107824 39142
rect 107848 39140 107904 39142
rect 107928 39140 107984 39142
rect 108008 39140 108064 39142
rect 107032 38650 107088 38652
rect 107112 38650 107168 38652
rect 107192 38650 107248 38652
rect 107272 38650 107328 38652
rect 107032 38598 107078 38650
rect 107078 38598 107088 38650
rect 107112 38598 107142 38650
rect 107142 38598 107154 38650
rect 107154 38598 107168 38650
rect 107192 38598 107206 38650
rect 107206 38598 107218 38650
rect 107218 38598 107248 38650
rect 107272 38598 107282 38650
rect 107282 38598 107328 38650
rect 107032 38596 107088 38598
rect 107112 38596 107168 38598
rect 107192 38596 107248 38598
rect 107272 38596 107328 38598
rect 107768 38106 107824 38108
rect 107848 38106 107904 38108
rect 107928 38106 107984 38108
rect 108008 38106 108064 38108
rect 107768 38054 107814 38106
rect 107814 38054 107824 38106
rect 107848 38054 107878 38106
rect 107878 38054 107890 38106
rect 107890 38054 107904 38106
rect 107928 38054 107942 38106
rect 107942 38054 107954 38106
rect 107954 38054 107984 38106
rect 108008 38054 108018 38106
rect 108018 38054 108064 38106
rect 107768 38052 107824 38054
rect 107848 38052 107904 38054
rect 107928 38052 107984 38054
rect 108008 38052 108064 38054
rect 107032 37562 107088 37564
rect 107112 37562 107168 37564
rect 107192 37562 107248 37564
rect 107272 37562 107328 37564
rect 107032 37510 107078 37562
rect 107078 37510 107088 37562
rect 107112 37510 107142 37562
rect 107142 37510 107154 37562
rect 107154 37510 107168 37562
rect 107192 37510 107206 37562
rect 107206 37510 107218 37562
rect 107218 37510 107248 37562
rect 107272 37510 107282 37562
rect 107282 37510 107328 37562
rect 107032 37508 107088 37510
rect 107112 37508 107168 37510
rect 107192 37508 107248 37510
rect 107272 37508 107328 37510
rect 107768 37018 107824 37020
rect 107848 37018 107904 37020
rect 107928 37018 107984 37020
rect 108008 37018 108064 37020
rect 107768 36966 107814 37018
rect 107814 36966 107824 37018
rect 107848 36966 107878 37018
rect 107878 36966 107890 37018
rect 107890 36966 107904 37018
rect 107928 36966 107942 37018
rect 107942 36966 107954 37018
rect 107954 36966 107984 37018
rect 108008 36966 108018 37018
rect 108018 36966 108064 37018
rect 107768 36964 107824 36966
rect 107848 36964 107904 36966
rect 107928 36964 107984 36966
rect 108008 36964 108064 36966
rect 107032 36474 107088 36476
rect 107112 36474 107168 36476
rect 107192 36474 107248 36476
rect 107272 36474 107328 36476
rect 107032 36422 107078 36474
rect 107078 36422 107088 36474
rect 107112 36422 107142 36474
rect 107142 36422 107154 36474
rect 107154 36422 107168 36474
rect 107192 36422 107206 36474
rect 107206 36422 107218 36474
rect 107218 36422 107248 36474
rect 107272 36422 107282 36474
rect 107282 36422 107328 36474
rect 107032 36420 107088 36422
rect 107112 36420 107168 36422
rect 107192 36420 107248 36422
rect 107272 36420 107328 36422
rect 107768 35930 107824 35932
rect 107848 35930 107904 35932
rect 107928 35930 107984 35932
rect 108008 35930 108064 35932
rect 107768 35878 107814 35930
rect 107814 35878 107824 35930
rect 107848 35878 107878 35930
rect 107878 35878 107890 35930
rect 107890 35878 107904 35930
rect 107928 35878 107942 35930
rect 107942 35878 107954 35930
rect 107954 35878 107984 35930
rect 108008 35878 108018 35930
rect 108018 35878 108064 35930
rect 107768 35876 107824 35878
rect 107848 35876 107904 35878
rect 107928 35876 107984 35878
rect 108008 35876 108064 35878
rect 107032 35386 107088 35388
rect 107112 35386 107168 35388
rect 107192 35386 107248 35388
rect 107272 35386 107328 35388
rect 107032 35334 107078 35386
rect 107078 35334 107088 35386
rect 107112 35334 107142 35386
rect 107142 35334 107154 35386
rect 107154 35334 107168 35386
rect 107192 35334 107206 35386
rect 107206 35334 107218 35386
rect 107218 35334 107248 35386
rect 107272 35334 107282 35386
rect 107282 35334 107328 35386
rect 107032 35332 107088 35334
rect 107112 35332 107168 35334
rect 107192 35332 107248 35334
rect 107272 35332 107328 35334
rect 107768 34842 107824 34844
rect 107848 34842 107904 34844
rect 107928 34842 107984 34844
rect 108008 34842 108064 34844
rect 107768 34790 107814 34842
rect 107814 34790 107824 34842
rect 107848 34790 107878 34842
rect 107878 34790 107890 34842
rect 107890 34790 107904 34842
rect 107928 34790 107942 34842
rect 107942 34790 107954 34842
rect 107954 34790 107984 34842
rect 108008 34790 108018 34842
rect 108018 34790 108064 34842
rect 107768 34788 107824 34790
rect 107848 34788 107904 34790
rect 107928 34788 107984 34790
rect 108008 34788 108064 34790
rect 107032 34298 107088 34300
rect 107112 34298 107168 34300
rect 107192 34298 107248 34300
rect 107272 34298 107328 34300
rect 107032 34246 107078 34298
rect 107078 34246 107088 34298
rect 107112 34246 107142 34298
rect 107142 34246 107154 34298
rect 107154 34246 107168 34298
rect 107192 34246 107206 34298
rect 107206 34246 107218 34298
rect 107218 34246 107248 34298
rect 107272 34246 107282 34298
rect 107282 34246 107328 34298
rect 107032 34244 107088 34246
rect 107112 34244 107168 34246
rect 107192 34244 107248 34246
rect 107272 34244 107328 34246
rect 107768 33754 107824 33756
rect 107848 33754 107904 33756
rect 107928 33754 107984 33756
rect 108008 33754 108064 33756
rect 107768 33702 107814 33754
rect 107814 33702 107824 33754
rect 107848 33702 107878 33754
rect 107878 33702 107890 33754
rect 107890 33702 107904 33754
rect 107928 33702 107942 33754
rect 107942 33702 107954 33754
rect 107954 33702 107984 33754
rect 108008 33702 108018 33754
rect 108018 33702 108064 33754
rect 107768 33700 107824 33702
rect 107848 33700 107904 33702
rect 107928 33700 107984 33702
rect 108008 33700 108064 33702
rect 107032 33210 107088 33212
rect 107112 33210 107168 33212
rect 107192 33210 107248 33212
rect 107272 33210 107328 33212
rect 107032 33158 107078 33210
rect 107078 33158 107088 33210
rect 107112 33158 107142 33210
rect 107142 33158 107154 33210
rect 107154 33158 107168 33210
rect 107192 33158 107206 33210
rect 107206 33158 107218 33210
rect 107218 33158 107248 33210
rect 107272 33158 107282 33210
rect 107282 33158 107328 33210
rect 107032 33156 107088 33158
rect 107112 33156 107168 33158
rect 107192 33156 107248 33158
rect 107272 33156 107328 33158
rect 104162 25064 104218 25120
rect 104346 23296 104402 23352
rect 16026 9832 16082 9888
rect 90362 9832 90418 9888
rect 31574 9696 31630 9752
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 23478 9560 23534 9616
rect 30470 9560 30526 9616
rect 25778 8064 25834 8120
rect 28998 8064 29054 8120
rect 24674 7540 24730 7576
rect 24674 7520 24676 7540
rect 24676 7520 24728 7540
rect 24728 7520 24730 7540
rect 26974 7540 27030 7576
rect 26974 7520 26976 7540
rect 26976 7520 27028 7540
rect 27028 7520 27030 7540
rect 28262 7540 28318 7576
rect 107768 32666 107824 32668
rect 107848 32666 107904 32668
rect 107928 32666 107984 32668
rect 108008 32666 108064 32668
rect 107768 32614 107814 32666
rect 107814 32614 107824 32666
rect 107848 32614 107878 32666
rect 107878 32614 107890 32666
rect 107890 32614 107904 32666
rect 107928 32614 107942 32666
rect 107942 32614 107954 32666
rect 107954 32614 107984 32666
rect 108008 32614 108018 32666
rect 108018 32614 108064 32666
rect 107768 32612 107824 32614
rect 107848 32612 107904 32614
rect 107928 32612 107984 32614
rect 108008 32612 108064 32614
rect 107032 32122 107088 32124
rect 107112 32122 107168 32124
rect 107192 32122 107248 32124
rect 107272 32122 107328 32124
rect 107032 32070 107078 32122
rect 107078 32070 107088 32122
rect 107112 32070 107142 32122
rect 107142 32070 107154 32122
rect 107154 32070 107168 32122
rect 107192 32070 107206 32122
rect 107206 32070 107218 32122
rect 107218 32070 107248 32122
rect 107272 32070 107282 32122
rect 107282 32070 107328 32122
rect 107032 32068 107088 32070
rect 107112 32068 107168 32070
rect 107192 32068 107248 32070
rect 107272 32068 107328 32070
rect 107768 31578 107824 31580
rect 107848 31578 107904 31580
rect 107928 31578 107984 31580
rect 108008 31578 108064 31580
rect 107768 31526 107814 31578
rect 107814 31526 107824 31578
rect 107848 31526 107878 31578
rect 107878 31526 107890 31578
rect 107890 31526 107904 31578
rect 107928 31526 107942 31578
rect 107942 31526 107954 31578
rect 107954 31526 107984 31578
rect 108008 31526 108018 31578
rect 108018 31526 108064 31578
rect 107768 31524 107824 31526
rect 107848 31524 107904 31526
rect 107928 31524 107984 31526
rect 108008 31524 108064 31526
rect 110510 31320 110566 31376
rect 107032 31034 107088 31036
rect 107112 31034 107168 31036
rect 107192 31034 107248 31036
rect 107272 31034 107328 31036
rect 107032 30982 107078 31034
rect 107078 30982 107088 31034
rect 107112 30982 107142 31034
rect 107142 30982 107154 31034
rect 107154 30982 107168 31034
rect 107192 30982 107206 31034
rect 107206 30982 107218 31034
rect 107218 30982 107248 31034
rect 107272 30982 107282 31034
rect 107282 30982 107328 31034
rect 107032 30980 107088 30982
rect 107112 30980 107168 30982
rect 107192 30980 107248 30982
rect 107272 30980 107328 30982
rect 107768 30490 107824 30492
rect 107848 30490 107904 30492
rect 107928 30490 107984 30492
rect 108008 30490 108064 30492
rect 107768 30438 107814 30490
rect 107814 30438 107824 30490
rect 107848 30438 107878 30490
rect 107878 30438 107890 30490
rect 107890 30438 107904 30490
rect 107928 30438 107942 30490
rect 107942 30438 107954 30490
rect 107954 30438 107984 30490
rect 108008 30438 108018 30490
rect 108018 30438 108064 30490
rect 107768 30436 107824 30438
rect 107848 30436 107904 30438
rect 107928 30436 107984 30438
rect 108008 30436 108064 30438
rect 107032 29946 107088 29948
rect 107112 29946 107168 29948
rect 107192 29946 107248 29948
rect 107272 29946 107328 29948
rect 107032 29894 107078 29946
rect 107078 29894 107088 29946
rect 107112 29894 107142 29946
rect 107142 29894 107154 29946
rect 107154 29894 107168 29946
rect 107192 29894 107206 29946
rect 107206 29894 107218 29946
rect 107218 29894 107248 29946
rect 107272 29894 107282 29946
rect 107282 29894 107328 29946
rect 107032 29892 107088 29894
rect 107112 29892 107168 29894
rect 107192 29892 107248 29894
rect 107272 29892 107328 29894
rect 107768 29402 107824 29404
rect 107848 29402 107904 29404
rect 107928 29402 107984 29404
rect 108008 29402 108064 29404
rect 107768 29350 107814 29402
rect 107814 29350 107824 29402
rect 107848 29350 107878 29402
rect 107878 29350 107890 29402
rect 107890 29350 107904 29402
rect 107928 29350 107942 29402
rect 107942 29350 107954 29402
rect 107954 29350 107984 29402
rect 108008 29350 108018 29402
rect 108018 29350 108064 29402
rect 107768 29348 107824 29350
rect 107848 29348 107904 29350
rect 107928 29348 107984 29350
rect 108008 29348 108064 29350
rect 107032 28858 107088 28860
rect 107112 28858 107168 28860
rect 107192 28858 107248 28860
rect 107272 28858 107328 28860
rect 107032 28806 107078 28858
rect 107078 28806 107088 28858
rect 107112 28806 107142 28858
rect 107142 28806 107154 28858
rect 107154 28806 107168 28858
rect 107192 28806 107206 28858
rect 107206 28806 107218 28858
rect 107218 28806 107248 28858
rect 107272 28806 107282 28858
rect 107282 28806 107328 28858
rect 107032 28804 107088 28806
rect 107112 28804 107168 28806
rect 107192 28804 107248 28806
rect 107272 28804 107328 28806
rect 107768 28314 107824 28316
rect 107848 28314 107904 28316
rect 107928 28314 107984 28316
rect 108008 28314 108064 28316
rect 107768 28262 107814 28314
rect 107814 28262 107824 28314
rect 107848 28262 107878 28314
rect 107878 28262 107890 28314
rect 107890 28262 107904 28314
rect 107928 28262 107942 28314
rect 107942 28262 107954 28314
rect 107954 28262 107984 28314
rect 108008 28262 108018 28314
rect 108018 28262 108064 28314
rect 107768 28260 107824 28262
rect 107848 28260 107904 28262
rect 107928 28260 107984 28262
rect 108008 28260 108064 28262
rect 107032 27770 107088 27772
rect 107112 27770 107168 27772
rect 107192 27770 107248 27772
rect 107272 27770 107328 27772
rect 107032 27718 107078 27770
rect 107078 27718 107088 27770
rect 107112 27718 107142 27770
rect 107142 27718 107154 27770
rect 107154 27718 107168 27770
rect 107192 27718 107206 27770
rect 107206 27718 107218 27770
rect 107218 27718 107248 27770
rect 107272 27718 107282 27770
rect 107282 27718 107328 27770
rect 107032 27716 107088 27718
rect 107112 27716 107168 27718
rect 107192 27716 107248 27718
rect 107272 27716 107328 27718
rect 107768 27226 107824 27228
rect 107848 27226 107904 27228
rect 107928 27226 107984 27228
rect 108008 27226 108064 27228
rect 107768 27174 107814 27226
rect 107814 27174 107824 27226
rect 107848 27174 107878 27226
rect 107878 27174 107890 27226
rect 107890 27174 107904 27226
rect 107928 27174 107942 27226
rect 107942 27174 107954 27226
rect 107954 27174 107984 27226
rect 108008 27174 108018 27226
rect 108018 27174 108064 27226
rect 107768 27172 107824 27174
rect 107848 27172 107904 27174
rect 107928 27172 107984 27174
rect 108008 27172 108064 27174
rect 107032 26682 107088 26684
rect 107112 26682 107168 26684
rect 107192 26682 107248 26684
rect 107272 26682 107328 26684
rect 107032 26630 107078 26682
rect 107078 26630 107088 26682
rect 107112 26630 107142 26682
rect 107142 26630 107154 26682
rect 107154 26630 107168 26682
rect 107192 26630 107206 26682
rect 107206 26630 107218 26682
rect 107218 26630 107248 26682
rect 107272 26630 107282 26682
rect 107282 26630 107328 26682
rect 107032 26628 107088 26630
rect 107112 26628 107168 26630
rect 107192 26628 107248 26630
rect 107272 26628 107328 26630
rect 104530 22208 104586 22264
rect 107768 26138 107824 26140
rect 107848 26138 107904 26140
rect 107928 26138 107984 26140
rect 108008 26138 108064 26140
rect 107768 26086 107814 26138
rect 107814 26086 107824 26138
rect 107848 26086 107878 26138
rect 107878 26086 107890 26138
rect 107890 26086 107904 26138
rect 107928 26086 107942 26138
rect 107942 26086 107954 26138
rect 107954 26086 107984 26138
rect 108008 26086 108018 26138
rect 108018 26086 108064 26138
rect 107768 26084 107824 26086
rect 107848 26084 107904 26086
rect 107928 26084 107984 26086
rect 108008 26084 108064 26086
rect 107032 25594 107088 25596
rect 107112 25594 107168 25596
rect 107192 25594 107248 25596
rect 107272 25594 107328 25596
rect 107032 25542 107078 25594
rect 107078 25542 107088 25594
rect 107112 25542 107142 25594
rect 107142 25542 107154 25594
rect 107154 25542 107168 25594
rect 107192 25542 107206 25594
rect 107206 25542 107218 25594
rect 107218 25542 107248 25594
rect 107272 25542 107282 25594
rect 107282 25542 107328 25594
rect 107032 25540 107088 25542
rect 107112 25540 107168 25542
rect 107192 25540 107248 25542
rect 107272 25540 107328 25542
rect 107768 25050 107824 25052
rect 107848 25050 107904 25052
rect 107928 25050 107984 25052
rect 108008 25050 108064 25052
rect 107768 24998 107814 25050
rect 107814 24998 107824 25050
rect 107848 24998 107878 25050
rect 107878 24998 107890 25050
rect 107890 24998 107904 25050
rect 107928 24998 107942 25050
rect 107942 24998 107954 25050
rect 107954 24998 107984 25050
rect 108008 24998 108018 25050
rect 108018 24998 108064 25050
rect 107768 24996 107824 24998
rect 107848 24996 107904 24998
rect 107928 24996 107984 24998
rect 108008 24996 108064 24998
rect 107032 24506 107088 24508
rect 107112 24506 107168 24508
rect 107192 24506 107248 24508
rect 107272 24506 107328 24508
rect 107032 24454 107078 24506
rect 107078 24454 107088 24506
rect 107112 24454 107142 24506
rect 107142 24454 107154 24506
rect 107154 24454 107168 24506
rect 107192 24454 107206 24506
rect 107206 24454 107218 24506
rect 107218 24454 107248 24506
rect 107272 24454 107282 24506
rect 107282 24454 107328 24506
rect 107032 24452 107088 24454
rect 107112 24452 107168 24454
rect 107192 24452 107248 24454
rect 107272 24452 107328 24454
rect 107768 23962 107824 23964
rect 107848 23962 107904 23964
rect 107928 23962 107984 23964
rect 108008 23962 108064 23964
rect 107768 23910 107814 23962
rect 107814 23910 107824 23962
rect 107848 23910 107878 23962
rect 107878 23910 107890 23962
rect 107890 23910 107904 23962
rect 107928 23910 107942 23962
rect 107942 23910 107954 23962
rect 107954 23910 107984 23962
rect 108008 23910 108018 23962
rect 108018 23910 108064 23962
rect 107768 23908 107824 23910
rect 107848 23908 107904 23910
rect 107928 23908 107984 23910
rect 108008 23908 108064 23910
rect 107032 23418 107088 23420
rect 107112 23418 107168 23420
rect 107192 23418 107248 23420
rect 107272 23418 107328 23420
rect 107032 23366 107078 23418
rect 107078 23366 107088 23418
rect 107112 23366 107142 23418
rect 107142 23366 107154 23418
rect 107154 23366 107168 23418
rect 107192 23366 107206 23418
rect 107206 23366 107218 23418
rect 107218 23366 107248 23418
rect 107272 23366 107282 23418
rect 107282 23366 107328 23418
rect 107032 23364 107088 23366
rect 107112 23364 107168 23366
rect 107192 23364 107248 23366
rect 107272 23364 107328 23366
rect 107768 22874 107824 22876
rect 107848 22874 107904 22876
rect 107928 22874 107984 22876
rect 108008 22874 108064 22876
rect 107768 22822 107814 22874
rect 107814 22822 107824 22874
rect 107848 22822 107878 22874
rect 107878 22822 107890 22874
rect 107890 22822 107904 22874
rect 107928 22822 107942 22874
rect 107942 22822 107954 22874
rect 107954 22822 107984 22874
rect 108008 22822 108018 22874
rect 108018 22822 108064 22874
rect 107768 22820 107824 22822
rect 107848 22820 107904 22822
rect 107928 22820 107984 22822
rect 108008 22820 108064 22822
rect 107032 22330 107088 22332
rect 107112 22330 107168 22332
rect 107192 22330 107248 22332
rect 107272 22330 107328 22332
rect 107032 22278 107078 22330
rect 107078 22278 107088 22330
rect 107112 22278 107142 22330
rect 107142 22278 107154 22330
rect 107154 22278 107168 22330
rect 107192 22278 107206 22330
rect 107206 22278 107218 22330
rect 107218 22278 107248 22330
rect 107272 22278 107282 22330
rect 107282 22278 107328 22330
rect 107032 22276 107088 22278
rect 107112 22276 107168 22278
rect 107192 22276 107248 22278
rect 107272 22276 107328 22278
rect 107768 21786 107824 21788
rect 107848 21786 107904 21788
rect 107928 21786 107984 21788
rect 108008 21786 108064 21788
rect 107768 21734 107814 21786
rect 107814 21734 107824 21786
rect 107848 21734 107878 21786
rect 107878 21734 107890 21786
rect 107890 21734 107904 21786
rect 107928 21734 107942 21786
rect 107942 21734 107954 21786
rect 107954 21734 107984 21786
rect 108008 21734 108018 21786
rect 108018 21734 108064 21786
rect 107768 21732 107824 21734
rect 107848 21732 107904 21734
rect 107928 21732 107984 21734
rect 108008 21732 108064 21734
rect 107032 21242 107088 21244
rect 107112 21242 107168 21244
rect 107192 21242 107248 21244
rect 107272 21242 107328 21244
rect 107032 21190 107078 21242
rect 107078 21190 107088 21242
rect 107112 21190 107142 21242
rect 107142 21190 107154 21242
rect 107154 21190 107168 21242
rect 107192 21190 107206 21242
rect 107206 21190 107218 21242
rect 107218 21190 107248 21242
rect 107272 21190 107282 21242
rect 107282 21190 107328 21242
rect 107032 21188 107088 21190
rect 107112 21188 107168 21190
rect 107192 21188 107248 21190
rect 107272 21188 107328 21190
rect 107768 20698 107824 20700
rect 107848 20698 107904 20700
rect 107928 20698 107984 20700
rect 108008 20698 108064 20700
rect 107768 20646 107814 20698
rect 107814 20646 107824 20698
rect 107848 20646 107878 20698
rect 107878 20646 107890 20698
rect 107890 20646 107904 20698
rect 107928 20646 107942 20698
rect 107942 20646 107954 20698
rect 107954 20646 107984 20698
rect 108008 20646 108018 20698
rect 108018 20646 108064 20698
rect 107768 20644 107824 20646
rect 107848 20644 107904 20646
rect 107928 20644 107984 20646
rect 108008 20644 108064 20646
rect 107032 20154 107088 20156
rect 107112 20154 107168 20156
rect 107192 20154 107248 20156
rect 107272 20154 107328 20156
rect 107032 20102 107078 20154
rect 107078 20102 107088 20154
rect 107112 20102 107142 20154
rect 107142 20102 107154 20154
rect 107154 20102 107168 20154
rect 107192 20102 107206 20154
rect 107206 20102 107218 20154
rect 107218 20102 107248 20154
rect 107272 20102 107282 20154
rect 107282 20102 107328 20154
rect 107032 20100 107088 20102
rect 107112 20100 107168 20102
rect 107192 20100 107248 20102
rect 107272 20100 107328 20102
rect 107768 19610 107824 19612
rect 107848 19610 107904 19612
rect 107928 19610 107984 19612
rect 108008 19610 108064 19612
rect 107768 19558 107814 19610
rect 107814 19558 107824 19610
rect 107848 19558 107878 19610
rect 107878 19558 107890 19610
rect 107890 19558 107904 19610
rect 107928 19558 107942 19610
rect 107942 19558 107954 19610
rect 107954 19558 107984 19610
rect 108008 19558 108018 19610
rect 108018 19558 108064 19610
rect 107768 19556 107824 19558
rect 107848 19556 107904 19558
rect 107928 19556 107984 19558
rect 108008 19556 108064 19558
rect 107032 19066 107088 19068
rect 107112 19066 107168 19068
rect 107192 19066 107248 19068
rect 107272 19066 107328 19068
rect 107032 19014 107078 19066
rect 107078 19014 107088 19066
rect 107112 19014 107142 19066
rect 107142 19014 107154 19066
rect 107154 19014 107168 19066
rect 107192 19014 107206 19066
rect 107206 19014 107218 19066
rect 107218 19014 107248 19066
rect 107272 19014 107282 19066
rect 107282 19014 107328 19066
rect 107032 19012 107088 19014
rect 107112 19012 107168 19014
rect 107192 19012 107248 19014
rect 107272 19012 107328 19014
rect 107768 18522 107824 18524
rect 107848 18522 107904 18524
rect 107928 18522 107984 18524
rect 108008 18522 108064 18524
rect 107768 18470 107814 18522
rect 107814 18470 107824 18522
rect 107848 18470 107878 18522
rect 107878 18470 107890 18522
rect 107890 18470 107904 18522
rect 107928 18470 107942 18522
rect 107942 18470 107954 18522
rect 107954 18470 107984 18522
rect 108008 18470 108018 18522
rect 108018 18470 108064 18522
rect 107768 18468 107824 18470
rect 107848 18468 107904 18470
rect 107928 18468 107984 18470
rect 108008 18468 108064 18470
rect 107032 17978 107088 17980
rect 107112 17978 107168 17980
rect 107192 17978 107248 17980
rect 107272 17978 107328 17980
rect 107032 17926 107078 17978
rect 107078 17926 107088 17978
rect 107112 17926 107142 17978
rect 107142 17926 107154 17978
rect 107154 17926 107168 17978
rect 107192 17926 107206 17978
rect 107206 17926 107218 17978
rect 107218 17926 107248 17978
rect 107272 17926 107282 17978
rect 107282 17926 107328 17978
rect 107032 17924 107088 17926
rect 107112 17924 107168 17926
rect 107192 17924 107248 17926
rect 107272 17924 107328 17926
rect 107768 17434 107824 17436
rect 107848 17434 107904 17436
rect 107928 17434 107984 17436
rect 108008 17434 108064 17436
rect 107768 17382 107814 17434
rect 107814 17382 107824 17434
rect 107848 17382 107878 17434
rect 107878 17382 107890 17434
rect 107890 17382 107904 17434
rect 107928 17382 107942 17434
rect 107942 17382 107954 17434
rect 107954 17382 107984 17434
rect 108008 17382 108018 17434
rect 108018 17382 108064 17434
rect 107768 17380 107824 17382
rect 107848 17380 107904 17382
rect 107928 17380 107984 17382
rect 108008 17380 108064 17382
rect 107032 16890 107088 16892
rect 107112 16890 107168 16892
rect 107192 16890 107248 16892
rect 107272 16890 107328 16892
rect 107032 16838 107078 16890
rect 107078 16838 107088 16890
rect 107112 16838 107142 16890
rect 107142 16838 107154 16890
rect 107154 16838 107168 16890
rect 107192 16838 107206 16890
rect 107206 16838 107218 16890
rect 107218 16838 107248 16890
rect 107272 16838 107282 16890
rect 107282 16838 107328 16890
rect 107032 16836 107088 16838
rect 107112 16836 107168 16838
rect 107192 16836 107248 16838
rect 107272 16836 107328 16838
rect 107768 16346 107824 16348
rect 107848 16346 107904 16348
rect 107928 16346 107984 16348
rect 108008 16346 108064 16348
rect 107768 16294 107814 16346
rect 107814 16294 107824 16346
rect 107848 16294 107878 16346
rect 107878 16294 107890 16346
rect 107890 16294 107904 16346
rect 107928 16294 107942 16346
rect 107942 16294 107954 16346
rect 107954 16294 107984 16346
rect 108008 16294 108018 16346
rect 108018 16294 108064 16346
rect 107768 16292 107824 16294
rect 107848 16292 107904 16294
rect 107928 16292 107984 16294
rect 108008 16292 108064 16294
rect 107032 15802 107088 15804
rect 107112 15802 107168 15804
rect 107192 15802 107248 15804
rect 107272 15802 107328 15804
rect 107032 15750 107078 15802
rect 107078 15750 107088 15802
rect 107112 15750 107142 15802
rect 107142 15750 107154 15802
rect 107154 15750 107168 15802
rect 107192 15750 107206 15802
rect 107206 15750 107218 15802
rect 107218 15750 107248 15802
rect 107272 15750 107282 15802
rect 107282 15750 107328 15802
rect 107032 15748 107088 15750
rect 107112 15748 107168 15750
rect 107192 15748 107248 15750
rect 107272 15748 107328 15750
rect 107768 15258 107824 15260
rect 107848 15258 107904 15260
rect 107928 15258 107984 15260
rect 108008 15258 108064 15260
rect 107768 15206 107814 15258
rect 107814 15206 107824 15258
rect 107848 15206 107878 15258
rect 107878 15206 107890 15258
rect 107890 15206 107904 15258
rect 107928 15206 107942 15258
rect 107942 15206 107954 15258
rect 107954 15206 107984 15258
rect 108008 15206 108018 15258
rect 108018 15206 108064 15258
rect 107768 15204 107824 15206
rect 107848 15204 107904 15206
rect 107928 15204 107984 15206
rect 108008 15204 108064 15206
rect 107032 14714 107088 14716
rect 107112 14714 107168 14716
rect 107192 14714 107248 14716
rect 107272 14714 107328 14716
rect 107032 14662 107078 14714
rect 107078 14662 107088 14714
rect 107112 14662 107142 14714
rect 107142 14662 107154 14714
rect 107154 14662 107168 14714
rect 107192 14662 107206 14714
rect 107206 14662 107218 14714
rect 107218 14662 107248 14714
rect 107272 14662 107282 14714
rect 107282 14662 107328 14714
rect 107032 14660 107088 14662
rect 107112 14660 107168 14662
rect 107192 14660 107248 14662
rect 107272 14660 107328 14662
rect 107768 14170 107824 14172
rect 107848 14170 107904 14172
rect 107928 14170 107984 14172
rect 108008 14170 108064 14172
rect 107768 14118 107814 14170
rect 107814 14118 107824 14170
rect 107848 14118 107878 14170
rect 107878 14118 107890 14170
rect 107890 14118 107904 14170
rect 107928 14118 107942 14170
rect 107942 14118 107954 14170
rect 107954 14118 107984 14170
rect 108008 14118 108018 14170
rect 108018 14118 108064 14170
rect 107768 14116 107824 14118
rect 107848 14116 107904 14118
rect 107928 14116 107984 14118
rect 108008 14116 108064 14118
rect 107032 13626 107088 13628
rect 107112 13626 107168 13628
rect 107192 13626 107248 13628
rect 107272 13626 107328 13628
rect 107032 13574 107078 13626
rect 107078 13574 107088 13626
rect 107112 13574 107142 13626
rect 107142 13574 107154 13626
rect 107154 13574 107168 13626
rect 107192 13574 107206 13626
rect 107206 13574 107218 13626
rect 107218 13574 107248 13626
rect 107272 13574 107282 13626
rect 107282 13574 107328 13626
rect 107032 13572 107088 13574
rect 107112 13572 107168 13574
rect 107192 13572 107248 13574
rect 107272 13572 107328 13574
rect 107768 13082 107824 13084
rect 107848 13082 107904 13084
rect 107928 13082 107984 13084
rect 108008 13082 108064 13084
rect 107768 13030 107814 13082
rect 107814 13030 107824 13082
rect 107848 13030 107878 13082
rect 107878 13030 107890 13082
rect 107890 13030 107904 13082
rect 107928 13030 107942 13082
rect 107942 13030 107954 13082
rect 107954 13030 107984 13082
rect 108008 13030 108018 13082
rect 108018 13030 108064 13082
rect 107768 13028 107824 13030
rect 107848 13028 107904 13030
rect 107928 13028 107984 13030
rect 108008 13028 108064 13030
rect 107032 12538 107088 12540
rect 107112 12538 107168 12540
rect 107192 12538 107248 12540
rect 107272 12538 107328 12540
rect 107032 12486 107078 12538
rect 107078 12486 107088 12538
rect 107112 12486 107142 12538
rect 107142 12486 107154 12538
rect 107154 12486 107168 12538
rect 107192 12486 107206 12538
rect 107206 12486 107218 12538
rect 107218 12486 107248 12538
rect 107272 12486 107282 12538
rect 107282 12486 107328 12538
rect 107032 12484 107088 12486
rect 107112 12484 107168 12486
rect 107192 12484 107248 12486
rect 107272 12484 107328 12486
rect 107768 11994 107824 11996
rect 107848 11994 107904 11996
rect 107928 11994 107984 11996
rect 108008 11994 108064 11996
rect 107768 11942 107814 11994
rect 107814 11942 107824 11994
rect 107848 11942 107878 11994
rect 107878 11942 107890 11994
rect 107890 11942 107904 11994
rect 107928 11942 107942 11994
rect 107942 11942 107954 11994
rect 107954 11942 107984 11994
rect 108008 11942 108018 11994
rect 108018 11942 108064 11994
rect 107768 11940 107824 11942
rect 107848 11940 107904 11942
rect 107928 11940 107984 11942
rect 108008 11940 108064 11942
rect 107032 11450 107088 11452
rect 107112 11450 107168 11452
rect 107192 11450 107248 11452
rect 107272 11450 107328 11452
rect 107032 11398 107078 11450
rect 107078 11398 107088 11450
rect 107112 11398 107142 11450
rect 107142 11398 107154 11450
rect 107154 11398 107168 11450
rect 107192 11398 107206 11450
rect 107206 11398 107218 11450
rect 107218 11398 107248 11450
rect 107272 11398 107282 11450
rect 107282 11398 107328 11450
rect 107032 11396 107088 11398
rect 107112 11396 107168 11398
rect 107192 11396 107248 11398
rect 107272 11396 107328 11398
rect 107768 10906 107824 10908
rect 107848 10906 107904 10908
rect 107928 10906 107984 10908
rect 108008 10906 108064 10908
rect 107768 10854 107814 10906
rect 107814 10854 107824 10906
rect 107848 10854 107878 10906
rect 107878 10854 107890 10906
rect 107890 10854 107904 10906
rect 107928 10854 107942 10906
rect 107942 10854 107954 10906
rect 107954 10854 107984 10906
rect 108008 10854 108018 10906
rect 108018 10854 108064 10906
rect 107768 10852 107824 10854
rect 107848 10852 107904 10854
rect 107928 10852 107984 10854
rect 108008 10852 108064 10854
rect 107032 10362 107088 10364
rect 107112 10362 107168 10364
rect 107192 10362 107248 10364
rect 107272 10362 107328 10364
rect 107032 10310 107078 10362
rect 107078 10310 107088 10362
rect 107112 10310 107142 10362
rect 107142 10310 107154 10362
rect 107154 10310 107168 10362
rect 107192 10310 107206 10362
rect 107206 10310 107218 10362
rect 107218 10310 107248 10362
rect 107272 10310 107282 10362
rect 107282 10310 107328 10362
rect 107032 10308 107088 10310
rect 107112 10308 107168 10310
rect 107192 10308 107248 10310
rect 107272 10308 107328 10310
rect 110418 10240 110474 10296
rect 104254 9832 104310 9888
rect 107768 9818 107824 9820
rect 107848 9818 107904 9820
rect 107928 9818 107984 9820
rect 108008 9818 108064 9820
rect 107768 9766 107814 9818
rect 107814 9766 107824 9818
rect 107848 9766 107878 9818
rect 107878 9766 107890 9818
rect 107890 9766 107904 9818
rect 107928 9766 107942 9818
rect 107942 9766 107954 9818
rect 107954 9766 107984 9818
rect 108008 9766 108018 9818
rect 108018 9766 108064 9818
rect 107768 9764 107824 9766
rect 107848 9764 107904 9766
rect 107928 9764 107984 9766
rect 108008 9764 108064 9766
rect 90730 9424 90786 9480
rect 32862 8064 32918 8120
rect 35254 8064 35310 8120
rect 38658 8064 38714 8120
rect 28262 7520 28264 7540
rect 28264 7520 28316 7540
rect 28316 7520 28318 7540
rect 33966 7540 34022 7576
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 33966 7520 33968 7540
rect 33968 7520 34020 7540
rect 34020 7520 34022 7540
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36358 7540 36414 7576
rect 36358 7520 36360 7540
rect 36360 7520 36412 7540
rect 36412 7520 36414 7540
rect 37462 7540 37518 7576
rect 66320 7642 66376 7644
rect 66400 7642 66456 7644
rect 66480 7642 66536 7644
rect 66560 7642 66616 7644
rect 66320 7590 66366 7642
rect 66366 7590 66376 7642
rect 66400 7590 66430 7642
rect 66430 7590 66442 7642
rect 66442 7590 66456 7642
rect 66480 7590 66494 7642
rect 66494 7590 66506 7642
rect 66506 7590 66536 7642
rect 66560 7590 66570 7642
rect 66570 7590 66616 7642
rect 66320 7588 66376 7590
rect 66400 7588 66456 7590
rect 66480 7588 66536 7590
rect 66560 7588 66616 7590
rect 37462 7520 37464 7540
rect 37464 7520 37516 7540
rect 37516 7520 37518 7540
rect 39854 7540 39910 7576
rect 39854 7520 39856 7540
rect 39856 7520 39908 7540
rect 39908 7520 39910 7540
rect 41050 7540 41106 7576
rect 41050 7520 41052 7540
rect 41052 7520 41104 7540
rect 41104 7520 41106 7540
rect 42154 7540 42210 7576
rect 42154 7520 42156 7540
rect 42156 7520 42208 7540
rect 42208 7520 42210 7540
rect 43350 7540 43406 7576
rect 43350 7520 43352 7540
rect 43352 7520 43404 7540
rect 43404 7520 43406 7540
rect 90546 7540 90602 7576
rect 107032 9274 107088 9276
rect 107112 9274 107168 9276
rect 107192 9274 107248 9276
rect 107272 9274 107328 9276
rect 107032 9222 107078 9274
rect 107078 9222 107088 9274
rect 107112 9222 107142 9274
rect 107142 9222 107154 9274
rect 107154 9222 107168 9274
rect 107192 9222 107206 9274
rect 107206 9222 107218 9274
rect 107218 9222 107248 9274
rect 107272 9222 107282 9274
rect 107282 9222 107328 9274
rect 107032 9220 107088 9222
rect 107112 9220 107168 9222
rect 107192 9220 107248 9222
rect 107272 9220 107328 9222
rect 107768 8730 107824 8732
rect 107848 8730 107904 8732
rect 107928 8730 107984 8732
rect 108008 8730 108064 8732
rect 107768 8678 107814 8730
rect 107814 8678 107824 8730
rect 107848 8678 107878 8730
rect 107878 8678 107890 8730
rect 107890 8678 107904 8730
rect 107928 8678 107942 8730
rect 107942 8678 107954 8730
rect 107954 8678 107984 8730
rect 108008 8678 108018 8730
rect 108018 8678 108064 8730
rect 107768 8676 107824 8678
rect 107848 8676 107904 8678
rect 107928 8676 107984 8678
rect 108008 8676 108064 8678
rect 107032 8186 107088 8188
rect 107112 8186 107168 8188
rect 107192 8186 107248 8188
rect 107272 8186 107328 8188
rect 107032 8134 107078 8186
rect 107078 8134 107088 8186
rect 107112 8134 107142 8186
rect 107142 8134 107154 8186
rect 107154 8134 107168 8186
rect 107192 8134 107206 8186
rect 107206 8134 107218 8186
rect 107218 8134 107248 8186
rect 107272 8134 107282 8186
rect 107282 8134 107328 8186
rect 107032 8132 107088 8134
rect 107112 8132 107168 8134
rect 107192 8132 107248 8134
rect 107272 8132 107328 8134
rect 97040 7642 97096 7644
rect 97120 7642 97176 7644
rect 97200 7642 97256 7644
rect 97280 7642 97336 7644
rect 97040 7590 97086 7642
rect 97086 7590 97096 7642
rect 97120 7590 97150 7642
rect 97150 7590 97162 7642
rect 97162 7590 97176 7642
rect 97200 7590 97214 7642
rect 97214 7590 97226 7642
rect 97226 7590 97256 7642
rect 97280 7590 97290 7642
rect 97290 7590 97336 7642
rect 97040 7588 97096 7590
rect 97120 7588 97176 7590
rect 97200 7588 97256 7590
rect 97280 7588 97336 7590
rect 107768 7642 107824 7644
rect 107848 7642 107904 7644
rect 107928 7642 107984 7644
rect 108008 7642 108064 7644
rect 107768 7590 107814 7642
rect 107814 7590 107824 7642
rect 107848 7590 107878 7642
rect 107878 7590 107890 7642
rect 107890 7590 107904 7642
rect 107928 7590 107942 7642
rect 107942 7590 107954 7642
rect 107954 7590 107984 7642
rect 108008 7590 108018 7642
rect 108018 7590 108064 7642
rect 107768 7588 107824 7590
rect 107848 7588 107904 7590
rect 107928 7588 107984 7590
rect 108008 7588 108064 7590
rect 90546 7520 90548 7540
rect 90548 7520 90600 7540
rect 90600 7520 90602 7540
rect 91006 7540 91062 7576
rect 91006 7520 91008 7540
rect 91008 7520 91060 7540
rect 91060 7520 91062 7540
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 107032 7098 107088 7100
rect 107112 7098 107168 7100
rect 107192 7098 107248 7100
rect 107272 7098 107328 7100
rect 107032 7046 107078 7098
rect 107078 7046 107088 7098
rect 107112 7046 107142 7098
rect 107142 7046 107154 7098
rect 107154 7046 107168 7098
rect 107192 7046 107206 7098
rect 107206 7046 107218 7098
rect 107218 7046 107248 7098
rect 107272 7046 107282 7098
rect 107282 7046 107328 7098
rect 107032 7044 107088 7046
rect 107112 7044 107168 7046
rect 107192 7044 107248 7046
rect 107272 7044 107328 7046
rect 66320 6554 66376 6556
rect 66400 6554 66456 6556
rect 66480 6554 66536 6556
rect 66560 6554 66616 6556
rect 66320 6502 66366 6554
rect 66366 6502 66376 6554
rect 66400 6502 66430 6554
rect 66430 6502 66442 6554
rect 66442 6502 66456 6554
rect 66480 6502 66494 6554
rect 66494 6502 66506 6554
rect 66506 6502 66536 6554
rect 66560 6502 66570 6554
rect 66570 6502 66616 6554
rect 66320 6500 66376 6502
rect 66400 6500 66456 6502
rect 66480 6500 66536 6502
rect 66560 6500 66616 6502
rect 97040 6554 97096 6556
rect 97120 6554 97176 6556
rect 97200 6554 97256 6556
rect 97280 6554 97336 6556
rect 97040 6502 97086 6554
rect 97086 6502 97096 6554
rect 97120 6502 97150 6554
rect 97150 6502 97162 6554
rect 97162 6502 97176 6554
rect 97200 6502 97214 6554
rect 97214 6502 97226 6554
rect 97226 6502 97256 6554
rect 97280 6502 97290 6554
rect 97290 6502 97336 6554
rect 97040 6500 97096 6502
rect 97120 6500 97176 6502
rect 97200 6500 97256 6502
rect 97280 6500 97336 6502
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 66320 5466 66376 5468
rect 66400 5466 66456 5468
rect 66480 5466 66536 5468
rect 66560 5466 66616 5468
rect 66320 5414 66366 5466
rect 66366 5414 66376 5466
rect 66400 5414 66430 5466
rect 66430 5414 66442 5466
rect 66442 5414 66456 5466
rect 66480 5414 66494 5466
rect 66494 5414 66506 5466
rect 66506 5414 66536 5466
rect 66560 5414 66570 5466
rect 66570 5414 66616 5466
rect 66320 5412 66376 5414
rect 66400 5412 66456 5414
rect 66480 5412 66536 5414
rect 66560 5412 66616 5414
rect 97040 5466 97096 5468
rect 97120 5466 97176 5468
rect 97200 5466 97256 5468
rect 97280 5466 97336 5468
rect 97040 5414 97086 5466
rect 97086 5414 97096 5466
rect 97120 5414 97150 5466
rect 97150 5414 97162 5466
rect 97162 5414 97176 5466
rect 97200 5414 97214 5466
rect 97214 5414 97226 5466
rect 97226 5414 97256 5466
rect 97280 5414 97290 5466
rect 97290 5414 97336 5466
rect 97040 5412 97096 5414
rect 97120 5412 97176 5414
rect 97200 5412 97256 5414
rect 97280 5412 97336 5414
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 66320 4378 66376 4380
rect 66400 4378 66456 4380
rect 66480 4378 66536 4380
rect 66560 4378 66616 4380
rect 66320 4326 66366 4378
rect 66366 4326 66376 4378
rect 66400 4326 66430 4378
rect 66430 4326 66442 4378
rect 66442 4326 66456 4378
rect 66480 4326 66494 4378
rect 66494 4326 66506 4378
rect 66506 4326 66536 4378
rect 66560 4326 66570 4378
rect 66570 4326 66616 4378
rect 66320 4324 66376 4326
rect 66400 4324 66456 4326
rect 66480 4324 66536 4326
rect 66560 4324 66616 4326
rect 97040 4378 97096 4380
rect 97120 4378 97176 4380
rect 97200 4378 97256 4380
rect 97280 4378 97336 4380
rect 97040 4326 97086 4378
rect 97086 4326 97096 4378
rect 97120 4326 97150 4378
rect 97150 4326 97162 4378
rect 97162 4326 97176 4378
rect 97200 4326 97214 4378
rect 97214 4326 97226 4378
rect 97226 4326 97256 4378
rect 97280 4326 97290 4378
rect 97290 4326 97336 4378
rect 97040 4324 97096 4326
rect 97120 4324 97176 4326
rect 97200 4324 97256 4326
rect 97280 4324 97336 4326
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 66320 3290 66376 3292
rect 66400 3290 66456 3292
rect 66480 3290 66536 3292
rect 66560 3290 66616 3292
rect 66320 3238 66366 3290
rect 66366 3238 66376 3290
rect 66400 3238 66430 3290
rect 66430 3238 66442 3290
rect 66442 3238 66456 3290
rect 66480 3238 66494 3290
rect 66494 3238 66506 3290
rect 66506 3238 66536 3290
rect 66560 3238 66570 3290
rect 66570 3238 66616 3290
rect 66320 3236 66376 3238
rect 66400 3236 66456 3238
rect 66480 3236 66536 3238
rect 66560 3236 66616 3238
rect 97040 3290 97096 3292
rect 97120 3290 97176 3292
rect 97200 3290 97256 3292
rect 97280 3290 97336 3292
rect 97040 3238 97086 3290
rect 97086 3238 97096 3290
rect 97120 3238 97150 3290
rect 97150 3238 97162 3290
rect 97162 3238 97176 3290
rect 97200 3238 97214 3290
rect 97214 3238 97226 3290
rect 97226 3238 97256 3290
rect 97280 3238 97290 3290
rect 97290 3238 97336 3290
rect 97040 3236 97096 3238
rect 97120 3236 97176 3238
rect 97200 3236 97256 3238
rect 97280 3236 97336 3238
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 66320 2202 66376 2204
rect 66400 2202 66456 2204
rect 66480 2202 66536 2204
rect 66560 2202 66616 2204
rect 66320 2150 66366 2202
rect 66366 2150 66376 2202
rect 66400 2150 66430 2202
rect 66430 2150 66442 2202
rect 66442 2150 66456 2202
rect 66480 2150 66494 2202
rect 66494 2150 66506 2202
rect 66506 2150 66536 2202
rect 66560 2150 66570 2202
rect 66570 2150 66616 2202
rect 66320 2148 66376 2150
rect 66400 2148 66456 2150
rect 66480 2148 66536 2150
rect 66560 2148 66616 2150
rect 97040 2202 97096 2204
rect 97120 2202 97176 2204
rect 97200 2202 97256 2204
rect 97280 2202 97336 2204
rect 97040 2150 97086 2202
rect 97086 2150 97096 2202
rect 97120 2150 97150 2202
rect 97150 2150 97162 2202
rect 97162 2150 97176 2202
rect 97200 2150 97214 2202
rect 97214 2150 97226 2202
rect 97226 2150 97256 2202
rect 97280 2150 97290 2202
rect 97290 2150 97336 2202
rect 97040 2148 97096 2150
rect 97120 2148 97176 2150
rect 97200 2148 97256 2150
rect 97280 2148 97336 2150
<< metal3 >>
rect 4870 71840 5186 71841
rect 4870 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5186 71840
rect 4870 71775 5186 71776
rect 35590 71840 35906 71841
rect 35590 71776 35596 71840
rect 35660 71776 35676 71840
rect 35740 71776 35756 71840
rect 35820 71776 35836 71840
rect 35900 71776 35906 71840
rect 35590 71775 35906 71776
rect 66310 71840 66626 71841
rect 66310 71776 66316 71840
rect 66380 71776 66396 71840
rect 66460 71776 66476 71840
rect 66540 71776 66556 71840
rect 66620 71776 66626 71840
rect 66310 71775 66626 71776
rect 97030 71840 97346 71841
rect 97030 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97346 71840
rect 97030 71775 97346 71776
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 34930 71296 35246 71297
rect 34930 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35246 71296
rect 34930 71231 35246 71232
rect 65650 71296 65966 71297
rect 65650 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65966 71296
rect 65650 71231 65966 71232
rect 96370 71296 96686 71297
rect 96370 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96686 71296
rect 96370 71231 96686 71232
rect 4870 70752 5186 70753
rect 4870 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5186 70752
rect 4870 70687 5186 70688
rect 35590 70752 35906 70753
rect 35590 70688 35596 70752
rect 35660 70688 35676 70752
rect 35740 70688 35756 70752
rect 35820 70688 35836 70752
rect 35900 70688 35906 70752
rect 35590 70687 35906 70688
rect 66310 70752 66626 70753
rect 66310 70688 66316 70752
rect 66380 70688 66396 70752
rect 66460 70688 66476 70752
rect 66540 70688 66556 70752
rect 66620 70688 66626 70752
rect 66310 70687 66626 70688
rect 97030 70752 97346 70753
rect 97030 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97346 70752
rect 97030 70687 97346 70688
rect 4210 70208 4526 70209
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 34930 70208 35246 70209
rect 34930 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35246 70208
rect 34930 70143 35246 70144
rect 65650 70208 65966 70209
rect 65650 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65966 70208
rect 65650 70143 65966 70144
rect 96370 70208 96686 70209
rect 96370 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96686 70208
rect 96370 70143 96686 70144
rect 4870 69664 5186 69665
rect 4870 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5186 69664
rect 4870 69599 5186 69600
rect 35590 69664 35906 69665
rect 35590 69600 35596 69664
rect 35660 69600 35676 69664
rect 35740 69600 35756 69664
rect 35820 69600 35836 69664
rect 35900 69600 35906 69664
rect 35590 69599 35906 69600
rect 66310 69664 66626 69665
rect 66310 69600 66316 69664
rect 66380 69600 66396 69664
rect 66460 69600 66476 69664
rect 66540 69600 66556 69664
rect 66620 69600 66626 69664
rect 66310 69599 66626 69600
rect 97030 69664 97346 69665
rect 97030 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97346 69664
rect 97030 69599 97346 69600
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 34930 69120 35246 69121
rect 34930 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35246 69120
rect 34930 69055 35246 69056
rect 65650 69120 65966 69121
rect 65650 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65966 69120
rect 65650 69055 65966 69056
rect 96370 69120 96686 69121
rect 96370 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96686 69120
rect 96370 69055 96686 69056
rect 4870 68576 5186 68577
rect 4870 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5186 68576
rect 4870 68511 5186 68512
rect 35590 68576 35906 68577
rect 35590 68512 35596 68576
rect 35660 68512 35676 68576
rect 35740 68512 35756 68576
rect 35820 68512 35836 68576
rect 35900 68512 35906 68576
rect 35590 68511 35906 68512
rect 66310 68576 66626 68577
rect 66310 68512 66316 68576
rect 66380 68512 66396 68576
rect 66460 68512 66476 68576
rect 66540 68512 66556 68576
rect 66620 68512 66626 68576
rect 66310 68511 66626 68512
rect 97030 68576 97346 68577
rect 97030 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97346 68576
rect 97030 68511 97346 68512
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 34930 68032 35246 68033
rect 34930 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35246 68032
rect 34930 67967 35246 67968
rect 65650 68032 65966 68033
rect 65650 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65966 68032
rect 65650 67967 65966 67968
rect 96370 68032 96686 68033
rect 96370 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96686 68032
rect 96370 67967 96686 67968
rect 4870 67488 5186 67489
rect 4870 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5186 67488
rect 4870 67423 5186 67424
rect 35590 67488 35906 67489
rect 35590 67424 35596 67488
rect 35660 67424 35676 67488
rect 35740 67424 35756 67488
rect 35820 67424 35836 67488
rect 35900 67424 35906 67488
rect 35590 67423 35906 67424
rect 66310 67488 66626 67489
rect 66310 67424 66316 67488
rect 66380 67424 66396 67488
rect 66460 67424 66476 67488
rect 66540 67424 66556 67488
rect 66620 67424 66626 67488
rect 66310 67423 66626 67424
rect 97030 67488 97346 67489
rect 97030 67424 97036 67488
rect 97100 67424 97116 67488
rect 97180 67424 97196 67488
rect 97260 67424 97276 67488
rect 97340 67424 97346 67488
rect 97030 67423 97346 67424
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 96370 66944 96686 66945
rect 96370 66880 96376 66944
rect 96440 66880 96456 66944
rect 96520 66880 96536 66944
rect 96600 66880 96616 66944
rect 96680 66880 96686 66944
rect 96370 66879 96686 66880
rect 51022 66676 51028 66740
rect 51092 66738 51098 66740
rect 55673 66738 55739 66741
rect 51092 66736 55739 66738
rect 51092 66680 55678 66736
rect 55734 66680 55739 66736
rect 51092 66678 55739 66680
rect 51092 66676 51098 66678
rect 55673 66675 55739 66678
rect 66110 66540 66116 66604
rect 66180 66602 66186 66604
rect 68461 66602 68527 66605
rect 66180 66600 68527 66602
rect 66180 66544 68466 66600
rect 68522 66544 68527 66600
rect 66180 66542 68527 66544
rect 66180 66540 66186 66542
rect 68461 66539 68527 66542
rect 48630 66404 48636 66468
rect 48700 66466 48706 66468
rect 53649 66466 53715 66469
rect 48700 66464 53715 66466
rect 48700 66408 53654 66464
rect 53710 66408 53715 66464
rect 48700 66406 53715 66408
rect 48700 66404 48706 66406
rect 53649 66403 53715 66406
rect 55990 66404 55996 66468
rect 56060 66466 56066 66468
rect 59997 66466 60063 66469
rect 56060 66464 60063 66466
rect 56060 66408 60002 66464
rect 60058 66408 60063 66464
rect 56060 66406 60063 66408
rect 56060 66404 56066 66406
rect 59997 66403 60063 66406
rect 61142 66404 61148 66468
rect 61212 66466 61218 66468
rect 63953 66466 64019 66469
rect 61212 66464 64019 66466
rect 61212 66408 63958 66464
rect 64014 66408 64019 66464
rect 61212 66406 64019 66408
rect 61212 66404 61218 66406
rect 63953 66403 64019 66406
rect 4870 66400 5186 66401
rect 4870 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5186 66400
rect 4870 66335 5186 66336
rect 35590 66400 35906 66401
rect 35590 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35906 66400
rect 35590 66335 35906 66336
rect 66310 66400 66626 66401
rect 66310 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66626 66400
rect 66310 66335 66626 66336
rect 97030 66400 97346 66401
rect 97030 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97346 66400
rect 97030 66335 97346 66336
rect 107758 66400 108074 66401
rect 107758 66336 107764 66400
rect 107828 66336 107844 66400
rect 107908 66336 107924 66400
rect 107988 66336 108004 66400
rect 108068 66336 108074 66400
rect 107758 66335 108074 66336
rect 46054 66268 46060 66332
rect 46124 66330 46130 66332
rect 49693 66330 49759 66333
rect 46124 66328 49759 66330
rect 46124 66272 49698 66328
rect 49754 66272 49759 66328
rect 46124 66270 49759 66272
rect 46124 66268 46130 66270
rect 49693 66267 49759 66270
rect 58566 66268 58572 66332
rect 58636 66330 58642 66332
rect 61653 66330 61719 66333
rect 58636 66328 61719 66330
rect 58636 66272 61658 66328
rect 61714 66272 61719 66328
rect 58636 66270 61719 66272
rect 58636 66268 58642 66270
rect 61653 66267 61719 66270
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 96370 65856 96686 65857
rect 96370 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96686 65856
rect 96370 65791 96686 65792
rect 107022 65856 107338 65857
rect 107022 65792 107028 65856
rect 107092 65792 107108 65856
rect 107172 65792 107188 65856
rect 107252 65792 107268 65856
rect 107332 65792 107338 65856
rect 107022 65791 107338 65792
rect 63534 65452 63540 65516
rect 63604 65514 63610 65516
rect 64689 65514 64755 65517
rect 63604 65512 64755 65514
rect 63604 65456 64694 65512
rect 64750 65456 64755 65512
rect 63604 65454 64755 65456
rect 63604 65452 63610 65454
rect 64689 65451 64755 65454
rect 68502 65316 68508 65380
rect 68572 65378 68578 65380
rect 68737 65378 68803 65381
rect 68572 65376 68803 65378
rect 68572 65320 68742 65376
rect 68798 65320 68803 65376
rect 68572 65318 68803 65320
rect 68572 65316 68578 65318
rect 68737 65315 68803 65318
rect 73470 65316 73476 65380
rect 73540 65378 73546 65380
rect 74073 65378 74139 65381
rect 87321 65380 87387 65381
rect 87270 65378 87276 65380
rect 73540 65376 74139 65378
rect 73540 65320 74078 65376
rect 74134 65320 74139 65376
rect 73540 65318 74139 65320
rect 87230 65318 87276 65378
rect 87340 65376 87387 65380
rect 87382 65320 87387 65376
rect 73540 65316 73546 65318
rect 74073 65315 74139 65318
rect 87270 65316 87276 65318
rect 87340 65316 87387 65320
rect 87321 65315 87387 65316
rect 4870 65312 5186 65313
rect 4870 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5186 65312
rect 4870 65247 5186 65248
rect 107758 65312 108074 65313
rect 107758 65248 107764 65312
rect 107828 65248 107844 65312
rect 107908 65248 107924 65312
rect 107988 65248 108004 65312
rect 108068 65248 108074 65312
rect 107758 65247 108074 65248
rect 71078 65044 71084 65108
rect 71148 65106 71154 65108
rect 71221 65106 71287 65109
rect 71148 65104 71287 65106
rect 71148 65048 71226 65104
rect 71282 65048 71287 65104
rect 71148 65046 71287 65048
rect 71148 65044 71154 65046
rect 71221 65043 71287 65046
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 107022 64768 107338 64769
rect 107022 64704 107028 64768
rect 107092 64704 107108 64768
rect 107172 64704 107188 64768
rect 107252 64704 107268 64768
rect 107332 64704 107338 64768
rect 107022 64703 107338 64704
rect 4870 64224 5186 64225
rect 4870 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5186 64224
rect 4870 64159 5186 64160
rect 107758 64224 108074 64225
rect 107758 64160 107764 64224
rect 107828 64160 107844 64224
rect 107908 64160 107924 64224
rect 107988 64160 108004 64224
rect 108068 64160 108074 64224
rect 107758 64159 108074 64160
rect 36069 64092 36075 64156
rect 36139 64154 36145 64156
rect 43161 64154 43227 64157
rect 36139 64152 43227 64154
rect 36139 64096 43166 64152
rect 43222 64096 43227 64152
rect 36139 64094 43227 64096
rect 36139 64092 36145 64094
rect 43161 64091 43227 64094
rect 43570 64092 43576 64156
rect 43640 64154 43646 64156
rect 49969 64154 50035 64157
rect 43640 64152 50035 64154
rect 43640 64096 49974 64152
rect 50030 64096 50035 64152
rect 43640 64094 50035 64096
rect 43640 64092 43646 64094
rect 49969 64091 50035 64094
rect 87304 64092 87310 64156
rect 87374 64154 87380 64156
rect 104985 64154 105051 64157
rect 87374 64152 105051 64154
rect 87374 64096 104990 64152
rect 105046 64096 105051 64152
rect 87374 64094 105051 64096
rect 87374 64092 87380 64094
rect 104985 64091 105051 64094
rect 41061 63956 41067 64020
rect 41131 64018 41137 64020
rect 47577 64018 47643 64021
rect 41131 64016 47643 64018
rect 41131 63960 47582 64016
rect 47638 63960 47643 64016
rect 41131 63958 47643 63960
rect 41131 63956 41137 63958
rect 47577 63955 47643 63958
rect 86136 63956 86142 64020
rect 86206 64018 86212 64020
rect 86309 64018 86375 64021
rect 106181 64018 106247 64021
rect 86206 64016 106247 64018
rect 86206 63960 86314 64016
rect 86370 63960 106186 64016
rect 106242 63960 106247 64016
rect 86206 63958 106247 63960
rect 86206 63956 86212 63958
rect 86309 63955 86375 63958
rect 106181 63955 106247 63958
rect 38565 63820 38571 63884
rect 38635 63882 38641 63884
rect 45369 63882 45435 63885
rect 38635 63880 45435 63882
rect 38635 63824 45374 63880
rect 45430 63824 45435 63880
rect 38635 63822 45435 63824
rect 38635 63820 38641 63822
rect 45369 63819 45435 63822
rect 53541 63820 53547 63884
rect 53611 63882 53617 63884
rect 58157 63882 58223 63885
rect 95877 63884 95943 63885
rect 95852 63882 95858 63884
rect 53611 63880 58223 63882
rect 53611 63824 58162 63880
rect 58218 63824 58223 63880
rect 53611 63822 58223 63824
rect 95786 63822 95858 63882
rect 95922 63882 95943 63884
rect 104341 63882 104407 63885
rect 95922 63880 104407 63882
rect 95938 63824 104346 63880
rect 104402 63824 104407 63880
rect 53611 63820 53617 63822
rect 58157 63819 58223 63822
rect 95852 63820 95858 63822
rect 95922 63822 104407 63824
rect 95922 63820 95943 63822
rect 95877 63819 95943 63820
rect 104341 63819 104407 63822
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 107022 63680 107338 63681
rect 107022 63616 107028 63680
rect 107092 63616 107108 63680
rect 107172 63616 107188 63680
rect 107252 63616 107268 63680
rect 107332 63616 107338 63680
rect 107022 63615 107338 63616
rect 4870 63136 5186 63137
rect 4870 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5186 63136
rect 4870 63071 5186 63072
rect 107758 63136 108074 63137
rect 107758 63072 107764 63136
rect 107828 63072 107844 63136
rect 107908 63072 107924 63136
rect 107988 63072 108004 63136
rect 108068 63072 108074 63136
rect 107758 63071 108074 63072
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 107022 62592 107338 62593
rect 107022 62528 107028 62592
rect 107092 62528 107108 62592
rect 107172 62528 107188 62592
rect 107252 62528 107268 62592
rect 107332 62528 107338 62592
rect 107022 62527 107338 62528
rect 4870 62048 5186 62049
rect 4870 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5186 62048
rect 4870 61983 5186 61984
rect 107758 62048 108074 62049
rect 107758 61984 107764 62048
rect 107828 61984 107844 62048
rect 107908 61984 107924 62048
rect 107988 61984 108004 62048
rect 108068 61984 108074 62048
rect 107758 61983 108074 61984
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 107022 61504 107338 61505
rect 107022 61440 107028 61504
rect 107092 61440 107108 61504
rect 107172 61440 107188 61504
rect 107252 61440 107268 61504
rect 107332 61440 107338 61504
rect 107022 61439 107338 61440
rect 4870 60960 5186 60961
rect 4870 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5186 60960
rect 4870 60895 5186 60896
rect 107758 60960 108074 60961
rect 107758 60896 107764 60960
rect 107828 60896 107844 60960
rect 107908 60896 107924 60960
rect 107988 60896 108004 60960
rect 108068 60896 108074 60960
rect 107758 60895 108074 60896
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 107022 60416 107338 60417
rect 107022 60352 107028 60416
rect 107092 60352 107108 60416
rect 107172 60352 107188 60416
rect 107252 60352 107268 60416
rect 107332 60352 107338 60416
rect 107022 60351 107338 60352
rect 4870 59872 5186 59873
rect 4870 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5186 59872
rect 4870 59807 5186 59808
rect 107758 59872 108074 59873
rect 107758 59808 107764 59872
rect 107828 59808 107844 59872
rect 107908 59808 107924 59872
rect 107988 59808 108004 59872
rect 108068 59808 108074 59872
rect 107758 59807 108074 59808
rect 103697 59802 103763 59805
rect 102550 59800 103763 59802
rect 102550 59768 103702 59800
rect 101948 59744 103702 59768
rect 103758 59744 103763 59800
rect 101948 59742 103763 59744
rect 101948 59708 102610 59742
rect 103697 59739 103763 59742
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 107022 59328 107338 59329
rect 107022 59264 107028 59328
rect 107092 59264 107108 59328
rect 107172 59264 107188 59328
rect 107252 59264 107268 59328
rect 107332 59264 107338 59328
rect 107022 59263 107338 59264
rect 4870 58784 5186 58785
rect 4870 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5186 58784
rect 4870 58719 5186 58720
rect 107758 58784 108074 58785
rect 107758 58720 107764 58784
rect 107828 58720 107844 58784
rect 107908 58720 107924 58784
rect 107988 58720 108004 58784
rect 108068 58720 108074 58784
rect 107758 58719 108074 58720
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 107022 58240 107338 58241
rect 107022 58176 107028 58240
rect 107092 58176 107108 58240
rect 107172 58176 107188 58240
rect 107252 58176 107268 58240
rect 107332 58176 107338 58240
rect 107022 58175 107338 58176
rect 4870 57696 5186 57697
rect 4870 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5186 57696
rect 4870 57631 5186 57632
rect 107758 57696 108074 57697
rect 107758 57632 107764 57696
rect 107828 57632 107844 57696
rect 107908 57632 107924 57696
rect 107988 57632 108004 57696
rect 108068 57632 108074 57696
rect 107758 57631 108074 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 107022 57152 107338 57153
rect 107022 57088 107028 57152
rect 107092 57088 107108 57152
rect 107172 57088 107188 57152
rect 107252 57088 107268 57152
rect 107332 57088 107338 57152
rect 107022 57087 107338 57088
rect 4870 56608 5186 56609
rect 4870 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5186 56608
rect 4870 56543 5186 56544
rect 107758 56608 108074 56609
rect 107758 56544 107764 56608
rect 107828 56544 107844 56608
rect 107908 56544 107924 56608
rect 107988 56544 108004 56608
rect 108068 56544 108074 56608
rect 107758 56543 108074 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 107022 56064 107338 56065
rect 107022 56000 107028 56064
rect 107092 56000 107108 56064
rect 107172 56000 107188 56064
rect 107252 56000 107268 56064
rect 107332 56000 107338 56064
rect 107022 55999 107338 56000
rect 4870 55520 5186 55521
rect 4870 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5186 55520
rect 4870 55455 5186 55456
rect 107758 55520 108074 55521
rect 107758 55456 107764 55520
rect 107828 55456 107844 55520
rect 107908 55456 107924 55520
rect 107988 55456 108004 55520
rect 108068 55456 108074 55520
rect 107758 55455 108074 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 107022 54976 107338 54977
rect 107022 54912 107028 54976
rect 107092 54912 107108 54976
rect 107172 54912 107188 54976
rect 107252 54912 107268 54976
rect 107332 54912 107338 54976
rect 107022 54911 107338 54912
rect 4870 54432 5186 54433
rect 4870 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5186 54432
rect 4870 54367 5186 54368
rect 107758 54432 108074 54433
rect 107758 54368 107764 54432
rect 107828 54368 107844 54432
rect 107908 54368 107924 54432
rect 107988 54368 108004 54432
rect 108068 54368 108074 54432
rect 107758 54367 108074 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 107022 53888 107338 53889
rect 107022 53824 107028 53888
rect 107092 53824 107108 53888
rect 107172 53824 107188 53888
rect 107252 53824 107268 53888
rect 107332 53824 107338 53888
rect 107022 53823 107338 53824
rect 4870 53344 5186 53345
rect 4870 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5186 53344
rect 4870 53279 5186 53280
rect 107758 53344 108074 53345
rect 107758 53280 107764 53344
rect 107828 53280 107844 53344
rect 107908 53280 107924 53344
rect 107988 53280 108004 53344
rect 108068 53280 108074 53344
rect 107758 53279 108074 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 107022 52800 107338 52801
rect 107022 52736 107028 52800
rect 107092 52736 107108 52800
rect 107172 52736 107188 52800
rect 107252 52736 107268 52800
rect 107332 52736 107338 52800
rect 107022 52735 107338 52736
rect 4870 52256 5186 52257
rect 4870 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5186 52256
rect 4870 52191 5186 52192
rect 107758 52256 108074 52257
rect 107758 52192 107764 52256
rect 107828 52192 107844 52256
rect 107908 52192 107924 52256
rect 107988 52192 108004 52256
rect 108068 52192 108074 52256
rect 107758 52191 108074 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 107022 51712 107338 51713
rect 107022 51648 107028 51712
rect 107092 51648 107108 51712
rect 107172 51648 107188 51712
rect 107252 51648 107268 51712
rect 107332 51648 107338 51712
rect 107022 51647 107338 51648
rect 4870 51168 5186 51169
rect 4870 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5186 51168
rect 4870 51103 5186 51104
rect 107758 51168 108074 51169
rect 107758 51104 107764 51168
rect 107828 51104 107844 51168
rect 107908 51104 107924 51168
rect 107988 51104 108004 51168
rect 108068 51104 108074 51168
rect 107758 51103 108074 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 107022 50624 107338 50625
rect 107022 50560 107028 50624
rect 107092 50560 107108 50624
rect 107172 50560 107188 50624
rect 107252 50560 107268 50624
rect 107332 50560 107338 50624
rect 107022 50559 107338 50560
rect 4870 50080 5186 50081
rect 4870 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5186 50080
rect 4870 50015 5186 50016
rect 107758 50080 108074 50081
rect 107758 50016 107764 50080
rect 107828 50016 107844 50080
rect 107908 50016 107924 50080
rect 107988 50016 108004 50080
rect 108068 50016 108074 50080
rect 107758 50015 108074 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 107022 49536 107338 49537
rect 107022 49472 107028 49536
rect 107092 49472 107108 49536
rect 107172 49472 107188 49536
rect 107252 49472 107268 49536
rect 107332 49472 107338 49536
rect 107022 49471 107338 49472
rect 4870 48992 5186 48993
rect 4870 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5186 48992
rect 4870 48927 5186 48928
rect 107758 48992 108074 48993
rect 107758 48928 107764 48992
rect 107828 48928 107844 48992
rect 107908 48928 107924 48992
rect 107988 48928 108004 48992
rect 108068 48928 108074 48992
rect 107758 48927 108074 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 107022 48448 107338 48449
rect 107022 48384 107028 48448
rect 107092 48384 107108 48448
rect 107172 48384 107188 48448
rect 107252 48384 107268 48448
rect 107332 48384 107338 48448
rect 107022 48383 107338 48384
rect 4870 47904 5186 47905
rect 4870 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5186 47904
rect 4870 47839 5186 47840
rect 107758 47904 108074 47905
rect 107758 47840 107764 47904
rect 107828 47840 107844 47904
rect 107908 47840 107924 47904
rect 107988 47840 108004 47904
rect 108068 47840 108074 47904
rect 107758 47839 108074 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 107022 47360 107338 47361
rect 107022 47296 107028 47360
rect 107092 47296 107108 47360
rect 107172 47296 107188 47360
rect 107252 47296 107268 47360
rect 107332 47296 107338 47360
rect 107022 47295 107338 47296
rect 4870 46816 5186 46817
rect 4870 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5186 46816
rect 4870 46751 5186 46752
rect 107758 46816 108074 46817
rect 107758 46752 107764 46816
rect 107828 46752 107844 46816
rect 107908 46752 107924 46816
rect 107988 46752 108004 46816
rect 108068 46752 108074 46816
rect 107758 46751 108074 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 107022 46272 107338 46273
rect 107022 46208 107028 46272
rect 107092 46208 107108 46272
rect 107172 46208 107188 46272
rect 107252 46208 107268 46272
rect 107332 46208 107338 46272
rect 107022 46207 107338 46208
rect 4870 45728 5186 45729
rect 4870 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5186 45728
rect 4870 45663 5186 45664
rect 107758 45728 108074 45729
rect 107758 45664 107764 45728
rect 107828 45664 107844 45728
rect 107908 45664 107924 45728
rect 107988 45664 108004 45728
rect 108068 45664 108074 45728
rect 107758 45663 108074 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 107022 45184 107338 45185
rect 107022 45120 107028 45184
rect 107092 45120 107108 45184
rect 107172 45120 107188 45184
rect 107252 45120 107268 45184
rect 107332 45120 107338 45184
rect 107022 45119 107338 45120
rect 4870 44640 5186 44641
rect 4870 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5186 44640
rect 4870 44575 5186 44576
rect 107758 44640 108074 44641
rect 107758 44576 107764 44640
rect 107828 44576 107844 44640
rect 107908 44576 107924 44640
rect 107988 44576 108004 44640
rect 108068 44576 108074 44640
rect 107758 44575 108074 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 107022 44096 107338 44097
rect 107022 44032 107028 44096
rect 107092 44032 107108 44096
rect 107172 44032 107188 44096
rect 107252 44032 107268 44096
rect 107332 44032 107338 44096
rect 107022 44031 107338 44032
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 107758 43552 108074 43553
rect 107758 43488 107764 43552
rect 107828 43488 107844 43552
rect 107908 43488 107924 43552
rect 107988 43488 108004 43552
rect 108068 43488 108074 43552
rect 107758 43487 108074 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 107022 43008 107338 43009
rect 107022 42944 107028 43008
rect 107092 42944 107108 43008
rect 107172 42944 107188 43008
rect 107252 42944 107268 43008
rect 107332 42944 107338 43008
rect 107022 42943 107338 42944
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 107758 42464 108074 42465
rect 107758 42400 107764 42464
rect 107828 42400 107844 42464
rect 107908 42400 107924 42464
rect 107988 42400 108004 42464
rect 108068 42400 108074 42464
rect 107758 42399 108074 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 107022 41920 107338 41921
rect 107022 41856 107028 41920
rect 107092 41856 107108 41920
rect 107172 41856 107188 41920
rect 107252 41856 107268 41920
rect 107332 41856 107338 41920
rect 107022 41855 107338 41856
rect 0 41578 800 41608
rect 0 41518 6930 41578
rect 0 41488 800 41518
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 6870 41306 6930 41518
rect 107758 41376 108074 41377
rect 107758 41312 107764 41376
rect 107828 41312 107844 41376
rect 107908 41312 107924 41376
rect 107988 41312 108004 41376
rect 108068 41312 108074 41376
rect 107758 41311 108074 41312
rect 7557 41306 7623 41309
rect 6870 41304 9506 41306
rect 6870 41248 7562 41304
rect 7618 41254 9506 41304
rect 7618 41248 10028 41254
rect 6870 41246 10028 41248
rect 7557 41243 7623 41246
rect 9446 41194 10028 41246
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 107022 40832 107338 40833
rect 107022 40768 107028 40832
rect 107092 40768 107108 40832
rect 107172 40768 107188 40832
rect 107252 40768 107268 40832
rect 107332 40768 107338 40832
rect 107022 40767 107338 40768
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 107758 40288 108074 40289
rect 107758 40224 107764 40288
rect 107828 40224 107844 40288
rect 107908 40224 107924 40288
rect 107988 40224 108004 40288
rect 108068 40224 108074 40288
rect 107758 40223 108074 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 107022 39744 107338 39745
rect 107022 39680 107028 39744
rect 107092 39680 107108 39744
rect 107172 39680 107188 39744
rect 107252 39680 107268 39744
rect 107332 39680 107338 39744
rect 107022 39679 107338 39680
rect 0 39538 800 39568
rect 7557 39538 7623 39541
rect 9446 39538 10028 39554
rect 0 39536 10028 39538
rect 0 39480 7562 39536
rect 7618 39494 10028 39536
rect 7618 39480 9506 39494
rect 0 39478 9506 39480
rect 0 39448 800 39478
rect 7557 39475 7623 39478
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 107758 39200 108074 39201
rect 107758 39136 107764 39200
rect 107828 39136 107844 39200
rect 107908 39136 107924 39200
rect 107988 39136 108004 39200
rect 108068 39136 108074 39200
rect 107758 39135 108074 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 107022 38656 107338 38657
rect 107022 38592 107028 38656
rect 107092 38592 107108 38656
rect 107172 38592 107188 38656
rect 107252 38592 107268 38656
rect 107332 38592 107338 38656
rect 107022 38591 107338 38592
rect 9446 38366 10028 38426
rect 7557 38314 7623 38317
rect 9446 38314 9506 38366
rect 3006 38312 9506 38314
rect 3006 38256 7562 38312
rect 7618 38256 9506 38312
rect 3006 38254 9506 38256
rect 0 38178 800 38208
rect 3006 38178 3066 38254
rect 7557 38251 7623 38254
rect 0 38118 3066 38178
rect 0 38088 800 38118
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 107758 38112 108074 38113
rect 107758 38048 107764 38112
rect 107828 38048 107844 38112
rect 107908 38048 107924 38112
rect 107988 38048 108004 38112
rect 108068 38048 108074 38112
rect 107758 38047 108074 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 107022 37568 107338 37569
rect 107022 37504 107028 37568
rect 107092 37504 107108 37568
rect 107172 37504 107188 37568
rect 107252 37504 107268 37568
rect 107332 37504 107338 37568
rect 107022 37503 107338 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 107758 37024 108074 37025
rect 107758 36960 107764 37024
rect 107828 36960 107844 37024
rect 107908 36960 107924 37024
rect 107988 36960 108004 37024
rect 108068 36960 108074 37024
rect 107758 36959 108074 36960
rect 0 36818 800 36848
rect 7557 36818 7623 36821
rect 0 36816 9506 36818
rect 0 36760 7562 36816
rect 7618 36760 9506 36816
rect 0 36758 9506 36760
rect 0 36728 800 36758
rect 7557 36755 7623 36758
rect 9446 36726 9506 36758
rect 9446 36666 10028 36726
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 107022 36480 107338 36481
rect 107022 36416 107028 36480
rect 107092 36416 107108 36480
rect 107172 36416 107188 36480
rect 107252 36416 107268 36480
rect 107332 36416 107338 36480
rect 107022 36415 107338 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 107758 35936 108074 35937
rect 107758 35872 107764 35936
rect 107828 35872 107844 35936
rect 107908 35872 107924 35936
rect 107988 35872 108004 35936
rect 108068 35872 108074 35936
rect 107758 35871 108074 35872
rect 7557 35594 7623 35597
rect 9446 35594 10028 35643
rect 3374 35592 10028 35594
rect 3374 35536 7562 35592
rect 7618 35583 10028 35592
rect 7618 35536 9506 35583
rect 3374 35534 9506 35536
rect 0 35458 800 35488
rect 3374 35458 3434 35534
rect 7557 35531 7623 35534
rect 0 35398 3434 35458
rect 0 35368 800 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 107022 35392 107338 35393
rect 107022 35328 107028 35392
rect 107092 35328 107108 35392
rect 107172 35328 107188 35392
rect 107252 35328 107268 35392
rect 107332 35328 107338 35392
rect 107022 35327 107338 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 107758 34848 108074 34849
rect 107758 34784 107764 34848
rect 107828 34784 107844 34848
rect 107908 34784 107924 34848
rect 107988 34784 108004 34848
rect 108068 34784 108074 34848
rect 107758 34783 108074 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 107022 34304 107338 34305
rect 107022 34240 107028 34304
rect 107092 34240 107108 34304
rect 107172 34240 107188 34304
rect 107252 34240 107268 34304
rect 107332 34240 107338 34304
rect 107022 34239 107338 34240
rect 0 34098 800 34128
rect 7557 34098 7623 34101
rect 0 34096 9506 34098
rect 0 34040 7562 34096
rect 7618 34040 9506 34096
rect 0 34038 9506 34040
rect 0 34008 800 34038
rect 7557 34035 7623 34038
rect 9446 33963 9506 34038
rect 9446 33903 10028 33963
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 107758 33760 108074 33761
rect 107758 33696 107764 33760
rect 107828 33696 107844 33760
rect 107908 33696 107924 33760
rect 107988 33696 108004 33760
rect 108068 33696 108074 33760
rect 107758 33695 108074 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 107022 33216 107338 33217
rect 107022 33152 107028 33216
rect 107092 33152 107108 33216
rect 107172 33152 107188 33216
rect 107252 33152 107268 33216
rect 107332 33152 107338 33216
rect 107022 33151 107338 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 107758 32672 108074 32673
rect 107758 32608 107764 32672
rect 107828 32608 107844 32672
rect 107908 32608 107924 32672
rect 107988 32608 108004 32672
rect 108068 32608 108074 32672
rect 107758 32607 108074 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 107022 32128 107338 32129
rect 107022 32064 107028 32128
rect 107092 32064 107108 32128
rect 107172 32064 107188 32128
rect 107252 32064 107268 32128
rect 107332 32064 107338 32128
rect 107022 32063 107338 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 107758 31584 108074 31585
rect 107758 31520 107764 31584
rect 107828 31520 107844 31584
rect 107908 31520 107924 31584
rect 107988 31520 108004 31584
rect 108068 31520 108074 31584
rect 107758 31519 108074 31520
rect 110505 31378 110571 31381
rect 111200 31378 112000 31408
rect 110505 31376 112000 31378
rect 110505 31320 110510 31376
rect 110566 31320 112000 31376
rect 110505 31318 112000 31320
rect 110505 31315 110571 31318
rect 111200 31288 112000 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 107022 31040 107338 31041
rect 107022 30976 107028 31040
rect 107092 30976 107108 31040
rect 107172 30976 107188 31040
rect 107252 30976 107268 31040
rect 107332 30976 107338 31040
rect 107022 30975 107338 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 107758 30496 108074 30497
rect 107758 30432 107764 30496
rect 107828 30432 107844 30496
rect 107908 30432 107924 30496
rect 107988 30432 108004 30496
rect 108068 30432 108074 30496
rect 107758 30431 108074 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 107022 29952 107338 29953
rect 107022 29888 107028 29952
rect 107092 29888 107108 29952
rect 107172 29888 107188 29952
rect 107252 29888 107268 29952
rect 107332 29888 107338 29952
rect 107022 29887 107338 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 107758 29408 108074 29409
rect 107758 29344 107764 29408
rect 107828 29344 107844 29408
rect 107908 29344 107924 29408
rect 107988 29344 108004 29408
rect 108068 29344 108074 29408
rect 107758 29343 108074 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 107022 28864 107338 28865
rect 107022 28800 107028 28864
rect 107092 28800 107108 28864
rect 107172 28800 107188 28864
rect 107252 28800 107268 28864
rect 107332 28800 107338 28864
rect 107022 28799 107338 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 107758 28320 108074 28321
rect 107758 28256 107764 28320
rect 107828 28256 107844 28320
rect 107908 28256 107924 28320
rect 107988 28256 108004 28320
rect 108068 28256 108074 28320
rect 107758 28255 108074 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 107022 27776 107338 27777
rect 107022 27712 107028 27776
rect 107092 27712 107108 27776
rect 107172 27712 107188 27776
rect 107252 27712 107268 27776
rect 107332 27712 107338 27776
rect 107022 27711 107338 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 107758 27232 108074 27233
rect 107758 27168 107764 27232
rect 107828 27168 107844 27232
rect 107908 27168 107924 27232
rect 107988 27168 108004 27232
rect 108068 27168 108074 27232
rect 107758 27167 108074 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 107022 26688 107338 26689
rect 107022 26624 107028 26688
rect 107092 26624 107108 26688
rect 107172 26624 107188 26688
rect 107252 26624 107268 26688
rect 107332 26624 107338 26688
rect 107022 26623 107338 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 107758 26144 108074 26145
rect 107758 26080 107764 26144
rect 107828 26080 107844 26144
rect 107908 26080 107924 26144
rect 107988 26080 108004 26144
rect 108068 26080 108074 26144
rect 107758 26079 108074 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 107022 25600 107338 25601
rect 107022 25536 107028 25600
rect 107092 25536 107108 25600
rect 107172 25536 107188 25600
rect 107252 25536 107268 25600
rect 107332 25536 107338 25600
rect 107022 25535 107338 25536
rect 104157 25122 104223 25125
rect 102550 25120 104223 25122
rect 102550 25090 104162 25120
rect 101948 25064 104162 25090
rect 104218 25064 104223 25120
rect 101948 25062 104223 25064
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 101948 25030 102610 25062
rect 104157 25059 104223 25062
rect 107758 25056 108074 25057
rect 4870 24991 5186 24992
rect 107758 24992 107764 25056
rect 107828 24992 107844 25056
rect 107908 24992 107924 25056
rect 107988 24992 108004 25056
rect 108068 24992 108074 25056
rect 107758 24991 108074 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 107022 24512 107338 24513
rect 107022 24448 107028 24512
rect 107092 24448 107108 24512
rect 107172 24448 107188 24512
rect 107252 24448 107268 24512
rect 107332 24448 107338 24512
rect 107022 24447 107338 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 107758 23968 108074 23969
rect 107758 23904 107764 23968
rect 107828 23904 107844 23968
rect 107908 23904 107924 23968
rect 107988 23904 108004 23968
rect 108068 23904 108074 23968
rect 107758 23903 108074 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 107022 23424 107338 23425
rect 4210 23359 4526 23360
rect 101948 23354 102610 23390
rect 107022 23360 107028 23424
rect 107092 23360 107108 23424
rect 107172 23360 107188 23424
rect 107252 23360 107268 23424
rect 107332 23360 107338 23424
rect 107022 23359 107338 23360
rect 104341 23354 104407 23357
rect 101948 23352 104407 23354
rect 101948 23330 104346 23352
rect 102550 23296 104346 23330
rect 104402 23296 104407 23352
rect 102550 23294 104407 23296
rect 104341 23291 104407 23294
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 107758 22880 108074 22881
rect 107758 22816 107764 22880
rect 107828 22816 107844 22880
rect 107908 22816 107924 22880
rect 107988 22816 108004 22880
rect 108068 22816 108074 22880
rect 107758 22815 108074 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 107022 22336 107338 22337
rect 107022 22272 107028 22336
rect 107092 22272 107108 22336
rect 107172 22272 107188 22336
rect 107252 22272 107268 22336
rect 107332 22272 107338 22336
rect 107022 22271 107338 22272
rect 104525 22266 104591 22269
rect 102550 22264 104591 22266
rect 102550 22262 104530 22264
rect 101948 22208 104530 22262
rect 104586 22208 104591 22264
rect 101948 22206 104591 22208
rect 101948 22202 102610 22206
rect 104525 22203 104591 22206
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 107758 21792 108074 21793
rect 107758 21728 107764 21792
rect 107828 21728 107844 21792
rect 107908 21728 107924 21792
rect 107988 21728 108004 21792
rect 108068 21728 108074 21792
rect 107758 21727 108074 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 107022 21248 107338 21249
rect 107022 21184 107028 21248
rect 107092 21184 107108 21248
rect 107172 21184 107188 21248
rect 107252 21184 107268 21248
rect 107332 21184 107338 21248
rect 107022 21183 107338 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 107758 20704 108074 20705
rect 107758 20640 107764 20704
rect 107828 20640 107844 20704
rect 107908 20640 107924 20704
rect 107988 20640 108004 20704
rect 108068 20640 108074 20704
rect 107758 20639 108074 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 107022 20160 107338 20161
rect 107022 20096 107028 20160
rect 107092 20096 107108 20160
rect 107172 20096 107188 20160
rect 107252 20096 107268 20160
rect 107332 20096 107338 20160
rect 107022 20095 107338 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 107758 19616 108074 19617
rect 107758 19552 107764 19616
rect 107828 19552 107844 19616
rect 107908 19552 107924 19616
rect 107988 19552 108004 19616
rect 108068 19552 108074 19616
rect 107758 19551 108074 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 107022 19072 107338 19073
rect 107022 19008 107028 19072
rect 107092 19008 107108 19072
rect 107172 19008 107188 19072
rect 107252 19008 107268 19072
rect 107332 19008 107338 19072
rect 107022 19007 107338 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 107758 18528 108074 18529
rect 107758 18464 107764 18528
rect 107828 18464 107844 18528
rect 107908 18464 107924 18528
rect 107988 18464 108004 18528
rect 108068 18464 108074 18528
rect 107758 18463 108074 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 107022 17984 107338 17985
rect 107022 17920 107028 17984
rect 107092 17920 107108 17984
rect 107172 17920 107188 17984
rect 107252 17920 107268 17984
rect 107332 17920 107338 17984
rect 107022 17919 107338 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 107758 17440 108074 17441
rect 107758 17376 107764 17440
rect 107828 17376 107844 17440
rect 107908 17376 107924 17440
rect 107988 17376 108004 17440
rect 108068 17376 108074 17440
rect 107758 17375 108074 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 107022 16896 107338 16897
rect 107022 16832 107028 16896
rect 107092 16832 107108 16896
rect 107172 16832 107188 16896
rect 107252 16832 107268 16896
rect 107332 16832 107338 16896
rect 107022 16831 107338 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 107758 16352 108074 16353
rect 107758 16288 107764 16352
rect 107828 16288 107844 16352
rect 107908 16288 107924 16352
rect 107988 16288 108004 16352
rect 108068 16288 108074 16352
rect 107758 16287 108074 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 107022 15808 107338 15809
rect 107022 15744 107028 15808
rect 107092 15744 107108 15808
rect 107172 15744 107188 15808
rect 107252 15744 107268 15808
rect 107332 15744 107338 15808
rect 107022 15743 107338 15744
rect 0 15678 3434 15738
rect 0 15648 800 15678
rect 3374 15602 3434 15678
rect 7557 15602 7623 15605
rect 3374 15600 9506 15602
rect 3374 15544 7562 15600
rect 7618 15544 9506 15600
rect 3374 15542 9506 15544
rect 7557 15539 7623 15542
rect 9446 15483 9506 15542
rect 9446 15423 10028 15483
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 107758 15264 108074 15265
rect 107758 15200 107764 15264
rect 107828 15200 107844 15264
rect 107908 15200 107924 15264
rect 107988 15200 108004 15264
rect 108068 15200 108074 15264
rect 107758 15199 108074 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 107022 14720 107338 14721
rect 107022 14656 107028 14720
rect 107092 14656 107108 14720
rect 107172 14656 107188 14720
rect 107252 14656 107268 14720
rect 107332 14656 107338 14720
rect 107022 14655 107338 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 107758 14176 108074 14177
rect 107758 14112 107764 14176
rect 107828 14112 107844 14176
rect 107908 14112 107924 14176
rect 107988 14112 108004 14176
rect 108068 14112 108074 14176
rect 107758 14111 108074 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 107022 13632 107338 13633
rect 107022 13568 107028 13632
rect 107092 13568 107108 13632
rect 107172 13568 107188 13632
rect 107252 13568 107268 13632
rect 107332 13568 107338 13632
rect 107022 13567 107338 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 107758 13088 108074 13089
rect 107758 13024 107764 13088
rect 107828 13024 107844 13088
rect 107908 13024 107924 13088
rect 107988 13024 108004 13088
rect 108068 13024 108074 13088
rect 107758 13023 108074 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 107022 12544 107338 12545
rect 107022 12480 107028 12544
rect 107092 12480 107108 12544
rect 107172 12480 107188 12544
rect 107252 12480 107268 12544
rect 107332 12480 107338 12544
rect 107022 12479 107338 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 107758 12000 108074 12001
rect 107758 11936 107764 12000
rect 107828 11936 107844 12000
rect 107908 11936 107924 12000
rect 107988 11936 108004 12000
rect 108068 11936 108074 12000
rect 107758 11935 108074 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 107022 11456 107338 11457
rect 107022 11392 107028 11456
rect 107092 11392 107108 11456
rect 107172 11392 107188 11456
rect 107252 11392 107268 11456
rect 107332 11392 107338 11456
rect 107022 11391 107338 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 107758 10912 108074 10913
rect 107758 10848 107764 10912
rect 107828 10848 107844 10912
rect 107908 10848 107924 10912
rect 107988 10848 108004 10912
rect 108068 10848 108074 10912
rect 107758 10847 108074 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 107022 10368 107338 10369
rect 107022 10304 107028 10368
rect 107092 10304 107108 10368
rect 107172 10304 107188 10368
rect 107252 10304 107268 10368
rect 107332 10304 107338 10368
rect 107022 10303 107338 10304
rect 110413 10298 110479 10301
rect 111200 10298 112000 10328
rect 110413 10296 112000 10298
rect 110413 10240 110418 10296
rect 110474 10240 112000 10296
rect 110413 10238 112000 10240
rect 110413 10235 110479 10238
rect 111200 10208 112000 10238
rect 16021 9892 16087 9893
rect 90357 9892 90423 9893
rect 16021 9888 16058 9892
rect 16122 9890 16128 9892
rect 90357 9890 90404 9892
rect 16021 9832 16026 9888
rect 16021 9828 16058 9832
rect 16122 9830 16178 9890
rect 90312 9888 90404 9890
rect 90312 9832 90362 9888
rect 90312 9830 90404 9832
rect 16122 9828 16128 9830
rect 90357 9828 90404 9830
rect 90468 9828 90474 9892
rect 90950 9828 90956 9892
rect 91020 9890 91026 9892
rect 104249 9890 104315 9893
rect 91020 9888 104315 9890
rect 91020 9832 104254 9888
rect 104310 9832 104315 9888
rect 91020 9830 104315 9832
rect 91020 9828 91026 9830
rect 16021 9827 16087 9828
rect 90357 9827 90423 9828
rect 104249 9827 104315 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 107758 9824 108074 9825
rect 107758 9760 107764 9824
rect 107828 9760 107844 9824
rect 107908 9760 107924 9824
rect 107988 9760 108004 9824
rect 108068 9760 108074 9824
rect 107758 9759 108074 9760
rect 31569 9756 31635 9757
rect 31569 9754 31614 9756
rect 31522 9752 31614 9754
rect 31522 9696 31574 9752
rect 31522 9694 31614 9696
rect 31569 9692 31614 9694
rect 31678 9692 31684 9756
rect 31569 9691 31635 9692
rect 23473 9620 23539 9621
rect 30465 9620 30531 9621
rect 23432 9556 23438 9620
rect 23502 9618 23539 9620
rect 23502 9616 23594 9618
rect 23534 9560 23594 9616
rect 23502 9558 23594 9560
rect 23502 9556 23539 9558
rect 30440 9556 30446 9620
rect 30510 9618 30531 9620
rect 30510 9616 30602 9618
rect 30526 9560 30602 9616
rect 30510 9558 30602 9560
rect 30510 9556 30531 9558
rect 23473 9555 23539 9556
rect 30465 9555 30531 9556
rect 90725 9484 90791 9485
rect 90674 9482 90680 9484
rect 90634 9422 90680 9482
rect 90744 9480 90791 9484
rect 90786 9424 90791 9480
rect 90674 9420 90680 9422
rect 90744 9420 90791 9424
rect 90725 9419 90791 9420
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 107022 9280 107338 9281
rect 107022 9216 107028 9280
rect 107092 9216 107108 9280
rect 107172 9216 107188 9280
rect 107252 9216 107268 9280
rect 107332 9216 107338 9280
rect 107022 9215 107338 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 107758 8736 108074 8737
rect 107758 8672 107764 8736
rect 107828 8672 107844 8736
rect 107908 8672 107924 8736
rect 107988 8672 108004 8736
rect 108068 8672 108074 8736
rect 107758 8671 108074 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 107022 8192 107338 8193
rect 107022 8128 107028 8192
rect 107092 8128 107108 8192
rect 107172 8128 107188 8192
rect 107252 8128 107268 8192
rect 107332 8128 107338 8192
rect 107022 8127 107338 8128
rect 25773 8124 25839 8125
rect 25773 8122 25820 8124
rect 25728 8120 25820 8122
rect 25728 8064 25778 8120
rect 25728 8062 25820 8064
rect 25773 8060 25820 8062
rect 25884 8060 25890 8124
rect 28993 8122 29059 8125
rect 32857 8124 32923 8125
rect 35249 8124 35315 8125
rect 29310 8122 29316 8124
rect 28993 8120 29316 8122
rect 28993 8064 28998 8120
rect 29054 8064 29316 8120
rect 28993 8062 29316 8064
rect 25773 8059 25839 8060
rect 28993 8059 29059 8062
rect 29310 8060 29316 8062
rect 29380 8060 29386 8124
rect 32806 8060 32812 8124
rect 32876 8122 32923 8124
rect 32876 8120 32968 8122
rect 32918 8064 32968 8120
rect 32876 8062 32968 8064
rect 32876 8060 32923 8062
rect 35198 8060 35204 8124
rect 35268 8122 35315 8124
rect 38653 8124 38719 8125
rect 38653 8122 38700 8124
rect 35268 8120 35360 8122
rect 35310 8064 35360 8120
rect 35268 8062 35360 8064
rect 38608 8120 38700 8122
rect 38608 8064 38658 8120
rect 38608 8062 38700 8064
rect 35268 8060 35315 8062
rect 32857 8059 32923 8060
rect 35249 8059 35315 8060
rect 38653 8060 38700 8062
rect 38764 8060 38770 8124
rect 38653 8059 38719 8060
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 66310 7648 66626 7649
rect 66310 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66626 7648
rect 66310 7583 66626 7584
rect 97030 7648 97346 7649
rect 97030 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97346 7648
rect 97030 7583 97346 7584
rect 107758 7648 108074 7649
rect 107758 7584 107764 7648
rect 107828 7584 107844 7648
rect 107908 7584 107924 7648
rect 107988 7584 108004 7648
rect 108068 7584 108074 7648
rect 107758 7583 108074 7584
rect 24669 7580 24735 7581
rect 26969 7580 27035 7581
rect 28257 7580 28323 7581
rect 33961 7580 34027 7581
rect 36353 7580 36419 7581
rect 37457 7580 37523 7581
rect 39849 7580 39915 7581
rect 24669 7578 24716 7580
rect 24624 7576 24716 7578
rect 24624 7520 24674 7576
rect 24624 7518 24716 7520
rect 24669 7516 24716 7518
rect 24780 7516 24786 7580
rect 26918 7516 26924 7580
rect 26988 7578 27035 7580
rect 26988 7576 27080 7578
rect 27030 7520 27080 7576
rect 26988 7518 27080 7520
rect 26988 7516 27035 7518
rect 28206 7516 28212 7580
rect 28276 7578 28323 7580
rect 28276 7576 28368 7578
rect 28318 7520 28368 7576
rect 28276 7518 28368 7520
rect 28276 7516 28323 7518
rect 33910 7516 33916 7580
rect 33980 7578 34027 7580
rect 33980 7576 34072 7578
rect 34022 7520 34072 7576
rect 33980 7518 34072 7520
rect 33980 7516 34027 7518
rect 36302 7516 36308 7580
rect 36372 7578 36419 7580
rect 36372 7576 36464 7578
rect 36414 7520 36464 7576
rect 36372 7518 36464 7520
rect 36372 7516 36419 7518
rect 37406 7516 37412 7580
rect 37476 7578 37523 7580
rect 37476 7576 37568 7578
rect 37518 7520 37568 7576
rect 37476 7518 37568 7520
rect 37476 7516 37523 7518
rect 39798 7516 39804 7580
rect 39868 7578 39915 7580
rect 39868 7576 39960 7578
rect 39910 7520 39960 7576
rect 39868 7518 39960 7520
rect 39868 7516 39915 7518
rect 40902 7516 40908 7580
rect 40972 7578 40978 7580
rect 41045 7578 41111 7581
rect 42149 7580 42215 7581
rect 43345 7580 43411 7581
rect 42149 7578 42196 7580
rect 40972 7576 41111 7578
rect 40972 7520 41050 7576
rect 41106 7520 41111 7576
rect 40972 7518 41111 7520
rect 42104 7576 42196 7578
rect 42104 7520 42154 7576
rect 42104 7518 42196 7520
rect 40972 7516 40978 7518
rect 24669 7515 24735 7516
rect 26969 7515 27035 7516
rect 28257 7515 28323 7516
rect 33961 7515 34027 7516
rect 36353 7515 36419 7516
rect 37457 7515 37523 7516
rect 39849 7515 39915 7516
rect 41045 7515 41111 7518
rect 42149 7516 42196 7518
rect 42260 7516 42266 7580
rect 43294 7516 43300 7580
rect 43364 7578 43411 7580
rect 43364 7576 43456 7578
rect 43406 7520 43456 7576
rect 43364 7518 43456 7520
rect 43364 7516 43411 7518
rect 90398 7516 90404 7580
rect 90468 7578 90474 7580
rect 90541 7578 90607 7581
rect 91001 7580 91067 7581
rect 90468 7576 90607 7578
rect 90468 7520 90546 7576
rect 90602 7520 90607 7576
rect 90468 7518 90607 7520
rect 90468 7516 90474 7518
rect 42149 7515 42215 7516
rect 43345 7515 43411 7516
rect 90541 7515 90607 7518
rect 90950 7516 90956 7580
rect 91020 7578 91067 7580
rect 91020 7576 91112 7578
rect 91062 7520 91112 7576
rect 91020 7518 91112 7520
rect 91020 7516 91067 7518
rect 91001 7515 91067 7516
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 96370 7104 96686 7105
rect 96370 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96686 7104
rect 96370 7039 96686 7040
rect 107022 7104 107338 7105
rect 107022 7040 107028 7104
rect 107092 7040 107108 7104
rect 107172 7040 107188 7104
rect 107252 7040 107268 7104
rect 107332 7040 107338 7104
rect 107022 7039 107338 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 66310 6560 66626 6561
rect 66310 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66626 6560
rect 66310 6495 66626 6496
rect 97030 6560 97346 6561
rect 97030 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97346 6560
rect 97030 6495 97346 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 96370 6016 96686 6017
rect 96370 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96686 6016
rect 96370 5951 96686 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 66310 5472 66626 5473
rect 66310 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66626 5472
rect 66310 5407 66626 5408
rect 97030 5472 97346 5473
rect 97030 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97346 5472
rect 97030 5407 97346 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 96370 4928 96686 4929
rect 96370 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96686 4928
rect 96370 4863 96686 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 66310 4384 66626 4385
rect 66310 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66626 4384
rect 66310 4319 66626 4320
rect 97030 4384 97346 4385
rect 97030 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97346 4384
rect 97030 4319 97346 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 96370 3840 96686 3841
rect 96370 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96686 3840
rect 96370 3775 96686 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 66310 3296 66626 3297
rect 66310 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66626 3296
rect 66310 3231 66626 3232
rect 97030 3296 97346 3297
rect 97030 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97346 3296
rect 97030 3231 97346 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 96370 2752 96686 2753
rect 96370 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96686 2752
rect 96370 2687 96686 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 66310 2208 66626 2209
rect 66310 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66626 2208
rect 66310 2143 66626 2144
rect 97030 2208 97346 2209
rect 97030 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97346 2208
rect 97030 2143 97346 2144
<< via3 >>
rect 4876 71836 4940 71840
rect 4876 71780 4880 71836
rect 4880 71780 4936 71836
rect 4936 71780 4940 71836
rect 4876 71776 4940 71780
rect 4956 71836 5020 71840
rect 4956 71780 4960 71836
rect 4960 71780 5016 71836
rect 5016 71780 5020 71836
rect 4956 71776 5020 71780
rect 5036 71836 5100 71840
rect 5036 71780 5040 71836
rect 5040 71780 5096 71836
rect 5096 71780 5100 71836
rect 5036 71776 5100 71780
rect 5116 71836 5180 71840
rect 5116 71780 5120 71836
rect 5120 71780 5176 71836
rect 5176 71780 5180 71836
rect 5116 71776 5180 71780
rect 35596 71836 35660 71840
rect 35596 71780 35600 71836
rect 35600 71780 35656 71836
rect 35656 71780 35660 71836
rect 35596 71776 35660 71780
rect 35676 71836 35740 71840
rect 35676 71780 35680 71836
rect 35680 71780 35736 71836
rect 35736 71780 35740 71836
rect 35676 71776 35740 71780
rect 35756 71836 35820 71840
rect 35756 71780 35760 71836
rect 35760 71780 35816 71836
rect 35816 71780 35820 71836
rect 35756 71776 35820 71780
rect 35836 71836 35900 71840
rect 35836 71780 35840 71836
rect 35840 71780 35896 71836
rect 35896 71780 35900 71836
rect 35836 71776 35900 71780
rect 66316 71836 66380 71840
rect 66316 71780 66320 71836
rect 66320 71780 66376 71836
rect 66376 71780 66380 71836
rect 66316 71776 66380 71780
rect 66396 71836 66460 71840
rect 66396 71780 66400 71836
rect 66400 71780 66456 71836
rect 66456 71780 66460 71836
rect 66396 71776 66460 71780
rect 66476 71836 66540 71840
rect 66476 71780 66480 71836
rect 66480 71780 66536 71836
rect 66536 71780 66540 71836
rect 66476 71776 66540 71780
rect 66556 71836 66620 71840
rect 66556 71780 66560 71836
rect 66560 71780 66616 71836
rect 66616 71780 66620 71836
rect 66556 71776 66620 71780
rect 97036 71836 97100 71840
rect 97036 71780 97040 71836
rect 97040 71780 97096 71836
rect 97096 71780 97100 71836
rect 97036 71776 97100 71780
rect 97116 71836 97180 71840
rect 97116 71780 97120 71836
rect 97120 71780 97176 71836
rect 97176 71780 97180 71836
rect 97116 71776 97180 71780
rect 97196 71836 97260 71840
rect 97196 71780 97200 71836
rect 97200 71780 97256 71836
rect 97256 71780 97260 71836
rect 97196 71776 97260 71780
rect 97276 71836 97340 71840
rect 97276 71780 97280 71836
rect 97280 71780 97336 71836
rect 97336 71780 97340 71836
rect 97276 71776 97340 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 34936 71292 35000 71296
rect 34936 71236 34940 71292
rect 34940 71236 34996 71292
rect 34996 71236 35000 71292
rect 34936 71232 35000 71236
rect 35016 71292 35080 71296
rect 35016 71236 35020 71292
rect 35020 71236 35076 71292
rect 35076 71236 35080 71292
rect 35016 71232 35080 71236
rect 35096 71292 35160 71296
rect 35096 71236 35100 71292
rect 35100 71236 35156 71292
rect 35156 71236 35160 71292
rect 35096 71232 35160 71236
rect 35176 71292 35240 71296
rect 35176 71236 35180 71292
rect 35180 71236 35236 71292
rect 35236 71236 35240 71292
rect 35176 71232 35240 71236
rect 65656 71292 65720 71296
rect 65656 71236 65660 71292
rect 65660 71236 65716 71292
rect 65716 71236 65720 71292
rect 65656 71232 65720 71236
rect 65736 71292 65800 71296
rect 65736 71236 65740 71292
rect 65740 71236 65796 71292
rect 65796 71236 65800 71292
rect 65736 71232 65800 71236
rect 65816 71292 65880 71296
rect 65816 71236 65820 71292
rect 65820 71236 65876 71292
rect 65876 71236 65880 71292
rect 65816 71232 65880 71236
rect 65896 71292 65960 71296
rect 65896 71236 65900 71292
rect 65900 71236 65956 71292
rect 65956 71236 65960 71292
rect 65896 71232 65960 71236
rect 96376 71292 96440 71296
rect 96376 71236 96380 71292
rect 96380 71236 96436 71292
rect 96436 71236 96440 71292
rect 96376 71232 96440 71236
rect 96456 71292 96520 71296
rect 96456 71236 96460 71292
rect 96460 71236 96516 71292
rect 96516 71236 96520 71292
rect 96456 71232 96520 71236
rect 96536 71292 96600 71296
rect 96536 71236 96540 71292
rect 96540 71236 96596 71292
rect 96596 71236 96600 71292
rect 96536 71232 96600 71236
rect 96616 71292 96680 71296
rect 96616 71236 96620 71292
rect 96620 71236 96676 71292
rect 96676 71236 96680 71292
rect 96616 71232 96680 71236
rect 4876 70748 4940 70752
rect 4876 70692 4880 70748
rect 4880 70692 4936 70748
rect 4936 70692 4940 70748
rect 4876 70688 4940 70692
rect 4956 70748 5020 70752
rect 4956 70692 4960 70748
rect 4960 70692 5016 70748
rect 5016 70692 5020 70748
rect 4956 70688 5020 70692
rect 5036 70748 5100 70752
rect 5036 70692 5040 70748
rect 5040 70692 5096 70748
rect 5096 70692 5100 70748
rect 5036 70688 5100 70692
rect 5116 70748 5180 70752
rect 5116 70692 5120 70748
rect 5120 70692 5176 70748
rect 5176 70692 5180 70748
rect 5116 70688 5180 70692
rect 35596 70748 35660 70752
rect 35596 70692 35600 70748
rect 35600 70692 35656 70748
rect 35656 70692 35660 70748
rect 35596 70688 35660 70692
rect 35676 70748 35740 70752
rect 35676 70692 35680 70748
rect 35680 70692 35736 70748
rect 35736 70692 35740 70748
rect 35676 70688 35740 70692
rect 35756 70748 35820 70752
rect 35756 70692 35760 70748
rect 35760 70692 35816 70748
rect 35816 70692 35820 70748
rect 35756 70688 35820 70692
rect 35836 70748 35900 70752
rect 35836 70692 35840 70748
rect 35840 70692 35896 70748
rect 35896 70692 35900 70748
rect 35836 70688 35900 70692
rect 66316 70748 66380 70752
rect 66316 70692 66320 70748
rect 66320 70692 66376 70748
rect 66376 70692 66380 70748
rect 66316 70688 66380 70692
rect 66396 70748 66460 70752
rect 66396 70692 66400 70748
rect 66400 70692 66456 70748
rect 66456 70692 66460 70748
rect 66396 70688 66460 70692
rect 66476 70748 66540 70752
rect 66476 70692 66480 70748
rect 66480 70692 66536 70748
rect 66536 70692 66540 70748
rect 66476 70688 66540 70692
rect 66556 70748 66620 70752
rect 66556 70692 66560 70748
rect 66560 70692 66616 70748
rect 66616 70692 66620 70748
rect 66556 70688 66620 70692
rect 97036 70748 97100 70752
rect 97036 70692 97040 70748
rect 97040 70692 97096 70748
rect 97096 70692 97100 70748
rect 97036 70688 97100 70692
rect 97116 70748 97180 70752
rect 97116 70692 97120 70748
rect 97120 70692 97176 70748
rect 97176 70692 97180 70748
rect 97116 70688 97180 70692
rect 97196 70748 97260 70752
rect 97196 70692 97200 70748
rect 97200 70692 97256 70748
rect 97256 70692 97260 70748
rect 97196 70688 97260 70692
rect 97276 70748 97340 70752
rect 97276 70692 97280 70748
rect 97280 70692 97336 70748
rect 97336 70692 97340 70748
rect 97276 70688 97340 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 34936 70204 35000 70208
rect 34936 70148 34940 70204
rect 34940 70148 34996 70204
rect 34996 70148 35000 70204
rect 34936 70144 35000 70148
rect 35016 70204 35080 70208
rect 35016 70148 35020 70204
rect 35020 70148 35076 70204
rect 35076 70148 35080 70204
rect 35016 70144 35080 70148
rect 35096 70204 35160 70208
rect 35096 70148 35100 70204
rect 35100 70148 35156 70204
rect 35156 70148 35160 70204
rect 35096 70144 35160 70148
rect 35176 70204 35240 70208
rect 35176 70148 35180 70204
rect 35180 70148 35236 70204
rect 35236 70148 35240 70204
rect 35176 70144 35240 70148
rect 65656 70204 65720 70208
rect 65656 70148 65660 70204
rect 65660 70148 65716 70204
rect 65716 70148 65720 70204
rect 65656 70144 65720 70148
rect 65736 70204 65800 70208
rect 65736 70148 65740 70204
rect 65740 70148 65796 70204
rect 65796 70148 65800 70204
rect 65736 70144 65800 70148
rect 65816 70204 65880 70208
rect 65816 70148 65820 70204
rect 65820 70148 65876 70204
rect 65876 70148 65880 70204
rect 65816 70144 65880 70148
rect 65896 70204 65960 70208
rect 65896 70148 65900 70204
rect 65900 70148 65956 70204
rect 65956 70148 65960 70204
rect 65896 70144 65960 70148
rect 96376 70204 96440 70208
rect 96376 70148 96380 70204
rect 96380 70148 96436 70204
rect 96436 70148 96440 70204
rect 96376 70144 96440 70148
rect 96456 70204 96520 70208
rect 96456 70148 96460 70204
rect 96460 70148 96516 70204
rect 96516 70148 96520 70204
rect 96456 70144 96520 70148
rect 96536 70204 96600 70208
rect 96536 70148 96540 70204
rect 96540 70148 96596 70204
rect 96596 70148 96600 70204
rect 96536 70144 96600 70148
rect 96616 70204 96680 70208
rect 96616 70148 96620 70204
rect 96620 70148 96676 70204
rect 96676 70148 96680 70204
rect 96616 70144 96680 70148
rect 4876 69660 4940 69664
rect 4876 69604 4880 69660
rect 4880 69604 4936 69660
rect 4936 69604 4940 69660
rect 4876 69600 4940 69604
rect 4956 69660 5020 69664
rect 4956 69604 4960 69660
rect 4960 69604 5016 69660
rect 5016 69604 5020 69660
rect 4956 69600 5020 69604
rect 5036 69660 5100 69664
rect 5036 69604 5040 69660
rect 5040 69604 5096 69660
rect 5096 69604 5100 69660
rect 5036 69600 5100 69604
rect 5116 69660 5180 69664
rect 5116 69604 5120 69660
rect 5120 69604 5176 69660
rect 5176 69604 5180 69660
rect 5116 69600 5180 69604
rect 35596 69660 35660 69664
rect 35596 69604 35600 69660
rect 35600 69604 35656 69660
rect 35656 69604 35660 69660
rect 35596 69600 35660 69604
rect 35676 69660 35740 69664
rect 35676 69604 35680 69660
rect 35680 69604 35736 69660
rect 35736 69604 35740 69660
rect 35676 69600 35740 69604
rect 35756 69660 35820 69664
rect 35756 69604 35760 69660
rect 35760 69604 35816 69660
rect 35816 69604 35820 69660
rect 35756 69600 35820 69604
rect 35836 69660 35900 69664
rect 35836 69604 35840 69660
rect 35840 69604 35896 69660
rect 35896 69604 35900 69660
rect 35836 69600 35900 69604
rect 66316 69660 66380 69664
rect 66316 69604 66320 69660
rect 66320 69604 66376 69660
rect 66376 69604 66380 69660
rect 66316 69600 66380 69604
rect 66396 69660 66460 69664
rect 66396 69604 66400 69660
rect 66400 69604 66456 69660
rect 66456 69604 66460 69660
rect 66396 69600 66460 69604
rect 66476 69660 66540 69664
rect 66476 69604 66480 69660
rect 66480 69604 66536 69660
rect 66536 69604 66540 69660
rect 66476 69600 66540 69604
rect 66556 69660 66620 69664
rect 66556 69604 66560 69660
rect 66560 69604 66616 69660
rect 66616 69604 66620 69660
rect 66556 69600 66620 69604
rect 97036 69660 97100 69664
rect 97036 69604 97040 69660
rect 97040 69604 97096 69660
rect 97096 69604 97100 69660
rect 97036 69600 97100 69604
rect 97116 69660 97180 69664
rect 97116 69604 97120 69660
rect 97120 69604 97176 69660
rect 97176 69604 97180 69660
rect 97116 69600 97180 69604
rect 97196 69660 97260 69664
rect 97196 69604 97200 69660
rect 97200 69604 97256 69660
rect 97256 69604 97260 69660
rect 97196 69600 97260 69604
rect 97276 69660 97340 69664
rect 97276 69604 97280 69660
rect 97280 69604 97336 69660
rect 97336 69604 97340 69660
rect 97276 69600 97340 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 96376 69116 96440 69120
rect 96376 69060 96380 69116
rect 96380 69060 96436 69116
rect 96436 69060 96440 69116
rect 96376 69056 96440 69060
rect 96456 69116 96520 69120
rect 96456 69060 96460 69116
rect 96460 69060 96516 69116
rect 96516 69060 96520 69116
rect 96456 69056 96520 69060
rect 96536 69116 96600 69120
rect 96536 69060 96540 69116
rect 96540 69060 96596 69116
rect 96596 69060 96600 69116
rect 96536 69056 96600 69060
rect 96616 69116 96680 69120
rect 96616 69060 96620 69116
rect 96620 69060 96676 69116
rect 96676 69060 96680 69116
rect 96616 69056 96680 69060
rect 4876 68572 4940 68576
rect 4876 68516 4880 68572
rect 4880 68516 4936 68572
rect 4936 68516 4940 68572
rect 4876 68512 4940 68516
rect 4956 68572 5020 68576
rect 4956 68516 4960 68572
rect 4960 68516 5016 68572
rect 5016 68516 5020 68572
rect 4956 68512 5020 68516
rect 5036 68572 5100 68576
rect 5036 68516 5040 68572
rect 5040 68516 5096 68572
rect 5096 68516 5100 68572
rect 5036 68512 5100 68516
rect 5116 68572 5180 68576
rect 5116 68516 5120 68572
rect 5120 68516 5176 68572
rect 5176 68516 5180 68572
rect 5116 68512 5180 68516
rect 35596 68572 35660 68576
rect 35596 68516 35600 68572
rect 35600 68516 35656 68572
rect 35656 68516 35660 68572
rect 35596 68512 35660 68516
rect 35676 68572 35740 68576
rect 35676 68516 35680 68572
rect 35680 68516 35736 68572
rect 35736 68516 35740 68572
rect 35676 68512 35740 68516
rect 35756 68572 35820 68576
rect 35756 68516 35760 68572
rect 35760 68516 35816 68572
rect 35816 68516 35820 68572
rect 35756 68512 35820 68516
rect 35836 68572 35900 68576
rect 35836 68516 35840 68572
rect 35840 68516 35896 68572
rect 35896 68516 35900 68572
rect 35836 68512 35900 68516
rect 66316 68572 66380 68576
rect 66316 68516 66320 68572
rect 66320 68516 66376 68572
rect 66376 68516 66380 68572
rect 66316 68512 66380 68516
rect 66396 68572 66460 68576
rect 66396 68516 66400 68572
rect 66400 68516 66456 68572
rect 66456 68516 66460 68572
rect 66396 68512 66460 68516
rect 66476 68572 66540 68576
rect 66476 68516 66480 68572
rect 66480 68516 66536 68572
rect 66536 68516 66540 68572
rect 66476 68512 66540 68516
rect 66556 68572 66620 68576
rect 66556 68516 66560 68572
rect 66560 68516 66616 68572
rect 66616 68516 66620 68572
rect 66556 68512 66620 68516
rect 97036 68572 97100 68576
rect 97036 68516 97040 68572
rect 97040 68516 97096 68572
rect 97096 68516 97100 68572
rect 97036 68512 97100 68516
rect 97116 68572 97180 68576
rect 97116 68516 97120 68572
rect 97120 68516 97176 68572
rect 97176 68516 97180 68572
rect 97116 68512 97180 68516
rect 97196 68572 97260 68576
rect 97196 68516 97200 68572
rect 97200 68516 97256 68572
rect 97256 68516 97260 68572
rect 97196 68512 97260 68516
rect 97276 68572 97340 68576
rect 97276 68516 97280 68572
rect 97280 68516 97336 68572
rect 97336 68516 97340 68572
rect 97276 68512 97340 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 96376 68028 96440 68032
rect 96376 67972 96380 68028
rect 96380 67972 96436 68028
rect 96436 67972 96440 68028
rect 96376 67968 96440 67972
rect 96456 68028 96520 68032
rect 96456 67972 96460 68028
rect 96460 67972 96516 68028
rect 96516 67972 96520 68028
rect 96456 67968 96520 67972
rect 96536 68028 96600 68032
rect 96536 67972 96540 68028
rect 96540 67972 96596 68028
rect 96596 67972 96600 68028
rect 96536 67968 96600 67972
rect 96616 68028 96680 68032
rect 96616 67972 96620 68028
rect 96620 67972 96676 68028
rect 96676 67972 96680 68028
rect 96616 67968 96680 67972
rect 4876 67484 4940 67488
rect 4876 67428 4880 67484
rect 4880 67428 4936 67484
rect 4936 67428 4940 67484
rect 4876 67424 4940 67428
rect 4956 67484 5020 67488
rect 4956 67428 4960 67484
rect 4960 67428 5016 67484
rect 5016 67428 5020 67484
rect 4956 67424 5020 67428
rect 5036 67484 5100 67488
rect 5036 67428 5040 67484
rect 5040 67428 5096 67484
rect 5096 67428 5100 67484
rect 5036 67424 5100 67428
rect 5116 67484 5180 67488
rect 5116 67428 5120 67484
rect 5120 67428 5176 67484
rect 5176 67428 5180 67484
rect 5116 67424 5180 67428
rect 35596 67484 35660 67488
rect 35596 67428 35600 67484
rect 35600 67428 35656 67484
rect 35656 67428 35660 67484
rect 35596 67424 35660 67428
rect 35676 67484 35740 67488
rect 35676 67428 35680 67484
rect 35680 67428 35736 67484
rect 35736 67428 35740 67484
rect 35676 67424 35740 67428
rect 35756 67484 35820 67488
rect 35756 67428 35760 67484
rect 35760 67428 35816 67484
rect 35816 67428 35820 67484
rect 35756 67424 35820 67428
rect 35836 67484 35900 67488
rect 35836 67428 35840 67484
rect 35840 67428 35896 67484
rect 35896 67428 35900 67484
rect 35836 67424 35900 67428
rect 66316 67484 66380 67488
rect 66316 67428 66320 67484
rect 66320 67428 66376 67484
rect 66376 67428 66380 67484
rect 66316 67424 66380 67428
rect 66396 67484 66460 67488
rect 66396 67428 66400 67484
rect 66400 67428 66456 67484
rect 66456 67428 66460 67484
rect 66396 67424 66460 67428
rect 66476 67484 66540 67488
rect 66476 67428 66480 67484
rect 66480 67428 66536 67484
rect 66536 67428 66540 67484
rect 66476 67424 66540 67428
rect 66556 67484 66620 67488
rect 66556 67428 66560 67484
rect 66560 67428 66616 67484
rect 66616 67428 66620 67484
rect 66556 67424 66620 67428
rect 97036 67484 97100 67488
rect 97036 67428 97040 67484
rect 97040 67428 97096 67484
rect 97096 67428 97100 67484
rect 97036 67424 97100 67428
rect 97116 67484 97180 67488
rect 97116 67428 97120 67484
rect 97120 67428 97176 67484
rect 97176 67428 97180 67484
rect 97116 67424 97180 67428
rect 97196 67484 97260 67488
rect 97196 67428 97200 67484
rect 97200 67428 97256 67484
rect 97256 67428 97260 67484
rect 97196 67424 97260 67428
rect 97276 67484 97340 67488
rect 97276 67428 97280 67484
rect 97280 67428 97336 67484
rect 97336 67428 97340 67484
rect 97276 67424 97340 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 96376 66940 96440 66944
rect 96376 66884 96380 66940
rect 96380 66884 96436 66940
rect 96436 66884 96440 66940
rect 96376 66880 96440 66884
rect 96456 66940 96520 66944
rect 96456 66884 96460 66940
rect 96460 66884 96516 66940
rect 96516 66884 96520 66940
rect 96456 66880 96520 66884
rect 96536 66940 96600 66944
rect 96536 66884 96540 66940
rect 96540 66884 96596 66940
rect 96596 66884 96600 66940
rect 96536 66880 96600 66884
rect 96616 66940 96680 66944
rect 96616 66884 96620 66940
rect 96620 66884 96676 66940
rect 96676 66884 96680 66940
rect 96616 66880 96680 66884
rect 51028 66676 51092 66740
rect 66116 66540 66180 66604
rect 48636 66404 48700 66468
rect 55996 66404 56060 66468
rect 61148 66404 61212 66468
rect 4876 66396 4940 66400
rect 4876 66340 4880 66396
rect 4880 66340 4936 66396
rect 4936 66340 4940 66396
rect 4876 66336 4940 66340
rect 4956 66396 5020 66400
rect 4956 66340 4960 66396
rect 4960 66340 5016 66396
rect 5016 66340 5020 66396
rect 4956 66336 5020 66340
rect 5036 66396 5100 66400
rect 5036 66340 5040 66396
rect 5040 66340 5096 66396
rect 5096 66340 5100 66396
rect 5036 66336 5100 66340
rect 5116 66396 5180 66400
rect 5116 66340 5120 66396
rect 5120 66340 5176 66396
rect 5176 66340 5180 66396
rect 5116 66336 5180 66340
rect 35596 66396 35660 66400
rect 35596 66340 35600 66396
rect 35600 66340 35656 66396
rect 35656 66340 35660 66396
rect 35596 66336 35660 66340
rect 35676 66396 35740 66400
rect 35676 66340 35680 66396
rect 35680 66340 35736 66396
rect 35736 66340 35740 66396
rect 35676 66336 35740 66340
rect 35756 66396 35820 66400
rect 35756 66340 35760 66396
rect 35760 66340 35816 66396
rect 35816 66340 35820 66396
rect 35756 66336 35820 66340
rect 35836 66396 35900 66400
rect 35836 66340 35840 66396
rect 35840 66340 35896 66396
rect 35896 66340 35900 66396
rect 35836 66336 35900 66340
rect 66316 66396 66380 66400
rect 66316 66340 66320 66396
rect 66320 66340 66376 66396
rect 66376 66340 66380 66396
rect 66316 66336 66380 66340
rect 66396 66396 66460 66400
rect 66396 66340 66400 66396
rect 66400 66340 66456 66396
rect 66456 66340 66460 66396
rect 66396 66336 66460 66340
rect 66476 66396 66540 66400
rect 66476 66340 66480 66396
rect 66480 66340 66536 66396
rect 66536 66340 66540 66396
rect 66476 66336 66540 66340
rect 66556 66396 66620 66400
rect 66556 66340 66560 66396
rect 66560 66340 66616 66396
rect 66616 66340 66620 66396
rect 66556 66336 66620 66340
rect 97036 66396 97100 66400
rect 97036 66340 97040 66396
rect 97040 66340 97096 66396
rect 97096 66340 97100 66396
rect 97036 66336 97100 66340
rect 97116 66396 97180 66400
rect 97116 66340 97120 66396
rect 97120 66340 97176 66396
rect 97176 66340 97180 66396
rect 97116 66336 97180 66340
rect 97196 66396 97260 66400
rect 97196 66340 97200 66396
rect 97200 66340 97256 66396
rect 97256 66340 97260 66396
rect 97196 66336 97260 66340
rect 97276 66396 97340 66400
rect 97276 66340 97280 66396
rect 97280 66340 97336 66396
rect 97336 66340 97340 66396
rect 97276 66336 97340 66340
rect 107764 66396 107828 66400
rect 107764 66340 107768 66396
rect 107768 66340 107824 66396
rect 107824 66340 107828 66396
rect 107764 66336 107828 66340
rect 107844 66396 107908 66400
rect 107844 66340 107848 66396
rect 107848 66340 107904 66396
rect 107904 66340 107908 66396
rect 107844 66336 107908 66340
rect 107924 66396 107988 66400
rect 107924 66340 107928 66396
rect 107928 66340 107984 66396
rect 107984 66340 107988 66396
rect 107924 66336 107988 66340
rect 108004 66396 108068 66400
rect 108004 66340 108008 66396
rect 108008 66340 108064 66396
rect 108064 66340 108068 66396
rect 108004 66336 108068 66340
rect 46060 66268 46124 66332
rect 58572 66268 58636 66332
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 96376 65852 96440 65856
rect 96376 65796 96380 65852
rect 96380 65796 96436 65852
rect 96436 65796 96440 65852
rect 96376 65792 96440 65796
rect 96456 65852 96520 65856
rect 96456 65796 96460 65852
rect 96460 65796 96516 65852
rect 96516 65796 96520 65852
rect 96456 65792 96520 65796
rect 96536 65852 96600 65856
rect 96536 65796 96540 65852
rect 96540 65796 96596 65852
rect 96596 65796 96600 65852
rect 96536 65792 96600 65796
rect 96616 65852 96680 65856
rect 96616 65796 96620 65852
rect 96620 65796 96676 65852
rect 96676 65796 96680 65852
rect 96616 65792 96680 65796
rect 107028 65852 107092 65856
rect 107028 65796 107032 65852
rect 107032 65796 107088 65852
rect 107088 65796 107092 65852
rect 107028 65792 107092 65796
rect 107108 65852 107172 65856
rect 107108 65796 107112 65852
rect 107112 65796 107168 65852
rect 107168 65796 107172 65852
rect 107108 65792 107172 65796
rect 107188 65852 107252 65856
rect 107188 65796 107192 65852
rect 107192 65796 107248 65852
rect 107248 65796 107252 65852
rect 107188 65792 107252 65796
rect 107268 65852 107332 65856
rect 107268 65796 107272 65852
rect 107272 65796 107328 65852
rect 107328 65796 107332 65852
rect 107268 65792 107332 65796
rect 63540 65452 63604 65516
rect 68508 65316 68572 65380
rect 73476 65316 73540 65380
rect 87276 65376 87340 65380
rect 87276 65320 87326 65376
rect 87326 65320 87340 65376
rect 87276 65316 87340 65320
rect 4876 65308 4940 65312
rect 4876 65252 4880 65308
rect 4880 65252 4936 65308
rect 4936 65252 4940 65308
rect 4876 65248 4940 65252
rect 4956 65308 5020 65312
rect 4956 65252 4960 65308
rect 4960 65252 5016 65308
rect 5016 65252 5020 65308
rect 4956 65248 5020 65252
rect 5036 65308 5100 65312
rect 5036 65252 5040 65308
rect 5040 65252 5096 65308
rect 5096 65252 5100 65308
rect 5036 65248 5100 65252
rect 5116 65308 5180 65312
rect 5116 65252 5120 65308
rect 5120 65252 5176 65308
rect 5176 65252 5180 65308
rect 5116 65248 5180 65252
rect 107764 65308 107828 65312
rect 107764 65252 107768 65308
rect 107768 65252 107824 65308
rect 107824 65252 107828 65308
rect 107764 65248 107828 65252
rect 107844 65308 107908 65312
rect 107844 65252 107848 65308
rect 107848 65252 107904 65308
rect 107904 65252 107908 65308
rect 107844 65248 107908 65252
rect 107924 65308 107988 65312
rect 107924 65252 107928 65308
rect 107928 65252 107984 65308
rect 107984 65252 107988 65308
rect 107924 65248 107988 65252
rect 108004 65308 108068 65312
rect 108004 65252 108008 65308
rect 108008 65252 108064 65308
rect 108064 65252 108068 65308
rect 108004 65248 108068 65252
rect 71084 65044 71148 65108
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 107028 64764 107092 64768
rect 107028 64708 107032 64764
rect 107032 64708 107088 64764
rect 107088 64708 107092 64764
rect 107028 64704 107092 64708
rect 107108 64764 107172 64768
rect 107108 64708 107112 64764
rect 107112 64708 107168 64764
rect 107168 64708 107172 64764
rect 107108 64704 107172 64708
rect 107188 64764 107252 64768
rect 107188 64708 107192 64764
rect 107192 64708 107248 64764
rect 107248 64708 107252 64764
rect 107188 64704 107252 64708
rect 107268 64764 107332 64768
rect 107268 64708 107272 64764
rect 107272 64708 107328 64764
rect 107328 64708 107332 64764
rect 107268 64704 107332 64708
rect 4876 64220 4940 64224
rect 4876 64164 4880 64220
rect 4880 64164 4936 64220
rect 4936 64164 4940 64220
rect 4876 64160 4940 64164
rect 4956 64220 5020 64224
rect 4956 64164 4960 64220
rect 4960 64164 5016 64220
rect 5016 64164 5020 64220
rect 4956 64160 5020 64164
rect 5036 64220 5100 64224
rect 5036 64164 5040 64220
rect 5040 64164 5096 64220
rect 5096 64164 5100 64220
rect 5036 64160 5100 64164
rect 5116 64220 5180 64224
rect 5116 64164 5120 64220
rect 5120 64164 5176 64220
rect 5176 64164 5180 64220
rect 5116 64160 5180 64164
rect 107764 64220 107828 64224
rect 107764 64164 107768 64220
rect 107768 64164 107824 64220
rect 107824 64164 107828 64220
rect 107764 64160 107828 64164
rect 107844 64220 107908 64224
rect 107844 64164 107848 64220
rect 107848 64164 107904 64220
rect 107904 64164 107908 64220
rect 107844 64160 107908 64164
rect 107924 64220 107988 64224
rect 107924 64164 107928 64220
rect 107928 64164 107984 64220
rect 107984 64164 107988 64220
rect 107924 64160 107988 64164
rect 108004 64220 108068 64224
rect 108004 64164 108008 64220
rect 108008 64164 108064 64220
rect 108064 64164 108068 64220
rect 108004 64160 108068 64164
rect 36075 64092 36139 64156
rect 43576 64092 43640 64156
rect 87310 64092 87374 64156
rect 41067 63956 41131 64020
rect 86142 63956 86206 64020
rect 38571 63820 38635 63884
rect 53547 63820 53611 63884
rect 95858 63880 95922 63884
rect 95858 63824 95882 63880
rect 95882 63824 95922 63880
rect 95858 63820 95922 63824
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 107028 63676 107092 63680
rect 107028 63620 107032 63676
rect 107032 63620 107088 63676
rect 107088 63620 107092 63676
rect 107028 63616 107092 63620
rect 107108 63676 107172 63680
rect 107108 63620 107112 63676
rect 107112 63620 107168 63676
rect 107168 63620 107172 63676
rect 107108 63616 107172 63620
rect 107188 63676 107252 63680
rect 107188 63620 107192 63676
rect 107192 63620 107248 63676
rect 107248 63620 107252 63676
rect 107188 63616 107252 63620
rect 107268 63676 107332 63680
rect 107268 63620 107272 63676
rect 107272 63620 107328 63676
rect 107328 63620 107332 63676
rect 107268 63616 107332 63620
rect 4876 63132 4940 63136
rect 4876 63076 4880 63132
rect 4880 63076 4936 63132
rect 4936 63076 4940 63132
rect 4876 63072 4940 63076
rect 4956 63132 5020 63136
rect 4956 63076 4960 63132
rect 4960 63076 5016 63132
rect 5016 63076 5020 63132
rect 4956 63072 5020 63076
rect 5036 63132 5100 63136
rect 5036 63076 5040 63132
rect 5040 63076 5096 63132
rect 5096 63076 5100 63132
rect 5036 63072 5100 63076
rect 5116 63132 5180 63136
rect 5116 63076 5120 63132
rect 5120 63076 5176 63132
rect 5176 63076 5180 63132
rect 5116 63072 5180 63076
rect 107764 63132 107828 63136
rect 107764 63076 107768 63132
rect 107768 63076 107824 63132
rect 107824 63076 107828 63132
rect 107764 63072 107828 63076
rect 107844 63132 107908 63136
rect 107844 63076 107848 63132
rect 107848 63076 107904 63132
rect 107904 63076 107908 63132
rect 107844 63072 107908 63076
rect 107924 63132 107988 63136
rect 107924 63076 107928 63132
rect 107928 63076 107984 63132
rect 107984 63076 107988 63132
rect 107924 63072 107988 63076
rect 108004 63132 108068 63136
rect 108004 63076 108008 63132
rect 108008 63076 108064 63132
rect 108064 63076 108068 63132
rect 108004 63072 108068 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 107028 62588 107092 62592
rect 107028 62532 107032 62588
rect 107032 62532 107088 62588
rect 107088 62532 107092 62588
rect 107028 62528 107092 62532
rect 107108 62588 107172 62592
rect 107108 62532 107112 62588
rect 107112 62532 107168 62588
rect 107168 62532 107172 62588
rect 107108 62528 107172 62532
rect 107188 62588 107252 62592
rect 107188 62532 107192 62588
rect 107192 62532 107248 62588
rect 107248 62532 107252 62588
rect 107188 62528 107252 62532
rect 107268 62588 107332 62592
rect 107268 62532 107272 62588
rect 107272 62532 107328 62588
rect 107328 62532 107332 62588
rect 107268 62528 107332 62532
rect 4876 62044 4940 62048
rect 4876 61988 4880 62044
rect 4880 61988 4936 62044
rect 4936 61988 4940 62044
rect 4876 61984 4940 61988
rect 4956 62044 5020 62048
rect 4956 61988 4960 62044
rect 4960 61988 5016 62044
rect 5016 61988 5020 62044
rect 4956 61984 5020 61988
rect 5036 62044 5100 62048
rect 5036 61988 5040 62044
rect 5040 61988 5096 62044
rect 5096 61988 5100 62044
rect 5036 61984 5100 61988
rect 5116 62044 5180 62048
rect 5116 61988 5120 62044
rect 5120 61988 5176 62044
rect 5176 61988 5180 62044
rect 5116 61984 5180 61988
rect 107764 62044 107828 62048
rect 107764 61988 107768 62044
rect 107768 61988 107824 62044
rect 107824 61988 107828 62044
rect 107764 61984 107828 61988
rect 107844 62044 107908 62048
rect 107844 61988 107848 62044
rect 107848 61988 107904 62044
rect 107904 61988 107908 62044
rect 107844 61984 107908 61988
rect 107924 62044 107988 62048
rect 107924 61988 107928 62044
rect 107928 61988 107984 62044
rect 107984 61988 107988 62044
rect 107924 61984 107988 61988
rect 108004 62044 108068 62048
rect 108004 61988 108008 62044
rect 108008 61988 108064 62044
rect 108064 61988 108068 62044
rect 108004 61984 108068 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 107028 61500 107092 61504
rect 107028 61444 107032 61500
rect 107032 61444 107088 61500
rect 107088 61444 107092 61500
rect 107028 61440 107092 61444
rect 107108 61500 107172 61504
rect 107108 61444 107112 61500
rect 107112 61444 107168 61500
rect 107168 61444 107172 61500
rect 107108 61440 107172 61444
rect 107188 61500 107252 61504
rect 107188 61444 107192 61500
rect 107192 61444 107248 61500
rect 107248 61444 107252 61500
rect 107188 61440 107252 61444
rect 107268 61500 107332 61504
rect 107268 61444 107272 61500
rect 107272 61444 107328 61500
rect 107328 61444 107332 61500
rect 107268 61440 107332 61444
rect 4876 60956 4940 60960
rect 4876 60900 4880 60956
rect 4880 60900 4936 60956
rect 4936 60900 4940 60956
rect 4876 60896 4940 60900
rect 4956 60956 5020 60960
rect 4956 60900 4960 60956
rect 4960 60900 5016 60956
rect 5016 60900 5020 60956
rect 4956 60896 5020 60900
rect 5036 60956 5100 60960
rect 5036 60900 5040 60956
rect 5040 60900 5096 60956
rect 5096 60900 5100 60956
rect 5036 60896 5100 60900
rect 5116 60956 5180 60960
rect 5116 60900 5120 60956
rect 5120 60900 5176 60956
rect 5176 60900 5180 60956
rect 5116 60896 5180 60900
rect 107764 60956 107828 60960
rect 107764 60900 107768 60956
rect 107768 60900 107824 60956
rect 107824 60900 107828 60956
rect 107764 60896 107828 60900
rect 107844 60956 107908 60960
rect 107844 60900 107848 60956
rect 107848 60900 107904 60956
rect 107904 60900 107908 60956
rect 107844 60896 107908 60900
rect 107924 60956 107988 60960
rect 107924 60900 107928 60956
rect 107928 60900 107984 60956
rect 107984 60900 107988 60956
rect 107924 60896 107988 60900
rect 108004 60956 108068 60960
rect 108004 60900 108008 60956
rect 108008 60900 108064 60956
rect 108064 60900 108068 60956
rect 108004 60896 108068 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 107028 60412 107092 60416
rect 107028 60356 107032 60412
rect 107032 60356 107088 60412
rect 107088 60356 107092 60412
rect 107028 60352 107092 60356
rect 107108 60412 107172 60416
rect 107108 60356 107112 60412
rect 107112 60356 107168 60412
rect 107168 60356 107172 60412
rect 107108 60352 107172 60356
rect 107188 60412 107252 60416
rect 107188 60356 107192 60412
rect 107192 60356 107248 60412
rect 107248 60356 107252 60412
rect 107188 60352 107252 60356
rect 107268 60412 107332 60416
rect 107268 60356 107272 60412
rect 107272 60356 107328 60412
rect 107328 60356 107332 60412
rect 107268 60352 107332 60356
rect 4876 59868 4940 59872
rect 4876 59812 4880 59868
rect 4880 59812 4936 59868
rect 4936 59812 4940 59868
rect 4876 59808 4940 59812
rect 4956 59868 5020 59872
rect 4956 59812 4960 59868
rect 4960 59812 5016 59868
rect 5016 59812 5020 59868
rect 4956 59808 5020 59812
rect 5036 59868 5100 59872
rect 5036 59812 5040 59868
rect 5040 59812 5096 59868
rect 5096 59812 5100 59868
rect 5036 59808 5100 59812
rect 5116 59868 5180 59872
rect 5116 59812 5120 59868
rect 5120 59812 5176 59868
rect 5176 59812 5180 59868
rect 5116 59808 5180 59812
rect 107764 59868 107828 59872
rect 107764 59812 107768 59868
rect 107768 59812 107824 59868
rect 107824 59812 107828 59868
rect 107764 59808 107828 59812
rect 107844 59868 107908 59872
rect 107844 59812 107848 59868
rect 107848 59812 107904 59868
rect 107904 59812 107908 59868
rect 107844 59808 107908 59812
rect 107924 59868 107988 59872
rect 107924 59812 107928 59868
rect 107928 59812 107984 59868
rect 107984 59812 107988 59868
rect 107924 59808 107988 59812
rect 108004 59868 108068 59872
rect 108004 59812 108008 59868
rect 108008 59812 108064 59868
rect 108064 59812 108068 59868
rect 108004 59808 108068 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 107028 59324 107092 59328
rect 107028 59268 107032 59324
rect 107032 59268 107088 59324
rect 107088 59268 107092 59324
rect 107028 59264 107092 59268
rect 107108 59324 107172 59328
rect 107108 59268 107112 59324
rect 107112 59268 107168 59324
rect 107168 59268 107172 59324
rect 107108 59264 107172 59268
rect 107188 59324 107252 59328
rect 107188 59268 107192 59324
rect 107192 59268 107248 59324
rect 107248 59268 107252 59324
rect 107188 59264 107252 59268
rect 107268 59324 107332 59328
rect 107268 59268 107272 59324
rect 107272 59268 107328 59324
rect 107328 59268 107332 59324
rect 107268 59264 107332 59268
rect 4876 58780 4940 58784
rect 4876 58724 4880 58780
rect 4880 58724 4936 58780
rect 4936 58724 4940 58780
rect 4876 58720 4940 58724
rect 4956 58780 5020 58784
rect 4956 58724 4960 58780
rect 4960 58724 5016 58780
rect 5016 58724 5020 58780
rect 4956 58720 5020 58724
rect 5036 58780 5100 58784
rect 5036 58724 5040 58780
rect 5040 58724 5096 58780
rect 5096 58724 5100 58780
rect 5036 58720 5100 58724
rect 5116 58780 5180 58784
rect 5116 58724 5120 58780
rect 5120 58724 5176 58780
rect 5176 58724 5180 58780
rect 5116 58720 5180 58724
rect 107764 58780 107828 58784
rect 107764 58724 107768 58780
rect 107768 58724 107824 58780
rect 107824 58724 107828 58780
rect 107764 58720 107828 58724
rect 107844 58780 107908 58784
rect 107844 58724 107848 58780
rect 107848 58724 107904 58780
rect 107904 58724 107908 58780
rect 107844 58720 107908 58724
rect 107924 58780 107988 58784
rect 107924 58724 107928 58780
rect 107928 58724 107984 58780
rect 107984 58724 107988 58780
rect 107924 58720 107988 58724
rect 108004 58780 108068 58784
rect 108004 58724 108008 58780
rect 108008 58724 108064 58780
rect 108064 58724 108068 58780
rect 108004 58720 108068 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 107028 58236 107092 58240
rect 107028 58180 107032 58236
rect 107032 58180 107088 58236
rect 107088 58180 107092 58236
rect 107028 58176 107092 58180
rect 107108 58236 107172 58240
rect 107108 58180 107112 58236
rect 107112 58180 107168 58236
rect 107168 58180 107172 58236
rect 107108 58176 107172 58180
rect 107188 58236 107252 58240
rect 107188 58180 107192 58236
rect 107192 58180 107248 58236
rect 107248 58180 107252 58236
rect 107188 58176 107252 58180
rect 107268 58236 107332 58240
rect 107268 58180 107272 58236
rect 107272 58180 107328 58236
rect 107328 58180 107332 58236
rect 107268 58176 107332 58180
rect 4876 57692 4940 57696
rect 4876 57636 4880 57692
rect 4880 57636 4936 57692
rect 4936 57636 4940 57692
rect 4876 57632 4940 57636
rect 4956 57692 5020 57696
rect 4956 57636 4960 57692
rect 4960 57636 5016 57692
rect 5016 57636 5020 57692
rect 4956 57632 5020 57636
rect 5036 57692 5100 57696
rect 5036 57636 5040 57692
rect 5040 57636 5096 57692
rect 5096 57636 5100 57692
rect 5036 57632 5100 57636
rect 5116 57692 5180 57696
rect 5116 57636 5120 57692
rect 5120 57636 5176 57692
rect 5176 57636 5180 57692
rect 5116 57632 5180 57636
rect 107764 57692 107828 57696
rect 107764 57636 107768 57692
rect 107768 57636 107824 57692
rect 107824 57636 107828 57692
rect 107764 57632 107828 57636
rect 107844 57692 107908 57696
rect 107844 57636 107848 57692
rect 107848 57636 107904 57692
rect 107904 57636 107908 57692
rect 107844 57632 107908 57636
rect 107924 57692 107988 57696
rect 107924 57636 107928 57692
rect 107928 57636 107984 57692
rect 107984 57636 107988 57692
rect 107924 57632 107988 57636
rect 108004 57692 108068 57696
rect 108004 57636 108008 57692
rect 108008 57636 108064 57692
rect 108064 57636 108068 57692
rect 108004 57632 108068 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 107028 57148 107092 57152
rect 107028 57092 107032 57148
rect 107032 57092 107088 57148
rect 107088 57092 107092 57148
rect 107028 57088 107092 57092
rect 107108 57148 107172 57152
rect 107108 57092 107112 57148
rect 107112 57092 107168 57148
rect 107168 57092 107172 57148
rect 107108 57088 107172 57092
rect 107188 57148 107252 57152
rect 107188 57092 107192 57148
rect 107192 57092 107248 57148
rect 107248 57092 107252 57148
rect 107188 57088 107252 57092
rect 107268 57148 107332 57152
rect 107268 57092 107272 57148
rect 107272 57092 107328 57148
rect 107328 57092 107332 57148
rect 107268 57088 107332 57092
rect 4876 56604 4940 56608
rect 4876 56548 4880 56604
rect 4880 56548 4936 56604
rect 4936 56548 4940 56604
rect 4876 56544 4940 56548
rect 4956 56604 5020 56608
rect 4956 56548 4960 56604
rect 4960 56548 5016 56604
rect 5016 56548 5020 56604
rect 4956 56544 5020 56548
rect 5036 56604 5100 56608
rect 5036 56548 5040 56604
rect 5040 56548 5096 56604
rect 5096 56548 5100 56604
rect 5036 56544 5100 56548
rect 5116 56604 5180 56608
rect 5116 56548 5120 56604
rect 5120 56548 5176 56604
rect 5176 56548 5180 56604
rect 5116 56544 5180 56548
rect 107764 56604 107828 56608
rect 107764 56548 107768 56604
rect 107768 56548 107824 56604
rect 107824 56548 107828 56604
rect 107764 56544 107828 56548
rect 107844 56604 107908 56608
rect 107844 56548 107848 56604
rect 107848 56548 107904 56604
rect 107904 56548 107908 56604
rect 107844 56544 107908 56548
rect 107924 56604 107988 56608
rect 107924 56548 107928 56604
rect 107928 56548 107984 56604
rect 107984 56548 107988 56604
rect 107924 56544 107988 56548
rect 108004 56604 108068 56608
rect 108004 56548 108008 56604
rect 108008 56548 108064 56604
rect 108064 56548 108068 56604
rect 108004 56544 108068 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 107028 56060 107092 56064
rect 107028 56004 107032 56060
rect 107032 56004 107088 56060
rect 107088 56004 107092 56060
rect 107028 56000 107092 56004
rect 107108 56060 107172 56064
rect 107108 56004 107112 56060
rect 107112 56004 107168 56060
rect 107168 56004 107172 56060
rect 107108 56000 107172 56004
rect 107188 56060 107252 56064
rect 107188 56004 107192 56060
rect 107192 56004 107248 56060
rect 107248 56004 107252 56060
rect 107188 56000 107252 56004
rect 107268 56060 107332 56064
rect 107268 56004 107272 56060
rect 107272 56004 107328 56060
rect 107328 56004 107332 56060
rect 107268 56000 107332 56004
rect 4876 55516 4940 55520
rect 4876 55460 4880 55516
rect 4880 55460 4936 55516
rect 4936 55460 4940 55516
rect 4876 55456 4940 55460
rect 4956 55516 5020 55520
rect 4956 55460 4960 55516
rect 4960 55460 5016 55516
rect 5016 55460 5020 55516
rect 4956 55456 5020 55460
rect 5036 55516 5100 55520
rect 5036 55460 5040 55516
rect 5040 55460 5096 55516
rect 5096 55460 5100 55516
rect 5036 55456 5100 55460
rect 5116 55516 5180 55520
rect 5116 55460 5120 55516
rect 5120 55460 5176 55516
rect 5176 55460 5180 55516
rect 5116 55456 5180 55460
rect 107764 55516 107828 55520
rect 107764 55460 107768 55516
rect 107768 55460 107824 55516
rect 107824 55460 107828 55516
rect 107764 55456 107828 55460
rect 107844 55516 107908 55520
rect 107844 55460 107848 55516
rect 107848 55460 107904 55516
rect 107904 55460 107908 55516
rect 107844 55456 107908 55460
rect 107924 55516 107988 55520
rect 107924 55460 107928 55516
rect 107928 55460 107984 55516
rect 107984 55460 107988 55516
rect 107924 55456 107988 55460
rect 108004 55516 108068 55520
rect 108004 55460 108008 55516
rect 108008 55460 108064 55516
rect 108064 55460 108068 55516
rect 108004 55456 108068 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 107028 54972 107092 54976
rect 107028 54916 107032 54972
rect 107032 54916 107088 54972
rect 107088 54916 107092 54972
rect 107028 54912 107092 54916
rect 107108 54972 107172 54976
rect 107108 54916 107112 54972
rect 107112 54916 107168 54972
rect 107168 54916 107172 54972
rect 107108 54912 107172 54916
rect 107188 54972 107252 54976
rect 107188 54916 107192 54972
rect 107192 54916 107248 54972
rect 107248 54916 107252 54972
rect 107188 54912 107252 54916
rect 107268 54972 107332 54976
rect 107268 54916 107272 54972
rect 107272 54916 107328 54972
rect 107328 54916 107332 54972
rect 107268 54912 107332 54916
rect 4876 54428 4940 54432
rect 4876 54372 4880 54428
rect 4880 54372 4936 54428
rect 4936 54372 4940 54428
rect 4876 54368 4940 54372
rect 4956 54428 5020 54432
rect 4956 54372 4960 54428
rect 4960 54372 5016 54428
rect 5016 54372 5020 54428
rect 4956 54368 5020 54372
rect 5036 54428 5100 54432
rect 5036 54372 5040 54428
rect 5040 54372 5096 54428
rect 5096 54372 5100 54428
rect 5036 54368 5100 54372
rect 5116 54428 5180 54432
rect 5116 54372 5120 54428
rect 5120 54372 5176 54428
rect 5176 54372 5180 54428
rect 5116 54368 5180 54372
rect 107764 54428 107828 54432
rect 107764 54372 107768 54428
rect 107768 54372 107824 54428
rect 107824 54372 107828 54428
rect 107764 54368 107828 54372
rect 107844 54428 107908 54432
rect 107844 54372 107848 54428
rect 107848 54372 107904 54428
rect 107904 54372 107908 54428
rect 107844 54368 107908 54372
rect 107924 54428 107988 54432
rect 107924 54372 107928 54428
rect 107928 54372 107984 54428
rect 107984 54372 107988 54428
rect 107924 54368 107988 54372
rect 108004 54428 108068 54432
rect 108004 54372 108008 54428
rect 108008 54372 108064 54428
rect 108064 54372 108068 54428
rect 108004 54368 108068 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 107028 53884 107092 53888
rect 107028 53828 107032 53884
rect 107032 53828 107088 53884
rect 107088 53828 107092 53884
rect 107028 53824 107092 53828
rect 107108 53884 107172 53888
rect 107108 53828 107112 53884
rect 107112 53828 107168 53884
rect 107168 53828 107172 53884
rect 107108 53824 107172 53828
rect 107188 53884 107252 53888
rect 107188 53828 107192 53884
rect 107192 53828 107248 53884
rect 107248 53828 107252 53884
rect 107188 53824 107252 53828
rect 107268 53884 107332 53888
rect 107268 53828 107272 53884
rect 107272 53828 107328 53884
rect 107328 53828 107332 53884
rect 107268 53824 107332 53828
rect 4876 53340 4940 53344
rect 4876 53284 4880 53340
rect 4880 53284 4936 53340
rect 4936 53284 4940 53340
rect 4876 53280 4940 53284
rect 4956 53340 5020 53344
rect 4956 53284 4960 53340
rect 4960 53284 5016 53340
rect 5016 53284 5020 53340
rect 4956 53280 5020 53284
rect 5036 53340 5100 53344
rect 5036 53284 5040 53340
rect 5040 53284 5096 53340
rect 5096 53284 5100 53340
rect 5036 53280 5100 53284
rect 5116 53340 5180 53344
rect 5116 53284 5120 53340
rect 5120 53284 5176 53340
rect 5176 53284 5180 53340
rect 5116 53280 5180 53284
rect 107764 53340 107828 53344
rect 107764 53284 107768 53340
rect 107768 53284 107824 53340
rect 107824 53284 107828 53340
rect 107764 53280 107828 53284
rect 107844 53340 107908 53344
rect 107844 53284 107848 53340
rect 107848 53284 107904 53340
rect 107904 53284 107908 53340
rect 107844 53280 107908 53284
rect 107924 53340 107988 53344
rect 107924 53284 107928 53340
rect 107928 53284 107984 53340
rect 107984 53284 107988 53340
rect 107924 53280 107988 53284
rect 108004 53340 108068 53344
rect 108004 53284 108008 53340
rect 108008 53284 108064 53340
rect 108064 53284 108068 53340
rect 108004 53280 108068 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 107028 52796 107092 52800
rect 107028 52740 107032 52796
rect 107032 52740 107088 52796
rect 107088 52740 107092 52796
rect 107028 52736 107092 52740
rect 107108 52796 107172 52800
rect 107108 52740 107112 52796
rect 107112 52740 107168 52796
rect 107168 52740 107172 52796
rect 107108 52736 107172 52740
rect 107188 52796 107252 52800
rect 107188 52740 107192 52796
rect 107192 52740 107248 52796
rect 107248 52740 107252 52796
rect 107188 52736 107252 52740
rect 107268 52796 107332 52800
rect 107268 52740 107272 52796
rect 107272 52740 107328 52796
rect 107328 52740 107332 52796
rect 107268 52736 107332 52740
rect 4876 52252 4940 52256
rect 4876 52196 4880 52252
rect 4880 52196 4936 52252
rect 4936 52196 4940 52252
rect 4876 52192 4940 52196
rect 4956 52252 5020 52256
rect 4956 52196 4960 52252
rect 4960 52196 5016 52252
rect 5016 52196 5020 52252
rect 4956 52192 5020 52196
rect 5036 52252 5100 52256
rect 5036 52196 5040 52252
rect 5040 52196 5096 52252
rect 5096 52196 5100 52252
rect 5036 52192 5100 52196
rect 5116 52252 5180 52256
rect 5116 52196 5120 52252
rect 5120 52196 5176 52252
rect 5176 52196 5180 52252
rect 5116 52192 5180 52196
rect 107764 52252 107828 52256
rect 107764 52196 107768 52252
rect 107768 52196 107824 52252
rect 107824 52196 107828 52252
rect 107764 52192 107828 52196
rect 107844 52252 107908 52256
rect 107844 52196 107848 52252
rect 107848 52196 107904 52252
rect 107904 52196 107908 52252
rect 107844 52192 107908 52196
rect 107924 52252 107988 52256
rect 107924 52196 107928 52252
rect 107928 52196 107984 52252
rect 107984 52196 107988 52252
rect 107924 52192 107988 52196
rect 108004 52252 108068 52256
rect 108004 52196 108008 52252
rect 108008 52196 108064 52252
rect 108064 52196 108068 52252
rect 108004 52192 108068 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 107028 51708 107092 51712
rect 107028 51652 107032 51708
rect 107032 51652 107088 51708
rect 107088 51652 107092 51708
rect 107028 51648 107092 51652
rect 107108 51708 107172 51712
rect 107108 51652 107112 51708
rect 107112 51652 107168 51708
rect 107168 51652 107172 51708
rect 107108 51648 107172 51652
rect 107188 51708 107252 51712
rect 107188 51652 107192 51708
rect 107192 51652 107248 51708
rect 107248 51652 107252 51708
rect 107188 51648 107252 51652
rect 107268 51708 107332 51712
rect 107268 51652 107272 51708
rect 107272 51652 107328 51708
rect 107328 51652 107332 51708
rect 107268 51648 107332 51652
rect 4876 51164 4940 51168
rect 4876 51108 4880 51164
rect 4880 51108 4936 51164
rect 4936 51108 4940 51164
rect 4876 51104 4940 51108
rect 4956 51164 5020 51168
rect 4956 51108 4960 51164
rect 4960 51108 5016 51164
rect 5016 51108 5020 51164
rect 4956 51104 5020 51108
rect 5036 51164 5100 51168
rect 5036 51108 5040 51164
rect 5040 51108 5096 51164
rect 5096 51108 5100 51164
rect 5036 51104 5100 51108
rect 5116 51164 5180 51168
rect 5116 51108 5120 51164
rect 5120 51108 5176 51164
rect 5176 51108 5180 51164
rect 5116 51104 5180 51108
rect 107764 51164 107828 51168
rect 107764 51108 107768 51164
rect 107768 51108 107824 51164
rect 107824 51108 107828 51164
rect 107764 51104 107828 51108
rect 107844 51164 107908 51168
rect 107844 51108 107848 51164
rect 107848 51108 107904 51164
rect 107904 51108 107908 51164
rect 107844 51104 107908 51108
rect 107924 51164 107988 51168
rect 107924 51108 107928 51164
rect 107928 51108 107984 51164
rect 107984 51108 107988 51164
rect 107924 51104 107988 51108
rect 108004 51164 108068 51168
rect 108004 51108 108008 51164
rect 108008 51108 108064 51164
rect 108064 51108 108068 51164
rect 108004 51104 108068 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 107028 50620 107092 50624
rect 107028 50564 107032 50620
rect 107032 50564 107088 50620
rect 107088 50564 107092 50620
rect 107028 50560 107092 50564
rect 107108 50620 107172 50624
rect 107108 50564 107112 50620
rect 107112 50564 107168 50620
rect 107168 50564 107172 50620
rect 107108 50560 107172 50564
rect 107188 50620 107252 50624
rect 107188 50564 107192 50620
rect 107192 50564 107248 50620
rect 107248 50564 107252 50620
rect 107188 50560 107252 50564
rect 107268 50620 107332 50624
rect 107268 50564 107272 50620
rect 107272 50564 107328 50620
rect 107328 50564 107332 50620
rect 107268 50560 107332 50564
rect 4876 50076 4940 50080
rect 4876 50020 4880 50076
rect 4880 50020 4936 50076
rect 4936 50020 4940 50076
rect 4876 50016 4940 50020
rect 4956 50076 5020 50080
rect 4956 50020 4960 50076
rect 4960 50020 5016 50076
rect 5016 50020 5020 50076
rect 4956 50016 5020 50020
rect 5036 50076 5100 50080
rect 5036 50020 5040 50076
rect 5040 50020 5096 50076
rect 5096 50020 5100 50076
rect 5036 50016 5100 50020
rect 5116 50076 5180 50080
rect 5116 50020 5120 50076
rect 5120 50020 5176 50076
rect 5176 50020 5180 50076
rect 5116 50016 5180 50020
rect 107764 50076 107828 50080
rect 107764 50020 107768 50076
rect 107768 50020 107824 50076
rect 107824 50020 107828 50076
rect 107764 50016 107828 50020
rect 107844 50076 107908 50080
rect 107844 50020 107848 50076
rect 107848 50020 107904 50076
rect 107904 50020 107908 50076
rect 107844 50016 107908 50020
rect 107924 50076 107988 50080
rect 107924 50020 107928 50076
rect 107928 50020 107984 50076
rect 107984 50020 107988 50076
rect 107924 50016 107988 50020
rect 108004 50076 108068 50080
rect 108004 50020 108008 50076
rect 108008 50020 108064 50076
rect 108064 50020 108068 50076
rect 108004 50016 108068 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 107028 49532 107092 49536
rect 107028 49476 107032 49532
rect 107032 49476 107088 49532
rect 107088 49476 107092 49532
rect 107028 49472 107092 49476
rect 107108 49532 107172 49536
rect 107108 49476 107112 49532
rect 107112 49476 107168 49532
rect 107168 49476 107172 49532
rect 107108 49472 107172 49476
rect 107188 49532 107252 49536
rect 107188 49476 107192 49532
rect 107192 49476 107248 49532
rect 107248 49476 107252 49532
rect 107188 49472 107252 49476
rect 107268 49532 107332 49536
rect 107268 49476 107272 49532
rect 107272 49476 107328 49532
rect 107328 49476 107332 49532
rect 107268 49472 107332 49476
rect 4876 48988 4940 48992
rect 4876 48932 4880 48988
rect 4880 48932 4936 48988
rect 4936 48932 4940 48988
rect 4876 48928 4940 48932
rect 4956 48988 5020 48992
rect 4956 48932 4960 48988
rect 4960 48932 5016 48988
rect 5016 48932 5020 48988
rect 4956 48928 5020 48932
rect 5036 48988 5100 48992
rect 5036 48932 5040 48988
rect 5040 48932 5096 48988
rect 5096 48932 5100 48988
rect 5036 48928 5100 48932
rect 5116 48988 5180 48992
rect 5116 48932 5120 48988
rect 5120 48932 5176 48988
rect 5176 48932 5180 48988
rect 5116 48928 5180 48932
rect 107764 48988 107828 48992
rect 107764 48932 107768 48988
rect 107768 48932 107824 48988
rect 107824 48932 107828 48988
rect 107764 48928 107828 48932
rect 107844 48988 107908 48992
rect 107844 48932 107848 48988
rect 107848 48932 107904 48988
rect 107904 48932 107908 48988
rect 107844 48928 107908 48932
rect 107924 48988 107988 48992
rect 107924 48932 107928 48988
rect 107928 48932 107984 48988
rect 107984 48932 107988 48988
rect 107924 48928 107988 48932
rect 108004 48988 108068 48992
rect 108004 48932 108008 48988
rect 108008 48932 108064 48988
rect 108064 48932 108068 48988
rect 108004 48928 108068 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 107028 48444 107092 48448
rect 107028 48388 107032 48444
rect 107032 48388 107088 48444
rect 107088 48388 107092 48444
rect 107028 48384 107092 48388
rect 107108 48444 107172 48448
rect 107108 48388 107112 48444
rect 107112 48388 107168 48444
rect 107168 48388 107172 48444
rect 107108 48384 107172 48388
rect 107188 48444 107252 48448
rect 107188 48388 107192 48444
rect 107192 48388 107248 48444
rect 107248 48388 107252 48444
rect 107188 48384 107252 48388
rect 107268 48444 107332 48448
rect 107268 48388 107272 48444
rect 107272 48388 107328 48444
rect 107328 48388 107332 48444
rect 107268 48384 107332 48388
rect 4876 47900 4940 47904
rect 4876 47844 4880 47900
rect 4880 47844 4936 47900
rect 4936 47844 4940 47900
rect 4876 47840 4940 47844
rect 4956 47900 5020 47904
rect 4956 47844 4960 47900
rect 4960 47844 5016 47900
rect 5016 47844 5020 47900
rect 4956 47840 5020 47844
rect 5036 47900 5100 47904
rect 5036 47844 5040 47900
rect 5040 47844 5096 47900
rect 5096 47844 5100 47900
rect 5036 47840 5100 47844
rect 5116 47900 5180 47904
rect 5116 47844 5120 47900
rect 5120 47844 5176 47900
rect 5176 47844 5180 47900
rect 5116 47840 5180 47844
rect 107764 47900 107828 47904
rect 107764 47844 107768 47900
rect 107768 47844 107824 47900
rect 107824 47844 107828 47900
rect 107764 47840 107828 47844
rect 107844 47900 107908 47904
rect 107844 47844 107848 47900
rect 107848 47844 107904 47900
rect 107904 47844 107908 47900
rect 107844 47840 107908 47844
rect 107924 47900 107988 47904
rect 107924 47844 107928 47900
rect 107928 47844 107984 47900
rect 107984 47844 107988 47900
rect 107924 47840 107988 47844
rect 108004 47900 108068 47904
rect 108004 47844 108008 47900
rect 108008 47844 108064 47900
rect 108064 47844 108068 47900
rect 108004 47840 108068 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 107028 47356 107092 47360
rect 107028 47300 107032 47356
rect 107032 47300 107088 47356
rect 107088 47300 107092 47356
rect 107028 47296 107092 47300
rect 107108 47356 107172 47360
rect 107108 47300 107112 47356
rect 107112 47300 107168 47356
rect 107168 47300 107172 47356
rect 107108 47296 107172 47300
rect 107188 47356 107252 47360
rect 107188 47300 107192 47356
rect 107192 47300 107248 47356
rect 107248 47300 107252 47356
rect 107188 47296 107252 47300
rect 107268 47356 107332 47360
rect 107268 47300 107272 47356
rect 107272 47300 107328 47356
rect 107328 47300 107332 47356
rect 107268 47296 107332 47300
rect 4876 46812 4940 46816
rect 4876 46756 4880 46812
rect 4880 46756 4936 46812
rect 4936 46756 4940 46812
rect 4876 46752 4940 46756
rect 4956 46812 5020 46816
rect 4956 46756 4960 46812
rect 4960 46756 5016 46812
rect 5016 46756 5020 46812
rect 4956 46752 5020 46756
rect 5036 46812 5100 46816
rect 5036 46756 5040 46812
rect 5040 46756 5096 46812
rect 5096 46756 5100 46812
rect 5036 46752 5100 46756
rect 5116 46812 5180 46816
rect 5116 46756 5120 46812
rect 5120 46756 5176 46812
rect 5176 46756 5180 46812
rect 5116 46752 5180 46756
rect 107764 46812 107828 46816
rect 107764 46756 107768 46812
rect 107768 46756 107824 46812
rect 107824 46756 107828 46812
rect 107764 46752 107828 46756
rect 107844 46812 107908 46816
rect 107844 46756 107848 46812
rect 107848 46756 107904 46812
rect 107904 46756 107908 46812
rect 107844 46752 107908 46756
rect 107924 46812 107988 46816
rect 107924 46756 107928 46812
rect 107928 46756 107984 46812
rect 107984 46756 107988 46812
rect 107924 46752 107988 46756
rect 108004 46812 108068 46816
rect 108004 46756 108008 46812
rect 108008 46756 108064 46812
rect 108064 46756 108068 46812
rect 108004 46752 108068 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 107028 46268 107092 46272
rect 107028 46212 107032 46268
rect 107032 46212 107088 46268
rect 107088 46212 107092 46268
rect 107028 46208 107092 46212
rect 107108 46268 107172 46272
rect 107108 46212 107112 46268
rect 107112 46212 107168 46268
rect 107168 46212 107172 46268
rect 107108 46208 107172 46212
rect 107188 46268 107252 46272
rect 107188 46212 107192 46268
rect 107192 46212 107248 46268
rect 107248 46212 107252 46268
rect 107188 46208 107252 46212
rect 107268 46268 107332 46272
rect 107268 46212 107272 46268
rect 107272 46212 107328 46268
rect 107328 46212 107332 46268
rect 107268 46208 107332 46212
rect 4876 45724 4940 45728
rect 4876 45668 4880 45724
rect 4880 45668 4936 45724
rect 4936 45668 4940 45724
rect 4876 45664 4940 45668
rect 4956 45724 5020 45728
rect 4956 45668 4960 45724
rect 4960 45668 5016 45724
rect 5016 45668 5020 45724
rect 4956 45664 5020 45668
rect 5036 45724 5100 45728
rect 5036 45668 5040 45724
rect 5040 45668 5096 45724
rect 5096 45668 5100 45724
rect 5036 45664 5100 45668
rect 5116 45724 5180 45728
rect 5116 45668 5120 45724
rect 5120 45668 5176 45724
rect 5176 45668 5180 45724
rect 5116 45664 5180 45668
rect 107764 45724 107828 45728
rect 107764 45668 107768 45724
rect 107768 45668 107824 45724
rect 107824 45668 107828 45724
rect 107764 45664 107828 45668
rect 107844 45724 107908 45728
rect 107844 45668 107848 45724
rect 107848 45668 107904 45724
rect 107904 45668 107908 45724
rect 107844 45664 107908 45668
rect 107924 45724 107988 45728
rect 107924 45668 107928 45724
rect 107928 45668 107984 45724
rect 107984 45668 107988 45724
rect 107924 45664 107988 45668
rect 108004 45724 108068 45728
rect 108004 45668 108008 45724
rect 108008 45668 108064 45724
rect 108064 45668 108068 45724
rect 108004 45664 108068 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 107028 45180 107092 45184
rect 107028 45124 107032 45180
rect 107032 45124 107088 45180
rect 107088 45124 107092 45180
rect 107028 45120 107092 45124
rect 107108 45180 107172 45184
rect 107108 45124 107112 45180
rect 107112 45124 107168 45180
rect 107168 45124 107172 45180
rect 107108 45120 107172 45124
rect 107188 45180 107252 45184
rect 107188 45124 107192 45180
rect 107192 45124 107248 45180
rect 107248 45124 107252 45180
rect 107188 45120 107252 45124
rect 107268 45180 107332 45184
rect 107268 45124 107272 45180
rect 107272 45124 107328 45180
rect 107328 45124 107332 45180
rect 107268 45120 107332 45124
rect 4876 44636 4940 44640
rect 4876 44580 4880 44636
rect 4880 44580 4936 44636
rect 4936 44580 4940 44636
rect 4876 44576 4940 44580
rect 4956 44636 5020 44640
rect 4956 44580 4960 44636
rect 4960 44580 5016 44636
rect 5016 44580 5020 44636
rect 4956 44576 5020 44580
rect 5036 44636 5100 44640
rect 5036 44580 5040 44636
rect 5040 44580 5096 44636
rect 5096 44580 5100 44636
rect 5036 44576 5100 44580
rect 5116 44636 5180 44640
rect 5116 44580 5120 44636
rect 5120 44580 5176 44636
rect 5176 44580 5180 44636
rect 5116 44576 5180 44580
rect 107764 44636 107828 44640
rect 107764 44580 107768 44636
rect 107768 44580 107824 44636
rect 107824 44580 107828 44636
rect 107764 44576 107828 44580
rect 107844 44636 107908 44640
rect 107844 44580 107848 44636
rect 107848 44580 107904 44636
rect 107904 44580 107908 44636
rect 107844 44576 107908 44580
rect 107924 44636 107988 44640
rect 107924 44580 107928 44636
rect 107928 44580 107984 44636
rect 107984 44580 107988 44636
rect 107924 44576 107988 44580
rect 108004 44636 108068 44640
rect 108004 44580 108008 44636
rect 108008 44580 108064 44636
rect 108064 44580 108068 44636
rect 108004 44576 108068 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 107028 44092 107092 44096
rect 107028 44036 107032 44092
rect 107032 44036 107088 44092
rect 107088 44036 107092 44092
rect 107028 44032 107092 44036
rect 107108 44092 107172 44096
rect 107108 44036 107112 44092
rect 107112 44036 107168 44092
rect 107168 44036 107172 44092
rect 107108 44032 107172 44036
rect 107188 44092 107252 44096
rect 107188 44036 107192 44092
rect 107192 44036 107248 44092
rect 107248 44036 107252 44092
rect 107188 44032 107252 44036
rect 107268 44092 107332 44096
rect 107268 44036 107272 44092
rect 107272 44036 107328 44092
rect 107328 44036 107332 44092
rect 107268 44032 107332 44036
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 107764 43548 107828 43552
rect 107764 43492 107768 43548
rect 107768 43492 107824 43548
rect 107824 43492 107828 43548
rect 107764 43488 107828 43492
rect 107844 43548 107908 43552
rect 107844 43492 107848 43548
rect 107848 43492 107904 43548
rect 107904 43492 107908 43548
rect 107844 43488 107908 43492
rect 107924 43548 107988 43552
rect 107924 43492 107928 43548
rect 107928 43492 107984 43548
rect 107984 43492 107988 43548
rect 107924 43488 107988 43492
rect 108004 43548 108068 43552
rect 108004 43492 108008 43548
rect 108008 43492 108064 43548
rect 108064 43492 108068 43548
rect 108004 43488 108068 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 107028 43004 107092 43008
rect 107028 42948 107032 43004
rect 107032 42948 107088 43004
rect 107088 42948 107092 43004
rect 107028 42944 107092 42948
rect 107108 43004 107172 43008
rect 107108 42948 107112 43004
rect 107112 42948 107168 43004
rect 107168 42948 107172 43004
rect 107108 42944 107172 42948
rect 107188 43004 107252 43008
rect 107188 42948 107192 43004
rect 107192 42948 107248 43004
rect 107248 42948 107252 43004
rect 107188 42944 107252 42948
rect 107268 43004 107332 43008
rect 107268 42948 107272 43004
rect 107272 42948 107328 43004
rect 107328 42948 107332 43004
rect 107268 42944 107332 42948
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 107764 42460 107828 42464
rect 107764 42404 107768 42460
rect 107768 42404 107824 42460
rect 107824 42404 107828 42460
rect 107764 42400 107828 42404
rect 107844 42460 107908 42464
rect 107844 42404 107848 42460
rect 107848 42404 107904 42460
rect 107904 42404 107908 42460
rect 107844 42400 107908 42404
rect 107924 42460 107988 42464
rect 107924 42404 107928 42460
rect 107928 42404 107984 42460
rect 107984 42404 107988 42460
rect 107924 42400 107988 42404
rect 108004 42460 108068 42464
rect 108004 42404 108008 42460
rect 108008 42404 108064 42460
rect 108064 42404 108068 42460
rect 108004 42400 108068 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 107028 41916 107092 41920
rect 107028 41860 107032 41916
rect 107032 41860 107088 41916
rect 107088 41860 107092 41916
rect 107028 41856 107092 41860
rect 107108 41916 107172 41920
rect 107108 41860 107112 41916
rect 107112 41860 107168 41916
rect 107168 41860 107172 41916
rect 107108 41856 107172 41860
rect 107188 41916 107252 41920
rect 107188 41860 107192 41916
rect 107192 41860 107248 41916
rect 107248 41860 107252 41916
rect 107188 41856 107252 41860
rect 107268 41916 107332 41920
rect 107268 41860 107272 41916
rect 107272 41860 107328 41916
rect 107328 41860 107332 41916
rect 107268 41856 107332 41860
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 107764 41372 107828 41376
rect 107764 41316 107768 41372
rect 107768 41316 107824 41372
rect 107824 41316 107828 41372
rect 107764 41312 107828 41316
rect 107844 41372 107908 41376
rect 107844 41316 107848 41372
rect 107848 41316 107904 41372
rect 107904 41316 107908 41372
rect 107844 41312 107908 41316
rect 107924 41372 107988 41376
rect 107924 41316 107928 41372
rect 107928 41316 107984 41372
rect 107984 41316 107988 41372
rect 107924 41312 107988 41316
rect 108004 41372 108068 41376
rect 108004 41316 108008 41372
rect 108008 41316 108064 41372
rect 108064 41316 108068 41372
rect 108004 41312 108068 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 107028 40828 107092 40832
rect 107028 40772 107032 40828
rect 107032 40772 107088 40828
rect 107088 40772 107092 40828
rect 107028 40768 107092 40772
rect 107108 40828 107172 40832
rect 107108 40772 107112 40828
rect 107112 40772 107168 40828
rect 107168 40772 107172 40828
rect 107108 40768 107172 40772
rect 107188 40828 107252 40832
rect 107188 40772 107192 40828
rect 107192 40772 107248 40828
rect 107248 40772 107252 40828
rect 107188 40768 107252 40772
rect 107268 40828 107332 40832
rect 107268 40772 107272 40828
rect 107272 40772 107328 40828
rect 107328 40772 107332 40828
rect 107268 40768 107332 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 107764 40284 107828 40288
rect 107764 40228 107768 40284
rect 107768 40228 107824 40284
rect 107824 40228 107828 40284
rect 107764 40224 107828 40228
rect 107844 40284 107908 40288
rect 107844 40228 107848 40284
rect 107848 40228 107904 40284
rect 107904 40228 107908 40284
rect 107844 40224 107908 40228
rect 107924 40284 107988 40288
rect 107924 40228 107928 40284
rect 107928 40228 107984 40284
rect 107984 40228 107988 40284
rect 107924 40224 107988 40228
rect 108004 40284 108068 40288
rect 108004 40228 108008 40284
rect 108008 40228 108064 40284
rect 108064 40228 108068 40284
rect 108004 40224 108068 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 107028 39740 107092 39744
rect 107028 39684 107032 39740
rect 107032 39684 107088 39740
rect 107088 39684 107092 39740
rect 107028 39680 107092 39684
rect 107108 39740 107172 39744
rect 107108 39684 107112 39740
rect 107112 39684 107168 39740
rect 107168 39684 107172 39740
rect 107108 39680 107172 39684
rect 107188 39740 107252 39744
rect 107188 39684 107192 39740
rect 107192 39684 107248 39740
rect 107248 39684 107252 39740
rect 107188 39680 107252 39684
rect 107268 39740 107332 39744
rect 107268 39684 107272 39740
rect 107272 39684 107328 39740
rect 107328 39684 107332 39740
rect 107268 39680 107332 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 107764 39196 107828 39200
rect 107764 39140 107768 39196
rect 107768 39140 107824 39196
rect 107824 39140 107828 39196
rect 107764 39136 107828 39140
rect 107844 39196 107908 39200
rect 107844 39140 107848 39196
rect 107848 39140 107904 39196
rect 107904 39140 107908 39196
rect 107844 39136 107908 39140
rect 107924 39196 107988 39200
rect 107924 39140 107928 39196
rect 107928 39140 107984 39196
rect 107984 39140 107988 39196
rect 107924 39136 107988 39140
rect 108004 39196 108068 39200
rect 108004 39140 108008 39196
rect 108008 39140 108064 39196
rect 108064 39140 108068 39196
rect 108004 39136 108068 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 107028 38652 107092 38656
rect 107028 38596 107032 38652
rect 107032 38596 107088 38652
rect 107088 38596 107092 38652
rect 107028 38592 107092 38596
rect 107108 38652 107172 38656
rect 107108 38596 107112 38652
rect 107112 38596 107168 38652
rect 107168 38596 107172 38652
rect 107108 38592 107172 38596
rect 107188 38652 107252 38656
rect 107188 38596 107192 38652
rect 107192 38596 107248 38652
rect 107248 38596 107252 38652
rect 107188 38592 107252 38596
rect 107268 38652 107332 38656
rect 107268 38596 107272 38652
rect 107272 38596 107328 38652
rect 107328 38596 107332 38652
rect 107268 38592 107332 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 107764 38108 107828 38112
rect 107764 38052 107768 38108
rect 107768 38052 107824 38108
rect 107824 38052 107828 38108
rect 107764 38048 107828 38052
rect 107844 38108 107908 38112
rect 107844 38052 107848 38108
rect 107848 38052 107904 38108
rect 107904 38052 107908 38108
rect 107844 38048 107908 38052
rect 107924 38108 107988 38112
rect 107924 38052 107928 38108
rect 107928 38052 107984 38108
rect 107984 38052 107988 38108
rect 107924 38048 107988 38052
rect 108004 38108 108068 38112
rect 108004 38052 108008 38108
rect 108008 38052 108064 38108
rect 108064 38052 108068 38108
rect 108004 38048 108068 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 107028 37564 107092 37568
rect 107028 37508 107032 37564
rect 107032 37508 107088 37564
rect 107088 37508 107092 37564
rect 107028 37504 107092 37508
rect 107108 37564 107172 37568
rect 107108 37508 107112 37564
rect 107112 37508 107168 37564
rect 107168 37508 107172 37564
rect 107108 37504 107172 37508
rect 107188 37564 107252 37568
rect 107188 37508 107192 37564
rect 107192 37508 107248 37564
rect 107248 37508 107252 37564
rect 107188 37504 107252 37508
rect 107268 37564 107332 37568
rect 107268 37508 107272 37564
rect 107272 37508 107328 37564
rect 107328 37508 107332 37564
rect 107268 37504 107332 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 107764 37020 107828 37024
rect 107764 36964 107768 37020
rect 107768 36964 107824 37020
rect 107824 36964 107828 37020
rect 107764 36960 107828 36964
rect 107844 37020 107908 37024
rect 107844 36964 107848 37020
rect 107848 36964 107904 37020
rect 107904 36964 107908 37020
rect 107844 36960 107908 36964
rect 107924 37020 107988 37024
rect 107924 36964 107928 37020
rect 107928 36964 107984 37020
rect 107984 36964 107988 37020
rect 107924 36960 107988 36964
rect 108004 37020 108068 37024
rect 108004 36964 108008 37020
rect 108008 36964 108064 37020
rect 108064 36964 108068 37020
rect 108004 36960 108068 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 107028 36476 107092 36480
rect 107028 36420 107032 36476
rect 107032 36420 107088 36476
rect 107088 36420 107092 36476
rect 107028 36416 107092 36420
rect 107108 36476 107172 36480
rect 107108 36420 107112 36476
rect 107112 36420 107168 36476
rect 107168 36420 107172 36476
rect 107108 36416 107172 36420
rect 107188 36476 107252 36480
rect 107188 36420 107192 36476
rect 107192 36420 107248 36476
rect 107248 36420 107252 36476
rect 107188 36416 107252 36420
rect 107268 36476 107332 36480
rect 107268 36420 107272 36476
rect 107272 36420 107328 36476
rect 107328 36420 107332 36476
rect 107268 36416 107332 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 107764 35932 107828 35936
rect 107764 35876 107768 35932
rect 107768 35876 107824 35932
rect 107824 35876 107828 35932
rect 107764 35872 107828 35876
rect 107844 35932 107908 35936
rect 107844 35876 107848 35932
rect 107848 35876 107904 35932
rect 107904 35876 107908 35932
rect 107844 35872 107908 35876
rect 107924 35932 107988 35936
rect 107924 35876 107928 35932
rect 107928 35876 107984 35932
rect 107984 35876 107988 35932
rect 107924 35872 107988 35876
rect 108004 35932 108068 35936
rect 108004 35876 108008 35932
rect 108008 35876 108064 35932
rect 108064 35876 108068 35932
rect 108004 35872 108068 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 107028 35388 107092 35392
rect 107028 35332 107032 35388
rect 107032 35332 107088 35388
rect 107088 35332 107092 35388
rect 107028 35328 107092 35332
rect 107108 35388 107172 35392
rect 107108 35332 107112 35388
rect 107112 35332 107168 35388
rect 107168 35332 107172 35388
rect 107108 35328 107172 35332
rect 107188 35388 107252 35392
rect 107188 35332 107192 35388
rect 107192 35332 107248 35388
rect 107248 35332 107252 35388
rect 107188 35328 107252 35332
rect 107268 35388 107332 35392
rect 107268 35332 107272 35388
rect 107272 35332 107328 35388
rect 107328 35332 107332 35388
rect 107268 35328 107332 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 107764 34844 107828 34848
rect 107764 34788 107768 34844
rect 107768 34788 107824 34844
rect 107824 34788 107828 34844
rect 107764 34784 107828 34788
rect 107844 34844 107908 34848
rect 107844 34788 107848 34844
rect 107848 34788 107904 34844
rect 107904 34788 107908 34844
rect 107844 34784 107908 34788
rect 107924 34844 107988 34848
rect 107924 34788 107928 34844
rect 107928 34788 107984 34844
rect 107984 34788 107988 34844
rect 107924 34784 107988 34788
rect 108004 34844 108068 34848
rect 108004 34788 108008 34844
rect 108008 34788 108064 34844
rect 108064 34788 108068 34844
rect 108004 34784 108068 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 107028 34300 107092 34304
rect 107028 34244 107032 34300
rect 107032 34244 107088 34300
rect 107088 34244 107092 34300
rect 107028 34240 107092 34244
rect 107108 34300 107172 34304
rect 107108 34244 107112 34300
rect 107112 34244 107168 34300
rect 107168 34244 107172 34300
rect 107108 34240 107172 34244
rect 107188 34300 107252 34304
rect 107188 34244 107192 34300
rect 107192 34244 107248 34300
rect 107248 34244 107252 34300
rect 107188 34240 107252 34244
rect 107268 34300 107332 34304
rect 107268 34244 107272 34300
rect 107272 34244 107328 34300
rect 107328 34244 107332 34300
rect 107268 34240 107332 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 107764 33756 107828 33760
rect 107764 33700 107768 33756
rect 107768 33700 107824 33756
rect 107824 33700 107828 33756
rect 107764 33696 107828 33700
rect 107844 33756 107908 33760
rect 107844 33700 107848 33756
rect 107848 33700 107904 33756
rect 107904 33700 107908 33756
rect 107844 33696 107908 33700
rect 107924 33756 107988 33760
rect 107924 33700 107928 33756
rect 107928 33700 107984 33756
rect 107984 33700 107988 33756
rect 107924 33696 107988 33700
rect 108004 33756 108068 33760
rect 108004 33700 108008 33756
rect 108008 33700 108064 33756
rect 108064 33700 108068 33756
rect 108004 33696 108068 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 107028 33212 107092 33216
rect 107028 33156 107032 33212
rect 107032 33156 107088 33212
rect 107088 33156 107092 33212
rect 107028 33152 107092 33156
rect 107108 33212 107172 33216
rect 107108 33156 107112 33212
rect 107112 33156 107168 33212
rect 107168 33156 107172 33212
rect 107108 33152 107172 33156
rect 107188 33212 107252 33216
rect 107188 33156 107192 33212
rect 107192 33156 107248 33212
rect 107248 33156 107252 33212
rect 107188 33152 107252 33156
rect 107268 33212 107332 33216
rect 107268 33156 107272 33212
rect 107272 33156 107328 33212
rect 107328 33156 107332 33212
rect 107268 33152 107332 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 107764 32668 107828 32672
rect 107764 32612 107768 32668
rect 107768 32612 107824 32668
rect 107824 32612 107828 32668
rect 107764 32608 107828 32612
rect 107844 32668 107908 32672
rect 107844 32612 107848 32668
rect 107848 32612 107904 32668
rect 107904 32612 107908 32668
rect 107844 32608 107908 32612
rect 107924 32668 107988 32672
rect 107924 32612 107928 32668
rect 107928 32612 107984 32668
rect 107984 32612 107988 32668
rect 107924 32608 107988 32612
rect 108004 32668 108068 32672
rect 108004 32612 108008 32668
rect 108008 32612 108064 32668
rect 108064 32612 108068 32668
rect 108004 32608 108068 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 107028 32124 107092 32128
rect 107028 32068 107032 32124
rect 107032 32068 107088 32124
rect 107088 32068 107092 32124
rect 107028 32064 107092 32068
rect 107108 32124 107172 32128
rect 107108 32068 107112 32124
rect 107112 32068 107168 32124
rect 107168 32068 107172 32124
rect 107108 32064 107172 32068
rect 107188 32124 107252 32128
rect 107188 32068 107192 32124
rect 107192 32068 107248 32124
rect 107248 32068 107252 32124
rect 107188 32064 107252 32068
rect 107268 32124 107332 32128
rect 107268 32068 107272 32124
rect 107272 32068 107328 32124
rect 107328 32068 107332 32124
rect 107268 32064 107332 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 107764 31580 107828 31584
rect 107764 31524 107768 31580
rect 107768 31524 107824 31580
rect 107824 31524 107828 31580
rect 107764 31520 107828 31524
rect 107844 31580 107908 31584
rect 107844 31524 107848 31580
rect 107848 31524 107904 31580
rect 107904 31524 107908 31580
rect 107844 31520 107908 31524
rect 107924 31580 107988 31584
rect 107924 31524 107928 31580
rect 107928 31524 107984 31580
rect 107984 31524 107988 31580
rect 107924 31520 107988 31524
rect 108004 31580 108068 31584
rect 108004 31524 108008 31580
rect 108008 31524 108064 31580
rect 108064 31524 108068 31580
rect 108004 31520 108068 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 107028 31036 107092 31040
rect 107028 30980 107032 31036
rect 107032 30980 107088 31036
rect 107088 30980 107092 31036
rect 107028 30976 107092 30980
rect 107108 31036 107172 31040
rect 107108 30980 107112 31036
rect 107112 30980 107168 31036
rect 107168 30980 107172 31036
rect 107108 30976 107172 30980
rect 107188 31036 107252 31040
rect 107188 30980 107192 31036
rect 107192 30980 107248 31036
rect 107248 30980 107252 31036
rect 107188 30976 107252 30980
rect 107268 31036 107332 31040
rect 107268 30980 107272 31036
rect 107272 30980 107328 31036
rect 107328 30980 107332 31036
rect 107268 30976 107332 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 107764 30492 107828 30496
rect 107764 30436 107768 30492
rect 107768 30436 107824 30492
rect 107824 30436 107828 30492
rect 107764 30432 107828 30436
rect 107844 30492 107908 30496
rect 107844 30436 107848 30492
rect 107848 30436 107904 30492
rect 107904 30436 107908 30492
rect 107844 30432 107908 30436
rect 107924 30492 107988 30496
rect 107924 30436 107928 30492
rect 107928 30436 107984 30492
rect 107984 30436 107988 30492
rect 107924 30432 107988 30436
rect 108004 30492 108068 30496
rect 108004 30436 108008 30492
rect 108008 30436 108064 30492
rect 108064 30436 108068 30492
rect 108004 30432 108068 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 107028 29948 107092 29952
rect 107028 29892 107032 29948
rect 107032 29892 107088 29948
rect 107088 29892 107092 29948
rect 107028 29888 107092 29892
rect 107108 29948 107172 29952
rect 107108 29892 107112 29948
rect 107112 29892 107168 29948
rect 107168 29892 107172 29948
rect 107108 29888 107172 29892
rect 107188 29948 107252 29952
rect 107188 29892 107192 29948
rect 107192 29892 107248 29948
rect 107248 29892 107252 29948
rect 107188 29888 107252 29892
rect 107268 29948 107332 29952
rect 107268 29892 107272 29948
rect 107272 29892 107328 29948
rect 107328 29892 107332 29948
rect 107268 29888 107332 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 107764 29404 107828 29408
rect 107764 29348 107768 29404
rect 107768 29348 107824 29404
rect 107824 29348 107828 29404
rect 107764 29344 107828 29348
rect 107844 29404 107908 29408
rect 107844 29348 107848 29404
rect 107848 29348 107904 29404
rect 107904 29348 107908 29404
rect 107844 29344 107908 29348
rect 107924 29404 107988 29408
rect 107924 29348 107928 29404
rect 107928 29348 107984 29404
rect 107984 29348 107988 29404
rect 107924 29344 107988 29348
rect 108004 29404 108068 29408
rect 108004 29348 108008 29404
rect 108008 29348 108064 29404
rect 108064 29348 108068 29404
rect 108004 29344 108068 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 107028 28860 107092 28864
rect 107028 28804 107032 28860
rect 107032 28804 107088 28860
rect 107088 28804 107092 28860
rect 107028 28800 107092 28804
rect 107108 28860 107172 28864
rect 107108 28804 107112 28860
rect 107112 28804 107168 28860
rect 107168 28804 107172 28860
rect 107108 28800 107172 28804
rect 107188 28860 107252 28864
rect 107188 28804 107192 28860
rect 107192 28804 107248 28860
rect 107248 28804 107252 28860
rect 107188 28800 107252 28804
rect 107268 28860 107332 28864
rect 107268 28804 107272 28860
rect 107272 28804 107328 28860
rect 107328 28804 107332 28860
rect 107268 28800 107332 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 107764 28316 107828 28320
rect 107764 28260 107768 28316
rect 107768 28260 107824 28316
rect 107824 28260 107828 28316
rect 107764 28256 107828 28260
rect 107844 28316 107908 28320
rect 107844 28260 107848 28316
rect 107848 28260 107904 28316
rect 107904 28260 107908 28316
rect 107844 28256 107908 28260
rect 107924 28316 107988 28320
rect 107924 28260 107928 28316
rect 107928 28260 107984 28316
rect 107984 28260 107988 28316
rect 107924 28256 107988 28260
rect 108004 28316 108068 28320
rect 108004 28260 108008 28316
rect 108008 28260 108064 28316
rect 108064 28260 108068 28316
rect 108004 28256 108068 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 107028 27772 107092 27776
rect 107028 27716 107032 27772
rect 107032 27716 107088 27772
rect 107088 27716 107092 27772
rect 107028 27712 107092 27716
rect 107108 27772 107172 27776
rect 107108 27716 107112 27772
rect 107112 27716 107168 27772
rect 107168 27716 107172 27772
rect 107108 27712 107172 27716
rect 107188 27772 107252 27776
rect 107188 27716 107192 27772
rect 107192 27716 107248 27772
rect 107248 27716 107252 27772
rect 107188 27712 107252 27716
rect 107268 27772 107332 27776
rect 107268 27716 107272 27772
rect 107272 27716 107328 27772
rect 107328 27716 107332 27772
rect 107268 27712 107332 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 107764 27228 107828 27232
rect 107764 27172 107768 27228
rect 107768 27172 107824 27228
rect 107824 27172 107828 27228
rect 107764 27168 107828 27172
rect 107844 27228 107908 27232
rect 107844 27172 107848 27228
rect 107848 27172 107904 27228
rect 107904 27172 107908 27228
rect 107844 27168 107908 27172
rect 107924 27228 107988 27232
rect 107924 27172 107928 27228
rect 107928 27172 107984 27228
rect 107984 27172 107988 27228
rect 107924 27168 107988 27172
rect 108004 27228 108068 27232
rect 108004 27172 108008 27228
rect 108008 27172 108064 27228
rect 108064 27172 108068 27228
rect 108004 27168 108068 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 107028 26684 107092 26688
rect 107028 26628 107032 26684
rect 107032 26628 107088 26684
rect 107088 26628 107092 26684
rect 107028 26624 107092 26628
rect 107108 26684 107172 26688
rect 107108 26628 107112 26684
rect 107112 26628 107168 26684
rect 107168 26628 107172 26684
rect 107108 26624 107172 26628
rect 107188 26684 107252 26688
rect 107188 26628 107192 26684
rect 107192 26628 107248 26684
rect 107248 26628 107252 26684
rect 107188 26624 107252 26628
rect 107268 26684 107332 26688
rect 107268 26628 107272 26684
rect 107272 26628 107328 26684
rect 107328 26628 107332 26684
rect 107268 26624 107332 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 107764 26140 107828 26144
rect 107764 26084 107768 26140
rect 107768 26084 107824 26140
rect 107824 26084 107828 26140
rect 107764 26080 107828 26084
rect 107844 26140 107908 26144
rect 107844 26084 107848 26140
rect 107848 26084 107904 26140
rect 107904 26084 107908 26140
rect 107844 26080 107908 26084
rect 107924 26140 107988 26144
rect 107924 26084 107928 26140
rect 107928 26084 107984 26140
rect 107984 26084 107988 26140
rect 107924 26080 107988 26084
rect 108004 26140 108068 26144
rect 108004 26084 108008 26140
rect 108008 26084 108064 26140
rect 108064 26084 108068 26140
rect 108004 26080 108068 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 107028 25596 107092 25600
rect 107028 25540 107032 25596
rect 107032 25540 107088 25596
rect 107088 25540 107092 25596
rect 107028 25536 107092 25540
rect 107108 25596 107172 25600
rect 107108 25540 107112 25596
rect 107112 25540 107168 25596
rect 107168 25540 107172 25596
rect 107108 25536 107172 25540
rect 107188 25596 107252 25600
rect 107188 25540 107192 25596
rect 107192 25540 107248 25596
rect 107248 25540 107252 25596
rect 107188 25536 107252 25540
rect 107268 25596 107332 25600
rect 107268 25540 107272 25596
rect 107272 25540 107328 25596
rect 107328 25540 107332 25596
rect 107268 25536 107332 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 107764 25052 107828 25056
rect 107764 24996 107768 25052
rect 107768 24996 107824 25052
rect 107824 24996 107828 25052
rect 107764 24992 107828 24996
rect 107844 25052 107908 25056
rect 107844 24996 107848 25052
rect 107848 24996 107904 25052
rect 107904 24996 107908 25052
rect 107844 24992 107908 24996
rect 107924 25052 107988 25056
rect 107924 24996 107928 25052
rect 107928 24996 107984 25052
rect 107984 24996 107988 25052
rect 107924 24992 107988 24996
rect 108004 25052 108068 25056
rect 108004 24996 108008 25052
rect 108008 24996 108064 25052
rect 108064 24996 108068 25052
rect 108004 24992 108068 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 107028 24508 107092 24512
rect 107028 24452 107032 24508
rect 107032 24452 107088 24508
rect 107088 24452 107092 24508
rect 107028 24448 107092 24452
rect 107108 24508 107172 24512
rect 107108 24452 107112 24508
rect 107112 24452 107168 24508
rect 107168 24452 107172 24508
rect 107108 24448 107172 24452
rect 107188 24508 107252 24512
rect 107188 24452 107192 24508
rect 107192 24452 107248 24508
rect 107248 24452 107252 24508
rect 107188 24448 107252 24452
rect 107268 24508 107332 24512
rect 107268 24452 107272 24508
rect 107272 24452 107328 24508
rect 107328 24452 107332 24508
rect 107268 24448 107332 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 107764 23964 107828 23968
rect 107764 23908 107768 23964
rect 107768 23908 107824 23964
rect 107824 23908 107828 23964
rect 107764 23904 107828 23908
rect 107844 23964 107908 23968
rect 107844 23908 107848 23964
rect 107848 23908 107904 23964
rect 107904 23908 107908 23964
rect 107844 23904 107908 23908
rect 107924 23964 107988 23968
rect 107924 23908 107928 23964
rect 107928 23908 107984 23964
rect 107984 23908 107988 23964
rect 107924 23904 107988 23908
rect 108004 23964 108068 23968
rect 108004 23908 108008 23964
rect 108008 23908 108064 23964
rect 108064 23908 108068 23964
rect 108004 23904 108068 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 107028 23420 107092 23424
rect 107028 23364 107032 23420
rect 107032 23364 107088 23420
rect 107088 23364 107092 23420
rect 107028 23360 107092 23364
rect 107108 23420 107172 23424
rect 107108 23364 107112 23420
rect 107112 23364 107168 23420
rect 107168 23364 107172 23420
rect 107108 23360 107172 23364
rect 107188 23420 107252 23424
rect 107188 23364 107192 23420
rect 107192 23364 107248 23420
rect 107248 23364 107252 23420
rect 107188 23360 107252 23364
rect 107268 23420 107332 23424
rect 107268 23364 107272 23420
rect 107272 23364 107328 23420
rect 107328 23364 107332 23420
rect 107268 23360 107332 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 107764 22876 107828 22880
rect 107764 22820 107768 22876
rect 107768 22820 107824 22876
rect 107824 22820 107828 22876
rect 107764 22816 107828 22820
rect 107844 22876 107908 22880
rect 107844 22820 107848 22876
rect 107848 22820 107904 22876
rect 107904 22820 107908 22876
rect 107844 22816 107908 22820
rect 107924 22876 107988 22880
rect 107924 22820 107928 22876
rect 107928 22820 107984 22876
rect 107984 22820 107988 22876
rect 107924 22816 107988 22820
rect 108004 22876 108068 22880
rect 108004 22820 108008 22876
rect 108008 22820 108064 22876
rect 108064 22820 108068 22876
rect 108004 22816 108068 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 107028 22332 107092 22336
rect 107028 22276 107032 22332
rect 107032 22276 107088 22332
rect 107088 22276 107092 22332
rect 107028 22272 107092 22276
rect 107108 22332 107172 22336
rect 107108 22276 107112 22332
rect 107112 22276 107168 22332
rect 107168 22276 107172 22332
rect 107108 22272 107172 22276
rect 107188 22332 107252 22336
rect 107188 22276 107192 22332
rect 107192 22276 107248 22332
rect 107248 22276 107252 22332
rect 107188 22272 107252 22276
rect 107268 22332 107332 22336
rect 107268 22276 107272 22332
rect 107272 22276 107328 22332
rect 107328 22276 107332 22332
rect 107268 22272 107332 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 107764 21788 107828 21792
rect 107764 21732 107768 21788
rect 107768 21732 107824 21788
rect 107824 21732 107828 21788
rect 107764 21728 107828 21732
rect 107844 21788 107908 21792
rect 107844 21732 107848 21788
rect 107848 21732 107904 21788
rect 107904 21732 107908 21788
rect 107844 21728 107908 21732
rect 107924 21788 107988 21792
rect 107924 21732 107928 21788
rect 107928 21732 107984 21788
rect 107984 21732 107988 21788
rect 107924 21728 107988 21732
rect 108004 21788 108068 21792
rect 108004 21732 108008 21788
rect 108008 21732 108064 21788
rect 108064 21732 108068 21788
rect 108004 21728 108068 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 107028 21244 107092 21248
rect 107028 21188 107032 21244
rect 107032 21188 107088 21244
rect 107088 21188 107092 21244
rect 107028 21184 107092 21188
rect 107108 21244 107172 21248
rect 107108 21188 107112 21244
rect 107112 21188 107168 21244
rect 107168 21188 107172 21244
rect 107108 21184 107172 21188
rect 107188 21244 107252 21248
rect 107188 21188 107192 21244
rect 107192 21188 107248 21244
rect 107248 21188 107252 21244
rect 107188 21184 107252 21188
rect 107268 21244 107332 21248
rect 107268 21188 107272 21244
rect 107272 21188 107328 21244
rect 107328 21188 107332 21244
rect 107268 21184 107332 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 107764 20700 107828 20704
rect 107764 20644 107768 20700
rect 107768 20644 107824 20700
rect 107824 20644 107828 20700
rect 107764 20640 107828 20644
rect 107844 20700 107908 20704
rect 107844 20644 107848 20700
rect 107848 20644 107904 20700
rect 107904 20644 107908 20700
rect 107844 20640 107908 20644
rect 107924 20700 107988 20704
rect 107924 20644 107928 20700
rect 107928 20644 107984 20700
rect 107984 20644 107988 20700
rect 107924 20640 107988 20644
rect 108004 20700 108068 20704
rect 108004 20644 108008 20700
rect 108008 20644 108064 20700
rect 108064 20644 108068 20700
rect 108004 20640 108068 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 107028 20156 107092 20160
rect 107028 20100 107032 20156
rect 107032 20100 107088 20156
rect 107088 20100 107092 20156
rect 107028 20096 107092 20100
rect 107108 20156 107172 20160
rect 107108 20100 107112 20156
rect 107112 20100 107168 20156
rect 107168 20100 107172 20156
rect 107108 20096 107172 20100
rect 107188 20156 107252 20160
rect 107188 20100 107192 20156
rect 107192 20100 107248 20156
rect 107248 20100 107252 20156
rect 107188 20096 107252 20100
rect 107268 20156 107332 20160
rect 107268 20100 107272 20156
rect 107272 20100 107328 20156
rect 107328 20100 107332 20156
rect 107268 20096 107332 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 107764 19612 107828 19616
rect 107764 19556 107768 19612
rect 107768 19556 107824 19612
rect 107824 19556 107828 19612
rect 107764 19552 107828 19556
rect 107844 19612 107908 19616
rect 107844 19556 107848 19612
rect 107848 19556 107904 19612
rect 107904 19556 107908 19612
rect 107844 19552 107908 19556
rect 107924 19612 107988 19616
rect 107924 19556 107928 19612
rect 107928 19556 107984 19612
rect 107984 19556 107988 19612
rect 107924 19552 107988 19556
rect 108004 19612 108068 19616
rect 108004 19556 108008 19612
rect 108008 19556 108064 19612
rect 108064 19556 108068 19612
rect 108004 19552 108068 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 107028 19068 107092 19072
rect 107028 19012 107032 19068
rect 107032 19012 107088 19068
rect 107088 19012 107092 19068
rect 107028 19008 107092 19012
rect 107108 19068 107172 19072
rect 107108 19012 107112 19068
rect 107112 19012 107168 19068
rect 107168 19012 107172 19068
rect 107108 19008 107172 19012
rect 107188 19068 107252 19072
rect 107188 19012 107192 19068
rect 107192 19012 107248 19068
rect 107248 19012 107252 19068
rect 107188 19008 107252 19012
rect 107268 19068 107332 19072
rect 107268 19012 107272 19068
rect 107272 19012 107328 19068
rect 107328 19012 107332 19068
rect 107268 19008 107332 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 107764 18524 107828 18528
rect 107764 18468 107768 18524
rect 107768 18468 107824 18524
rect 107824 18468 107828 18524
rect 107764 18464 107828 18468
rect 107844 18524 107908 18528
rect 107844 18468 107848 18524
rect 107848 18468 107904 18524
rect 107904 18468 107908 18524
rect 107844 18464 107908 18468
rect 107924 18524 107988 18528
rect 107924 18468 107928 18524
rect 107928 18468 107984 18524
rect 107984 18468 107988 18524
rect 107924 18464 107988 18468
rect 108004 18524 108068 18528
rect 108004 18468 108008 18524
rect 108008 18468 108064 18524
rect 108064 18468 108068 18524
rect 108004 18464 108068 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 107028 17980 107092 17984
rect 107028 17924 107032 17980
rect 107032 17924 107088 17980
rect 107088 17924 107092 17980
rect 107028 17920 107092 17924
rect 107108 17980 107172 17984
rect 107108 17924 107112 17980
rect 107112 17924 107168 17980
rect 107168 17924 107172 17980
rect 107108 17920 107172 17924
rect 107188 17980 107252 17984
rect 107188 17924 107192 17980
rect 107192 17924 107248 17980
rect 107248 17924 107252 17980
rect 107188 17920 107252 17924
rect 107268 17980 107332 17984
rect 107268 17924 107272 17980
rect 107272 17924 107328 17980
rect 107328 17924 107332 17980
rect 107268 17920 107332 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 107764 17436 107828 17440
rect 107764 17380 107768 17436
rect 107768 17380 107824 17436
rect 107824 17380 107828 17436
rect 107764 17376 107828 17380
rect 107844 17436 107908 17440
rect 107844 17380 107848 17436
rect 107848 17380 107904 17436
rect 107904 17380 107908 17436
rect 107844 17376 107908 17380
rect 107924 17436 107988 17440
rect 107924 17380 107928 17436
rect 107928 17380 107984 17436
rect 107984 17380 107988 17436
rect 107924 17376 107988 17380
rect 108004 17436 108068 17440
rect 108004 17380 108008 17436
rect 108008 17380 108064 17436
rect 108064 17380 108068 17436
rect 108004 17376 108068 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 107028 16892 107092 16896
rect 107028 16836 107032 16892
rect 107032 16836 107088 16892
rect 107088 16836 107092 16892
rect 107028 16832 107092 16836
rect 107108 16892 107172 16896
rect 107108 16836 107112 16892
rect 107112 16836 107168 16892
rect 107168 16836 107172 16892
rect 107108 16832 107172 16836
rect 107188 16892 107252 16896
rect 107188 16836 107192 16892
rect 107192 16836 107248 16892
rect 107248 16836 107252 16892
rect 107188 16832 107252 16836
rect 107268 16892 107332 16896
rect 107268 16836 107272 16892
rect 107272 16836 107328 16892
rect 107328 16836 107332 16892
rect 107268 16832 107332 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 107764 16348 107828 16352
rect 107764 16292 107768 16348
rect 107768 16292 107824 16348
rect 107824 16292 107828 16348
rect 107764 16288 107828 16292
rect 107844 16348 107908 16352
rect 107844 16292 107848 16348
rect 107848 16292 107904 16348
rect 107904 16292 107908 16348
rect 107844 16288 107908 16292
rect 107924 16348 107988 16352
rect 107924 16292 107928 16348
rect 107928 16292 107984 16348
rect 107984 16292 107988 16348
rect 107924 16288 107988 16292
rect 108004 16348 108068 16352
rect 108004 16292 108008 16348
rect 108008 16292 108064 16348
rect 108064 16292 108068 16348
rect 108004 16288 108068 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 107028 15804 107092 15808
rect 107028 15748 107032 15804
rect 107032 15748 107088 15804
rect 107088 15748 107092 15804
rect 107028 15744 107092 15748
rect 107108 15804 107172 15808
rect 107108 15748 107112 15804
rect 107112 15748 107168 15804
rect 107168 15748 107172 15804
rect 107108 15744 107172 15748
rect 107188 15804 107252 15808
rect 107188 15748 107192 15804
rect 107192 15748 107248 15804
rect 107248 15748 107252 15804
rect 107188 15744 107252 15748
rect 107268 15804 107332 15808
rect 107268 15748 107272 15804
rect 107272 15748 107328 15804
rect 107328 15748 107332 15804
rect 107268 15744 107332 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 107764 15260 107828 15264
rect 107764 15204 107768 15260
rect 107768 15204 107824 15260
rect 107824 15204 107828 15260
rect 107764 15200 107828 15204
rect 107844 15260 107908 15264
rect 107844 15204 107848 15260
rect 107848 15204 107904 15260
rect 107904 15204 107908 15260
rect 107844 15200 107908 15204
rect 107924 15260 107988 15264
rect 107924 15204 107928 15260
rect 107928 15204 107984 15260
rect 107984 15204 107988 15260
rect 107924 15200 107988 15204
rect 108004 15260 108068 15264
rect 108004 15204 108008 15260
rect 108008 15204 108064 15260
rect 108064 15204 108068 15260
rect 108004 15200 108068 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 107028 14716 107092 14720
rect 107028 14660 107032 14716
rect 107032 14660 107088 14716
rect 107088 14660 107092 14716
rect 107028 14656 107092 14660
rect 107108 14716 107172 14720
rect 107108 14660 107112 14716
rect 107112 14660 107168 14716
rect 107168 14660 107172 14716
rect 107108 14656 107172 14660
rect 107188 14716 107252 14720
rect 107188 14660 107192 14716
rect 107192 14660 107248 14716
rect 107248 14660 107252 14716
rect 107188 14656 107252 14660
rect 107268 14716 107332 14720
rect 107268 14660 107272 14716
rect 107272 14660 107328 14716
rect 107328 14660 107332 14716
rect 107268 14656 107332 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 107764 14172 107828 14176
rect 107764 14116 107768 14172
rect 107768 14116 107824 14172
rect 107824 14116 107828 14172
rect 107764 14112 107828 14116
rect 107844 14172 107908 14176
rect 107844 14116 107848 14172
rect 107848 14116 107904 14172
rect 107904 14116 107908 14172
rect 107844 14112 107908 14116
rect 107924 14172 107988 14176
rect 107924 14116 107928 14172
rect 107928 14116 107984 14172
rect 107984 14116 107988 14172
rect 107924 14112 107988 14116
rect 108004 14172 108068 14176
rect 108004 14116 108008 14172
rect 108008 14116 108064 14172
rect 108064 14116 108068 14172
rect 108004 14112 108068 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 107028 13628 107092 13632
rect 107028 13572 107032 13628
rect 107032 13572 107088 13628
rect 107088 13572 107092 13628
rect 107028 13568 107092 13572
rect 107108 13628 107172 13632
rect 107108 13572 107112 13628
rect 107112 13572 107168 13628
rect 107168 13572 107172 13628
rect 107108 13568 107172 13572
rect 107188 13628 107252 13632
rect 107188 13572 107192 13628
rect 107192 13572 107248 13628
rect 107248 13572 107252 13628
rect 107188 13568 107252 13572
rect 107268 13628 107332 13632
rect 107268 13572 107272 13628
rect 107272 13572 107328 13628
rect 107328 13572 107332 13628
rect 107268 13568 107332 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 107764 13084 107828 13088
rect 107764 13028 107768 13084
rect 107768 13028 107824 13084
rect 107824 13028 107828 13084
rect 107764 13024 107828 13028
rect 107844 13084 107908 13088
rect 107844 13028 107848 13084
rect 107848 13028 107904 13084
rect 107904 13028 107908 13084
rect 107844 13024 107908 13028
rect 107924 13084 107988 13088
rect 107924 13028 107928 13084
rect 107928 13028 107984 13084
rect 107984 13028 107988 13084
rect 107924 13024 107988 13028
rect 108004 13084 108068 13088
rect 108004 13028 108008 13084
rect 108008 13028 108064 13084
rect 108064 13028 108068 13084
rect 108004 13024 108068 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 107028 12540 107092 12544
rect 107028 12484 107032 12540
rect 107032 12484 107088 12540
rect 107088 12484 107092 12540
rect 107028 12480 107092 12484
rect 107108 12540 107172 12544
rect 107108 12484 107112 12540
rect 107112 12484 107168 12540
rect 107168 12484 107172 12540
rect 107108 12480 107172 12484
rect 107188 12540 107252 12544
rect 107188 12484 107192 12540
rect 107192 12484 107248 12540
rect 107248 12484 107252 12540
rect 107188 12480 107252 12484
rect 107268 12540 107332 12544
rect 107268 12484 107272 12540
rect 107272 12484 107328 12540
rect 107328 12484 107332 12540
rect 107268 12480 107332 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 107764 11996 107828 12000
rect 107764 11940 107768 11996
rect 107768 11940 107824 11996
rect 107824 11940 107828 11996
rect 107764 11936 107828 11940
rect 107844 11996 107908 12000
rect 107844 11940 107848 11996
rect 107848 11940 107904 11996
rect 107904 11940 107908 11996
rect 107844 11936 107908 11940
rect 107924 11996 107988 12000
rect 107924 11940 107928 11996
rect 107928 11940 107984 11996
rect 107984 11940 107988 11996
rect 107924 11936 107988 11940
rect 108004 11996 108068 12000
rect 108004 11940 108008 11996
rect 108008 11940 108064 11996
rect 108064 11940 108068 11996
rect 108004 11936 108068 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 107028 11452 107092 11456
rect 107028 11396 107032 11452
rect 107032 11396 107088 11452
rect 107088 11396 107092 11452
rect 107028 11392 107092 11396
rect 107108 11452 107172 11456
rect 107108 11396 107112 11452
rect 107112 11396 107168 11452
rect 107168 11396 107172 11452
rect 107108 11392 107172 11396
rect 107188 11452 107252 11456
rect 107188 11396 107192 11452
rect 107192 11396 107248 11452
rect 107248 11396 107252 11452
rect 107188 11392 107252 11396
rect 107268 11452 107332 11456
rect 107268 11396 107272 11452
rect 107272 11396 107328 11452
rect 107328 11396 107332 11452
rect 107268 11392 107332 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 107764 10908 107828 10912
rect 107764 10852 107768 10908
rect 107768 10852 107824 10908
rect 107824 10852 107828 10908
rect 107764 10848 107828 10852
rect 107844 10908 107908 10912
rect 107844 10852 107848 10908
rect 107848 10852 107904 10908
rect 107904 10852 107908 10908
rect 107844 10848 107908 10852
rect 107924 10908 107988 10912
rect 107924 10852 107928 10908
rect 107928 10852 107984 10908
rect 107984 10852 107988 10908
rect 107924 10848 107988 10852
rect 108004 10908 108068 10912
rect 108004 10852 108008 10908
rect 108008 10852 108064 10908
rect 108064 10852 108068 10908
rect 108004 10848 108068 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 107028 10364 107092 10368
rect 107028 10308 107032 10364
rect 107032 10308 107088 10364
rect 107088 10308 107092 10364
rect 107028 10304 107092 10308
rect 107108 10364 107172 10368
rect 107108 10308 107112 10364
rect 107112 10308 107168 10364
rect 107168 10308 107172 10364
rect 107108 10304 107172 10308
rect 107188 10364 107252 10368
rect 107188 10308 107192 10364
rect 107192 10308 107248 10364
rect 107248 10308 107252 10364
rect 107188 10304 107252 10308
rect 107268 10364 107332 10368
rect 107268 10308 107272 10364
rect 107272 10308 107328 10364
rect 107328 10308 107332 10364
rect 107268 10304 107332 10308
rect 16058 9888 16122 9892
rect 16058 9832 16082 9888
rect 16082 9832 16122 9888
rect 16058 9828 16122 9832
rect 90404 9888 90468 9892
rect 90404 9832 90418 9888
rect 90418 9832 90468 9888
rect 90404 9828 90468 9832
rect 90956 9828 91020 9892
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 107764 9820 107828 9824
rect 107764 9764 107768 9820
rect 107768 9764 107824 9820
rect 107824 9764 107828 9820
rect 107764 9760 107828 9764
rect 107844 9820 107908 9824
rect 107844 9764 107848 9820
rect 107848 9764 107904 9820
rect 107904 9764 107908 9820
rect 107844 9760 107908 9764
rect 107924 9820 107988 9824
rect 107924 9764 107928 9820
rect 107928 9764 107984 9820
rect 107984 9764 107988 9820
rect 107924 9760 107988 9764
rect 108004 9820 108068 9824
rect 108004 9764 108008 9820
rect 108008 9764 108064 9820
rect 108064 9764 108068 9820
rect 108004 9760 108068 9764
rect 31614 9752 31678 9756
rect 31614 9696 31630 9752
rect 31630 9696 31678 9752
rect 31614 9692 31678 9696
rect 23438 9616 23502 9620
rect 23438 9560 23478 9616
rect 23478 9560 23502 9616
rect 23438 9556 23502 9560
rect 30446 9616 30510 9620
rect 30446 9560 30470 9616
rect 30470 9560 30510 9616
rect 30446 9556 30510 9560
rect 90680 9480 90744 9484
rect 90680 9424 90730 9480
rect 90730 9424 90744 9480
rect 90680 9420 90744 9424
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 107028 9276 107092 9280
rect 107028 9220 107032 9276
rect 107032 9220 107088 9276
rect 107088 9220 107092 9276
rect 107028 9216 107092 9220
rect 107108 9276 107172 9280
rect 107108 9220 107112 9276
rect 107112 9220 107168 9276
rect 107168 9220 107172 9276
rect 107108 9216 107172 9220
rect 107188 9276 107252 9280
rect 107188 9220 107192 9276
rect 107192 9220 107248 9276
rect 107248 9220 107252 9276
rect 107188 9216 107252 9220
rect 107268 9276 107332 9280
rect 107268 9220 107272 9276
rect 107272 9220 107328 9276
rect 107328 9220 107332 9276
rect 107268 9216 107332 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 107764 8732 107828 8736
rect 107764 8676 107768 8732
rect 107768 8676 107824 8732
rect 107824 8676 107828 8732
rect 107764 8672 107828 8676
rect 107844 8732 107908 8736
rect 107844 8676 107848 8732
rect 107848 8676 107904 8732
rect 107904 8676 107908 8732
rect 107844 8672 107908 8676
rect 107924 8732 107988 8736
rect 107924 8676 107928 8732
rect 107928 8676 107984 8732
rect 107984 8676 107988 8732
rect 107924 8672 107988 8676
rect 108004 8732 108068 8736
rect 108004 8676 108008 8732
rect 108008 8676 108064 8732
rect 108064 8676 108068 8732
rect 108004 8672 108068 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 107028 8188 107092 8192
rect 107028 8132 107032 8188
rect 107032 8132 107088 8188
rect 107088 8132 107092 8188
rect 107028 8128 107092 8132
rect 107108 8188 107172 8192
rect 107108 8132 107112 8188
rect 107112 8132 107168 8188
rect 107168 8132 107172 8188
rect 107108 8128 107172 8132
rect 107188 8188 107252 8192
rect 107188 8132 107192 8188
rect 107192 8132 107248 8188
rect 107248 8132 107252 8188
rect 107188 8128 107252 8132
rect 107268 8188 107332 8192
rect 107268 8132 107272 8188
rect 107272 8132 107328 8188
rect 107328 8132 107332 8188
rect 107268 8128 107332 8132
rect 25820 8120 25884 8124
rect 25820 8064 25834 8120
rect 25834 8064 25884 8120
rect 25820 8060 25884 8064
rect 29316 8060 29380 8124
rect 32812 8120 32876 8124
rect 32812 8064 32862 8120
rect 32862 8064 32876 8120
rect 32812 8060 32876 8064
rect 35204 8120 35268 8124
rect 35204 8064 35254 8120
rect 35254 8064 35268 8120
rect 35204 8060 35268 8064
rect 38700 8120 38764 8124
rect 38700 8064 38714 8120
rect 38714 8064 38764 8120
rect 38700 8060 38764 8064
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 66316 7644 66380 7648
rect 66316 7588 66320 7644
rect 66320 7588 66376 7644
rect 66376 7588 66380 7644
rect 66316 7584 66380 7588
rect 66396 7644 66460 7648
rect 66396 7588 66400 7644
rect 66400 7588 66456 7644
rect 66456 7588 66460 7644
rect 66396 7584 66460 7588
rect 66476 7644 66540 7648
rect 66476 7588 66480 7644
rect 66480 7588 66536 7644
rect 66536 7588 66540 7644
rect 66476 7584 66540 7588
rect 66556 7644 66620 7648
rect 66556 7588 66560 7644
rect 66560 7588 66616 7644
rect 66616 7588 66620 7644
rect 66556 7584 66620 7588
rect 97036 7644 97100 7648
rect 97036 7588 97040 7644
rect 97040 7588 97096 7644
rect 97096 7588 97100 7644
rect 97036 7584 97100 7588
rect 97116 7644 97180 7648
rect 97116 7588 97120 7644
rect 97120 7588 97176 7644
rect 97176 7588 97180 7644
rect 97116 7584 97180 7588
rect 97196 7644 97260 7648
rect 97196 7588 97200 7644
rect 97200 7588 97256 7644
rect 97256 7588 97260 7644
rect 97196 7584 97260 7588
rect 97276 7644 97340 7648
rect 97276 7588 97280 7644
rect 97280 7588 97336 7644
rect 97336 7588 97340 7644
rect 97276 7584 97340 7588
rect 107764 7644 107828 7648
rect 107764 7588 107768 7644
rect 107768 7588 107824 7644
rect 107824 7588 107828 7644
rect 107764 7584 107828 7588
rect 107844 7644 107908 7648
rect 107844 7588 107848 7644
rect 107848 7588 107904 7644
rect 107904 7588 107908 7644
rect 107844 7584 107908 7588
rect 107924 7644 107988 7648
rect 107924 7588 107928 7644
rect 107928 7588 107984 7644
rect 107984 7588 107988 7644
rect 107924 7584 107988 7588
rect 108004 7644 108068 7648
rect 108004 7588 108008 7644
rect 108008 7588 108064 7644
rect 108064 7588 108068 7644
rect 108004 7584 108068 7588
rect 24716 7576 24780 7580
rect 24716 7520 24730 7576
rect 24730 7520 24780 7576
rect 24716 7516 24780 7520
rect 26924 7576 26988 7580
rect 26924 7520 26974 7576
rect 26974 7520 26988 7576
rect 26924 7516 26988 7520
rect 28212 7576 28276 7580
rect 28212 7520 28262 7576
rect 28262 7520 28276 7576
rect 28212 7516 28276 7520
rect 33916 7576 33980 7580
rect 33916 7520 33966 7576
rect 33966 7520 33980 7576
rect 33916 7516 33980 7520
rect 36308 7576 36372 7580
rect 36308 7520 36358 7576
rect 36358 7520 36372 7576
rect 36308 7516 36372 7520
rect 37412 7576 37476 7580
rect 37412 7520 37462 7576
rect 37462 7520 37476 7576
rect 37412 7516 37476 7520
rect 39804 7576 39868 7580
rect 39804 7520 39854 7576
rect 39854 7520 39868 7576
rect 39804 7516 39868 7520
rect 40908 7516 40972 7580
rect 42196 7576 42260 7580
rect 42196 7520 42210 7576
rect 42210 7520 42260 7576
rect 42196 7516 42260 7520
rect 43300 7576 43364 7580
rect 43300 7520 43350 7576
rect 43350 7520 43364 7576
rect 43300 7516 43364 7520
rect 90404 7516 90468 7580
rect 90956 7576 91020 7580
rect 90956 7520 91006 7576
rect 91006 7520 91020 7576
rect 90956 7516 91020 7520
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 107028 7100 107092 7104
rect 107028 7044 107032 7100
rect 107032 7044 107088 7100
rect 107088 7044 107092 7100
rect 107028 7040 107092 7044
rect 107108 7100 107172 7104
rect 107108 7044 107112 7100
rect 107112 7044 107168 7100
rect 107168 7044 107172 7100
rect 107108 7040 107172 7044
rect 107188 7100 107252 7104
rect 107188 7044 107192 7100
rect 107192 7044 107248 7100
rect 107248 7044 107252 7100
rect 107188 7040 107252 7044
rect 107268 7100 107332 7104
rect 107268 7044 107272 7100
rect 107272 7044 107328 7100
rect 107328 7044 107332 7100
rect 107268 7040 107332 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 66316 6556 66380 6560
rect 66316 6500 66320 6556
rect 66320 6500 66376 6556
rect 66376 6500 66380 6556
rect 66316 6496 66380 6500
rect 66396 6556 66460 6560
rect 66396 6500 66400 6556
rect 66400 6500 66456 6556
rect 66456 6500 66460 6556
rect 66396 6496 66460 6500
rect 66476 6556 66540 6560
rect 66476 6500 66480 6556
rect 66480 6500 66536 6556
rect 66536 6500 66540 6556
rect 66476 6496 66540 6500
rect 66556 6556 66620 6560
rect 66556 6500 66560 6556
rect 66560 6500 66616 6556
rect 66616 6500 66620 6556
rect 66556 6496 66620 6500
rect 97036 6556 97100 6560
rect 97036 6500 97040 6556
rect 97040 6500 97096 6556
rect 97096 6500 97100 6556
rect 97036 6496 97100 6500
rect 97116 6556 97180 6560
rect 97116 6500 97120 6556
rect 97120 6500 97176 6556
rect 97176 6500 97180 6556
rect 97116 6496 97180 6500
rect 97196 6556 97260 6560
rect 97196 6500 97200 6556
rect 97200 6500 97256 6556
rect 97256 6500 97260 6556
rect 97196 6496 97260 6500
rect 97276 6556 97340 6560
rect 97276 6500 97280 6556
rect 97280 6500 97336 6556
rect 97336 6500 97340 6556
rect 97276 6496 97340 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 66316 5468 66380 5472
rect 66316 5412 66320 5468
rect 66320 5412 66376 5468
rect 66376 5412 66380 5468
rect 66316 5408 66380 5412
rect 66396 5468 66460 5472
rect 66396 5412 66400 5468
rect 66400 5412 66456 5468
rect 66456 5412 66460 5468
rect 66396 5408 66460 5412
rect 66476 5468 66540 5472
rect 66476 5412 66480 5468
rect 66480 5412 66536 5468
rect 66536 5412 66540 5468
rect 66476 5408 66540 5412
rect 66556 5468 66620 5472
rect 66556 5412 66560 5468
rect 66560 5412 66616 5468
rect 66616 5412 66620 5468
rect 66556 5408 66620 5412
rect 97036 5468 97100 5472
rect 97036 5412 97040 5468
rect 97040 5412 97096 5468
rect 97096 5412 97100 5468
rect 97036 5408 97100 5412
rect 97116 5468 97180 5472
rect 97116 5412 97120 5468
rect 97120 5412 97176 5468
rect 97176 5412 97180 5468
rect 97116 5408 97180 5412
rect 97196 5468 97260 5472
rect 97196 5412 97200 5468
rect 97200 5412 97256 5468
rect 97256 5412 97260 5468
rect 97196 5408 97260 5412
rect 97276 5468 97340 5472
rect 97276 5412 97280 5468
rect 97280 5412 97336 5468
rect 97336 5412 97340 5468
rect 97276 5408 97340 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 66316 4380 66380 4384
rect 66316 4324 66320 4380
rect 66320 4324 66376 4380
rect 66376 4324 66380 4380
rect 66316 4320 66380 4324
rect 66396 4380 66460 4384
rect 66396 4324 66400 4380
rect 66400 4324 66456 4380
rect 66456 4324 66460 4380
rect 66396 4320 66460 4324
rect 66476 4380 66540 4384
rect 66476 4324 66480 4380
rect 66480 4324 66536 4380
rect 66536 4324 66540 4380
rect 66476 4320 66540 4324
rect 66556 4380 66620 4384
rect 66556 4324 66560 4380
rect 66560 4324 66616 4380
rect 66616 4324 66620 4380
rect 66556 4320 66620 4324
rect 97036 4380 97100 4384
rect 97036 4324 97040 4380
rect 97040 4324 97096 4380
rect 97096 4324 97100 4380
rect 97036 4320 97100 4324
rect 97116 4380 97180 4384
rect 97116 4324 97120 4380
rect 97120 4324 97176 4380
rect 97176 4324 97180 4380
rect 97116 4320 97180 4324
rect 97196 4380 97260 4384
rect 97196 4324 97200 4380
rect 97200 4324 97256 4380
rect 97256 4324 97260 4380
rect 97196 4320 97260 4324
rect 97276 4380 97340 4384
rect 97276 4324 97280 4380
rect 97280 4324 97336 4380
rect 97336 4324 97340 4380
rect 97276 4320 97340 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 66316 3292 66380 3296
rect 66316 3236 66320 3292
rect 66320 3236 66376 3292
rect 66376 3236 66380 3292
rect 66316 3232 66380 3236
rect 66396 3292 66460 3296
rect 66396 3236 66400 3292
rect 66400 3236 66456 3292
rect 66456 3236 66460 3292
rect 66396 3232 66460 3236
rect 66476 3292 66540 3296
rect 66476 3236 66480 3292
rect 66480 3236 66536 3292
rect 66536 3236 66540 3292
rect 66476 3232 66540 3236
rect 66556 3292 66620 3296
rect 66556 3236 66560 3292
rect 66560 3236 66616 3292
rect 66616 3236 66620 3292
rect 66556 3232 66620 3236
rect 97036 3292 97100 3296
rect 97036 3236 97040 3292
rect 97040 3236 97096 3292
rect 97096 3236 97100 3292
rect 97036 3232 97100 3236
rect 97116 3292 97180 3296
rect 97116 3236 97120 3292
rect 97120 3236 97176 3292
rect 97176 3236 97180 3292
rect 97116 3232 97180 3236
rect 97196 3292 97260 3296
rect 97196 3236 97200 3292
rect 97200 3236 97256 3292
rect 97256 3236 97260 3292
rect 97196 3232 97260 3236
rect 97276 3292 97340 3296
rect 97276 3236 97280 3292
rect 97280 3236 97336 3292
rect 97336 3236 97340 3292
rect 97276 3232 97340 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
rect 66316 2204 66380 2208
rect 66316 2148 66320 2204
rect 66320 2148 66376 2204
rect 66376 2148 66380 2204
rect 66316 2144 66380 2148
rect 66396 2204 66460 2208
rect 66396 2148 66400 2204
rect 66400 2148 66456 2204
rect 66456 2148 66460 2204
rect 66396 2144 66460 2148
rect 66476 2204 66540 2208
rect 66476 2148 66480 2204
rect 66480 2148 66536 2204
rect 66536 2148 66540 2204
rect 66476 2144 66540 2148
rect 66556 2204 66620 2208
rect 66556 2148 66560 2204
rect 66560 2148 66616 2204
rect 66616 2148 66620 2204
rect 66556 2144 66620 2148
rect 97036 2204 97100 2208
rect 97036 2148 97040 2204
rect 97040 2148 97096 2204
rect 97096 2148 97100 2204
rect 97036 2144 97100 2148
rect 97116 2204 97180 2208
rect 97116 2148 97120 2204
rect 97120 2148 97176 2204
rect 97176 2148 97180 2204
rect 97116 2144 97180 2148
rect 97196 2204 97260 2208
rect 97196 2148 97200 2204
rect 97200 2148 97256 2204
rect 97256 2148 97260 2204
rect 97196 2144 97260 2148
rect 97276 2204 97340 2208
rect 97276 2148 97280 2204
rect 97280 2148 97336 2204
rect 97336 2148 97340 2204
rect 97276 2144 97340 2148
<< metal4 >>
rect 4208 71296 4528 71856
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66896 4296 66944
rect 4360 66896 4376 66944
rect 4440 66896 4456 66944
rect 4520 66880 4528 66944
rect 4208 66660 4250 66880
rect 4486 66660 4528 66880
rect 4208 65856 4528 66660
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 71840 5188 71856
rect 4868 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5188 71840
rect 4868 70752 5188 71776
rect 4868 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5188 70752
rect 4868 69664 5188 70688
rect 4868 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5188 69664
rect 4868 68576 5188 69600
rect 4868 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5188 68576
rect 4868 67556 5188 68512
rect 4868 67488 4910 67556
rect 5146 67488 5188 67556
rect 4868 67424 4876 67488
rect 5180 67424 5188 67488
rect 4868 67320 4910 67424
rect 5146 67320 5188 67424
rect 4868 66400 5188 67320
rect 4868 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5188 66400
rect 4868 65312 5188 66336
rect 34928 71296 35248 71856
rect 34928 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35248 71296
rect 34928 70208 35248 71232
rect 34928 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35248 70208
rect 34928 69120 35248 70144
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66896 35016 66944
rect 35080 66896 35096 66944
rect 35160 66896 35176 66944
rect 35240 66880 35248 66944
rect 34928 66660 34970 66880
rect 35206 66660 35248 66880
rect 34928 65856 35248 66660
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 65650 35248 65792
rect 35588 71840 35908 71856
rect 35588 71776 35596 71840
rect 35660 71776 35676 71840
rect 35740 71776 35756 71840
rect 35820 71776 35836 71840
rect 35900 71776 35908 71840
rect 35588 70752 35908 71776
rect 35588 70688 35596 70752
rect 35660 70688 35676 70752
rect 35740 70688 35756 70752
rect 35820 70688 35836 70752
rect 35900 70688 35908 70752
rect 35588 69664 35908 70688
rect 35588 69600 35596 69664
rect 35660 69600 35676 69664
rect 35740 69600 35756 69664
rect 35820 69600 35836 69664
rect 35900 69600 35908 69664
rect 35588 68576 35908 69600
rect 35588 68512 35596 68576
rect 35660 68512 35676 68576
rect 35740 68512 35756 68576
rect 35820 68512 35836 68576
rect 35900 68512 35908 68576
rect 35588 67556 35908 68512
rect 35588 67488 35630 67556
rect 35866 67488 35908 67556
rect 35588 67424 35596 67488
rect 35900 67424 35908 67488
rect 35588 67320 35630 67424
rect 35866 67320 35908 67424
rect 35588 66400 35908 67320
rect 65648 71296 65968 71856
rect 65648 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65968 71296
rect 65648 70208 65968 71232
rect 65648 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65968 70208
rect 65648 69120 65968 70144
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66896 65736 66944
rect 65800 66896 65816 66944
rect 65880 66896 65896 66944
rect 65960 66880 65968 66944
rect 51027 66740 51093 66741
rect 51027 66676 51028 66740
rect 51092 66676 51093 66740
rect 51027 66675 51093 66676
rect 48635 66468 48701 66469
rect 48635 66404 48636 66468
rect 48700 66404 48701 66468
rect 48635 66403 48701 66404
rect 35588 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35908 66400
rect 35588 65650 35908 66336
rect 46059 66332 46125 66333
rect 46059 66268 46060 66332
rect 46124 66268 46125 66332
rect 46059 66267 46125 66268
rect 4868 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5188 65312
rect 4868 64224 5188 65248
rect 4868 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5188 64224
rect 4868 63136 5188 64160
rect 36074 64156 36140 64157
rect 36074 64092 36075 64156
rect 36139 64092 36140 64156
rect 36074 64091 36140 64092
rect 43575 64156 43641 64157
rect 43575 64092 43576 64156
rect 43640 64092 43641 64156
rect 43575 64091 43641 64092
rect 36077 63676 36137 64091
rect 41066 64020 41132 64021
rect 41066 63956 41067 64020
rect 41131 63956 41132 64020
rect 41066 63955 41132 63956
rect 38570 63884 38636 63885
rect 38570 63820 38571 63884
rect 38635 63820 38636 63884
rect 38570 63819 38636 63820
rect 38573 63676 38633 63819
rect 41069 63676 41129 63955
rect 43578 63676 43638 64091
rect 46062 63676 46122 66267
rect 48638 64290 48698 66403
rect 48557 64230 48698 64290
rect 51030 64290 51090 66675
rect 65648 66660 65690 66880
rect 65926 66660 65968 66880
rect 55995 66468 56061 66469
rect 55995 66404 55996 66468
rect 56060 66404 56061 66468
rect 55995 66403 56061 66404
rect 61147 66468 61213 66469
rect 61147 66404 61148 66468
rect 61212 66404 61213 66468
rect 61147 66403 61213 66404
rect 55998 64290 56058 66403
rect 58571 66332 58637 66333
rect 58571 66268 58572 66332
rect 58636 66268 58637 66332
rect 58571 66267 58637 66268
rect 58574 64290 58634 66267
rect 61150 64290 61210 66403
rect 65648 65856 65968 66660
rect 66308 71840 66628 71856
rect 66308 71776 66316 71840
rect 66380 71776 66396 71840
rect 66460 71776 66476 71840
rect 66540 71776 66556 71840
rect 66620 71776 66628 71840
rect 66308 70752 66628 71776
rect 66308 70688 66316 70752
rect 66380 70688 66396 70752
rect 66460 70688 66476 70752
rect 66540 70688 66556 70752
rect 66620 70688 66628 70752
rect 66308 69664 66628 70688
rect 66308 69600 66316 69664
rect 66380 69600 66396 69664
rect 66460 69600 66476 69664
rect 66540 69600 66556 69664
rect 66620 69600 66628 69664
rect 66308 68576 66628 69600
rect 66308 68512 66316 68576
rect 66380 68512 66396 68576
rect 66460 68512 66476 68576
rect 66540 68512 66556 68576
rect 66620 68512 66628 68576
rect 66308 67556 66628 68512
rect 66308 67488 66350 67556
rect 66586 67488 66628 67556
rect 66308 67424 66316 67488
rect 66620 67424 66628 67488
rect 66308 67320 66350 67424
rect 66586 67320 66628 67424
rect 66115 66604 66181 66605
rect 66115 66540 66116 66604
rect 66180 66540 66181 66604
rect 66115 66539 66181 66540
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 65776 65968 65792
rect 63539 65516 63605 65517
rect 63539 65452 63540 65516
rect 63604 65452 63605 65516
rect 63539 65451 63605 65452
rect 51030 64230 51113 64290
rect 55998 64230 56105 64290
rect 48557 63676 48617 64230
rect 51053 63676 51113 64230
rect 53546 63884 53612 63885
rect 53546 63820 53547 63884
rect 53611 63820 53612 63884
rect 53546 63819 53612 63820
rect 53549 63676 53609 63819
rect 56045 63676 56105 64230
rect 58541 64230 58634 64290
rect 61058 64230 61210 64290
rect 58541 63676 58601 64230
rect 61058 63676 61118 64230
rect 63542 63676 63602 65451
rect 66118 64290 66178 66539
rect 66308 66400 66628 67320
rect 66308 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66628 66400
rect 66308 65650 66628 66336
rect 96368 71296 96688 71856
rect 96368 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96688 71296
rect 96368 70208 96688 71232
rect 96368 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96688 70208
rect 96368 69120 96688 70144
rect 96368 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96688 69120
rect 96368 68032 96688 69056
rect 96368 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96688 68032
rect 96368 66944 96688 67968
rect 96368 66880 96376 66944
rect 96440 66896 96456 66944
rect 96520 66896 96536 66944
rect 96600 66896 96616 66944
rect 96680 66880 96688 66944
rect 96368 66660 96410 66880
rect 96646 66660 96688 66880
rect 96368 65856 96688 66660
rect 96368 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96688 65856
rect 96368 65650 96688 65792
rect 97028 71840 97348 71856
rect 97028 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97348 71840
rect 97028 70752 97348 71776
rect 97028 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97348 70752
rect 97028 69664 97348 70688
rect 97028 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97348 69664
rect 97028 68576 97348 69600
rect 97028 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97348 68576
rect 97028 67556 97348 68512
rect 97028 67488 97070 67556
rect 97306 67488 97348 67556
rect 97028 67424 97036 67488
rect 97340 67424 97348 67488
rect 97028 67320 97070 67424
rect 97306 67320 97348 67424
rect 97028 66400 97348 67320
rect 97028 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97348 66400
rect 97028 65650 97348 66336
rect 107020 65856 107340 66416
rect 107020 65792 107028 65856
rect 107092 65792 107108 65856
rect 107172 65792 107188 65856
rect 107252 65792 107268 65856
rect 107332 65792 107340 65856
rect 68507 65380 68573 65381
rect 68507 65316 68508 65380
rect 68572 65316 68573 65380
rect 68507 65315 68573 65316
rect 73475 65380 73541 65381
rect 73475 65316 73476 65380
rect 73540 65316 73541 65380
rect 73475 65315 73541 65316
rect 87275 65380 87341 65381
rect 87275 65316 87276 65380
rect 87340 65316 87341 65380
rect 87275 65315 87341 65316
rect 66029 64230 66178 64290
rect 66029 63676 66089 64230
rect 68510 63676 68570 65315
rect 71083 65108 71149 65109
rect 71083 65044 71084 65108
rect 71148 65044 71149 65108
rect 71083 65043 71149 65044
rect 71086 64290 71146 65043
rect 71021 64230 71146 64290
rect 73478 64290 73538 65315
rect 87278 64290 87338 65315
rect 107020 64768 107340 65792
rect 107020 64704 107028 64768
rect 107092 64704 107108 64768
rect 107172 64704 107188 64768
rect 107252 64704 107268 64768
rect 107332 64704 107340 64768
rect 73478 64230 73577 64290
rect 87278 64230 87372 64290
rect 71021 63676 71081 64230
rect 73517 63676 73577 64230
rect 87312 64157 87372 64230
rect 87309 64156 87375 64157
rect 87309 64092 87310 64156
rect 87374 64092 87375 64156
rect 87309 64091 87375 64092
rect 86141 64020 86207 64021
rect 86141 63956 86142 64020
rect 86206 63956 86207 64020
rect 86141 63955 86207 63956
rect 86144 63676 86204 63955
rect 87312 63676 87372 64091
rect 95857 63884 95923 63885
rect 95857 63820 95858 63884
rect 95922 63820 95923 63884
rect 95857 63819 95923 63820
rect 95860 63676 95920 63819
rect 107020 63680 107340 64704
rect 4868 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5188 63136
rect 4868 62048 5188 63072
rect 4868 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5188 62048
rect 4868 60960 5188 61984
rect 4868 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5188 60960
rect 4868 59872 5188 60896
rect 4868 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5188 59872
rect 4868 58784 5188 59808
rect 4868 58720 4876 58784
rect 4940 58720 4956 58784
rect 5020 58720 5036 58784
rect 5100 58720 5116 58784
rect 5180 58720 5188 58784
rect 4868 57696 5188 58720
rect 4868 57632 4876 57696
rect 4940 57632 4956 57696
rect 5020 57632 5036 57696
rect 5100 57632 5116 57696
rect 5180 57632 5188 57696
rect 4868 56608 5188 57632
rect 4868 56544 4876 56608
rect 4940 56544 4956 56608
rect 5020 56544 5036 56608
rect 5100 56544 5116 56608
rect 5180 56544 5188 56608
rect 4868 55520 5188 56544
rect 4868 55456 4876 55520
rect 4940 55456 4956 55520
rect 5020 55456 5036 55520
rect 5100 55456 5116 55520
rect 5180 55456 5188 55520
rect 4868 54432 5188 55456
rect 4868 54368 4876 54432
rect 4940 54368 4956 54432
rect 5020 54368 5036 54432
rect 5100 54368 5116 54432
rect 5180 54368 5188 54432
rect 4868 53344 5188 54368
rect 4868 53280 4876 53344
rect 4940 53280 4956 53344
rect 5020 53280 5036 53344
rect 5100 53280 5116 53344
rect 5180 53280 5188 53344
rect 4868 52256 5188 53280
rect 4868 52192 4876 52256
rect 4940 52192 4956 52256
rect 5020 52192 5036 52256
rect 5100 52192 5116 52256
rect 5180 52192 5188 52256
rect 4868 51168 5188 52192
rect 4868 51104 4876 51168
rect 4940 51104 4956 51168
rect 5020 51104 5036 51168
rect 5100 51104 5116 51168
rect 5180 51104 5188 51168
rect 4868 50080 5188 51104
rect 4868 50016 4876 50080
rect 4940 50016 4956 50080
rect 5020 50016 5036 50080
rect 5100 50016 5116 50080
rect 5180 50016 5188 50080
rect 4868 48992 5188 50016
rect 4868 48928 4876 48992
rect 4940 48928 4956 48992
rect 5020 48928 5036 48992
rect 5100 48928 5116 48992
rect 5180 48928 5188 48992
rect 4868 47904 5188 48928
rect 4868 47840 4876 47904
rect 4940 47840 4956 47904
rect 5020 47840 5036 47904
rect 5100 47840 5116 47904
rect 5180 47840 5188 47904
rect 4868 46816 5188 47840
rect 4868 46752 4876 46816
rect 4940 46752 4956 46816
rect 5020 46752 5036 46816
rect 5100 46752 5116 46816
rect 5180 46752 5188 46816
rect 4868 45728 5188 46752
rect 4868 45664 4876 45728
rect 4940 45664 4956 45728
rect 5020 45664 5036 45728
rect 5100 45664 5116 45728
rect 5180 45664 5188 45728
rect 4868 44640 5188 45664
rect 4868 44576 4876 44640
rect 4940 44576 4956 44640
rect 5020 44576 5036 44640
rect 5100 44576 5116 44640
rect 5180 44576 5188 44640
rect 4868 43552 5188 44576
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 107020 63616 107028 63680
rect 107092 63616 107108 63680
rect 107172 63616 107188 63680
rect 107252 63616 107268 63680
rect 107332 63616 107340 63680
rect 107020 62592 107340 63616
rect 107020 62528 107028 62592
rect 107092 62528 107108 62592
rect 107172 62528 107188 62592
rect 107252 62528 107268 62592
rect 107332 62528 107340 62592
rect 107020 61504 107340 62528
rect 107020 61440 107028 61504
rect 107092 61440 107108 61504
rect 107172 61440 107188 61504
rect 107252 61440 107268 61504
rect 107332 61440 107340 61504
rect 107020 60416 107340 61440
rect 107020 60352 107028 60416
rect 107092 60352 107108 60416
rect 107172 60352 107188 60416
rect 107252 60352 107268 60416
rect 107332 60352 107340 60416
rect 107020 59328 107340 60352
rect 107020 59264 107028 59328
rect 107092 59264 107108 59328
rect 107172 59264 107188 59328
rect 107252 59264 107268 59328
rect 107332 59264 107340 59328
rect 107020 58240 107340 59264
rect 107020 58176 107028 58240
rect 107092 58176 107108 58240
rect 107172 58176 107188 58240
rect 107252 58176 107268 58240
rect 107332 58176 107340 58240
rect 107020 57152 107340 58176
rect 107020 57088 107028 57152
rect 107092 57088 107108 57152
rect 107172 57088 107188 57152
rect 107252 57088 107268 57152
rect 107332 57088 107340 57152
rect 107020 56064 107340 57088
rect 107020 56000 107028 56064
rect 107092 56000 107108 56064
rect 107172 56000 107188 56064
rect 107252 56000 107268 56064
rect 107332 56000 107340 56064
rect 107020 54976 107340 56000
rect 107020 54912 107028 54976
rect 107092 54912 107108 54976
rect 107172 54912 107188 54976
rect 107252 54912 107268 54976
rect 107332 54912 107340 54976
rect 107020 53888 107340 54912
rect 107020 53824 107028 53888
rect 107092 53824 107108 53888
rect 107172 53824 107188 53888
rect 107252 53824 107268 53888
rect 107332 53824 107340 53888
rect 107020 52800 107340 53824
rect 107020 52736 107028 52800
rect 107092 52736 107108 52800
rect 107172 52736 107188 52800
rect 107252 52736 107268 52800
rect 107332 52736 107340 52800
rect 107020 51712 107340 52736
rect 107020 51648 107028 51712
rect 107092 51648 107108 51712
rect 107172 51648 107188 51712
rect 107252 51648 107268 51712
rect 107332 51648 107340 51712
rect 107020 50624 107340 51648
rect 107020 50560 107028 50624
rect 107092 50560 107108 50624
rect 107172 50560 107188 50624
rect 107252 50560 107268 50624
rect 107332 50560 107340 50624
rect 107020 49536 107340 50560
rect 107020 49472 107028 49536
rect 107092 49472 107108 49536
rect 107172 49472 107188 49536
rect 107252 49472 107268 49536
rect 107332 49472 107340 49536
rect 107020 48448 107340 49472
rect 107020 48384 107028 48448
rect 107092 48384 107108 48448
rect 107172 48384 107188 48448
rect 107252 48384 107268 48448
rect 107332 48384 107340 48448
rect 107020 47360 107340 48384
rect 107020 47296 107028 47360
rect 107092 47296 107108 47360
rect 107172 47296 107188 47360
rect 107252 47296 107268 47360
rect 107332 47296 107340 47360
rect 107020 46272 107340 47296
rect 107020 46208 107028 46272
rect 107092 46208 107108 46272
rect 107172 46208 107188 46272
rect 107252 46208 107268 46272
rect 107332 46208 107340 46272
rect 107020 45184 107340 46208
rect 107020 45120 107028 45184
rect 107092 45120 107108 45184
rect 107172 45120 107188 45184
rect 107252 45120 107268 45184
rect 107332 45120 107340 45184
rect 107020 44096 107340 45120
rect 107020 44032 107028 44096
rect 107092 44032 107108 44096
rect 107172 44032 107188 44096
rect 107252 44032 107268 44096
rect 107332 44032 107340 44096
rect 107020 43008 107340 44032
rect 107020 42944 107028 43008
rect 107092 42944 107108 43008
rect 107172 42944 107188 43008
rect 107252 42944 107268 43008
rect 107332 42944 107340 43008
rect 107020 41920 107340 42944
rect 107020 41856 107028 41920
rect 107092 41856 107108 41920
rect 107172 41856 107188 41920
rect 107252 41856 107268 41920
rect 107332 41856 107340 41920
rect 107020 40832 107340 41856
rect 107020 40768 107028 40832
rect 107092 40768 107108 40832
rect 107172 40768 107188 40832
rect 107252 40768 107268 40832
rect 107332 40768 107340 40832
rect 107020 39744 107340 40768
rect 107020 39680 107028 39744
rect 107092 39680 107108 39744
rect 107172 39680 107188 39744
rect 107252 39680 107268 39744
rect 107332 39680 107340 39744
rect 107020 38656 107340 39680
rect 107020 38592 107028 38656
rect 107092 38592 107108 38656
rect 107172 38592 107188 38656
rect 107252 38592 107268 38656
rect 107332 38592 107340 38656
rect 107020 37568 107340 38592
rect 107020 37504 107028 37568
rect 107092 37504 107108 37568
rect 107172 37504 107188 37568
rect 107252 37504 107268 37568
rect 107332 37504 107340 37568
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 10696 36920 11044 36962
rect 10696 36684 10752 36920
rect 10988 36684 11044 36920
rect 10696 36642 11044 36684
rect 100936 36920 101284 36962
rect 100936 36684 100992 36920
rect 101228 36684 101284 36920
rect 100936 36642 101284 36684
rect 107020 36480 107340 37504
rect 107020 36416 107028 36480
rect 107092 36416 107108 36480
rect 107172 36416 107188 36480
rect 107252 36416 107268 36480
rect 107332 36416 107340 36480
rect 10000 36260 10348 36302
rect 10000 36024 10056 36260
rect 10292 36024 10348 36260
rect 10000 35982 10348 36024
rect 101632 36260 101980 36302
rect 101632 36024 101688 36260
rect 101924 36024 101980 36260
rect 101632 35982 101980 36024
rect 107020 36260 107340 36416
rect 107020 36024 107062 36260
rect 107298 36024 107340 36260
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 107020 35392 107340 36024
rect 107020 35328 107028 35392
rect 107092 35328 107108 35392
rect 107172 35328 107188 35392
rect 107252 35328 107268 35392
rect 107332 35328 107340 35392
rect 107020 34304 107340 35328
rect 107020 34240 107028 34304
rect 107092 34240 107108 34304
rect 107172 34240 107188 34304
rect 107252 34240 107268 34304
rect 107332 34240 107340 34304
rect 107020 33216 107340 34240
rect 107020 33152 107028 33216
rect 107092 33152 107108 33216
rect 107172 33152 107188 33216
rect 107252 33152 107268 33216
rect 107332 33152 107340 33216
rect 107020 32128 107340 33152
rect 107020 32064 107028 32128
rect 107092 32064 107108 32128
rect 107172 32064 107188 32128
rect 107252 32064 107268 32128
rect 107332 32064 107340 32128
rect 107020 31040 107340 32064
rect 107020 30976 107028 31040
rect 107092 30976 107108 31040
rect 107172 30976 107188 31040
rect 107252 30976 107268 31040
rect 107332 30976 107340 31040
rect 107020 29952 107340 30976
rect 107020 29888 107028 29952
rect 107092 29888 107108 29952
rect 107172 29888 107188 29952
rect 107252 29888 107268 29952
rect 107332 29888 107340 29952
rect 107020 28864 107340 29888
rect 107020 28800 107028 28864
rect 107092 28800 107108 28864
rect 107172 28800 107188 28864
rect 107252 28800 107268 28864
rect 107332 28800 107340 28864
rect 107020 27776 107340 28800
rect 107020 27712 107028 27776
rect 107092 27712 107108 27776
rect 107172 27712 107188 27776
rect 107252 27712 107268 27776
rect 107332 27712 107340 27776
rect 107020 26688 107340 27712
rect 107020 26624 107028 26688
rect 107092 26624 107108 26688
rect 107172 26624 107188 26688
rect 107252 26624 107268 26688
rect 107332 26624 107340 26688
rect 107020 25600 107340 26624
rect 107020 25536 107028 25600
rect 107092 25536 107108 25600
rect 107172 25536 107188 25600
rect 107252 25536 107268 25600
rect 107332 25536 107340 25600
rect 107020 24512 107340 25536
rect 107020 24448 107028 24512
rect 107092 24448 107108 24512
rect 107172 24448 107188 24512
rect 107252 24448 107268 24512
rect 107332 24448 107340 24512
rect 107020 23424 107340 24448
rect 107020 23360 107028 23424
rect 107092 23360 107108 23424
rect 107172 23360 107188 23424
rect 107252 23360 107268 23424
rect 107332 23360 107340 23424
rect 107020 22336 107340 23360
rect 107020 22272 107028 22336
rect 107092 22272 107108 22336
rect 107172 22272 107188 22336
rect 107252 22272 107268 22336
rect 107332 22272 107340 22336
rect 107020 21248 107340 22272
rect 107020 21184 107028 21248
rect 107092 21184 107108 21248
rect 107172 21184 107188 21248
rect 107252 21184 107268 21248
rect 107332 21184 107340 21248
rect 107020 20160 107340 21184
rect 107020 20096 107028 20160
rect 107092 20096 107108 20160
rect 107172 20096 107188 20160
rect 107252 20096 107268 20160
rect 107332 20096 107340 20160
rect 107020 19072 107340 20096
rect 107020 19008 107028 19072
rect 107092 19008 107108 19072
rect 107172 19008 107188 19072
rect 107252 19008 107268 19072
rect 107332 19008 107340 19072
rect 107020 17984 107340 19008
rect 107020 17920 107028 17984
rect 107092 17920 107108 17984
rect 107172 17920 107188 17984
rect 107252 17920 107268 17984
rect 107332 17920 107340 17984
rect 107020 16896 107340 17920
rect 107020 16832 107028 16896
rect 107092 16832 107108 16896
rect 107172 16832 107188 16896
rect 107252 16832 107268 16896
rect 107332 16832 107340 16896
rect 107020 15808 107340 16832
rect 107020 15744 107028 15808
rect 107092 15744 107108 15808
rect 107172 15744 107188 15808
rect 107252 15744 107268 15808
rect 107332 15744 107340 15808
rect 107020 14720 107340 15744
rect 107020 14656 107028 14720
rect 107092 14656 107108 14720
rect 107172 14656 107188 14720
rect 107252 14656 107268 14720
rect 107332 14656 107340 14720
rect 107020 13632 107340 14656
rect 107020 13568 107028 13632
rect 107092 13568 107108 13632
rect 107172 13568 107188 13632
rect 107252 13568 107268 13632
rect 107332 13568 107340 13632
rect 107020 12544 107340 13568
rect 107020 12480 107028 12544
rect 107092 12480 107108 12544
rect 107172 12480 107188 12544
rect 107252 12480 107268 12544
rect 107332 12480 107340 12544
rect 107020 11456 107340 12480
rect 107020 11392 107028 11456
rect 107092 11392 107108 11456
rect 107172 11392 107188 11456
rect 107252 11392 107268 11456
rect 107332 11392 107340 11456
rect 107020 10368 107340 11392
rect 107020 10304 107028 10368
rect 107092 10304 107108 10368
rect 107172 10304 107188 10368
rect 107252 10304 107268 10368
rect 107332 10304 107340 10368
rect 16060 9893 16120 10038
rect 16057 9892 16123 9893
rect 16057 9828 16058 9892
rect 16122 9828 16123 9892
rect 16057 9827 16123 9828
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 23440 9621 23500 10038
rect 24626 9890 24686 10038
rect 25776 9890 25836 10038
rect 24626 9830 24778 9890
rect 25776 9830 25882 9890
rect 23437 9620 23503 9621
rect 23437 9556 23438 9620
rect 23502 9556 23503 9620
rect 23437 9555 23503 9556
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 24718 7581 24778 9830
rect 25822 8125 25882 9830
rect 25819 8124 25885 8125
rect 25819 8060 25820 8124
rect 25884 8060 25885 8124
rect 25819 8059 25885 8060
rect 26926 7581 26986 10038
rect 28122 9890 28182 10038
rect 29280 9890 29340 10038
rect 28122 9830 28274 9890
rect 29280 9830 29378 9890
rect 28214 7581 28274 9830
rect 29318 8125 29378 9830
rect 30448 9621 30508 10038
rect 31616 9757 31676 10038
rect 32784 9890 32844 10038
rect 33952 9890 34012 10038
rect 32784 9830 32874 9890
rect 31613 9756 31679 9757
rect 31613 9692 31614 9756
rect 31678 9692 31679 9756
rect 31613 9691 31679 9692
rect 30445 9620 30511 9621
rect 30445 9556 30446 9620
rect 30510 9556 30511 9620
rect 30445 9555 30511 9556
rect 32814 8125 32874 9830
rect 33918 9830 34012 9890
rect 35120 9890 35180 10038
rect 36288 9890 36348 10038
rect 37456 9890 37516 10038
rect 35120 9830 35266 9890
rect 36288 9830 36370 9890
rect 29315 8124 29381 8125
rect 29315 8060 29316 8124
rect 29380 8060 29381 8124
rect 29315 8059 29381 8060
rect 32811 8124 32877 8125
rect 32811 8060 32812 8124
rect 32876 8060 32877 8124
rect 32811 8059 32877 8060
rect 33918 7581 33978 9830
rect 35206 8125 35266 9830
rect 35203 8124 35269 8125
rect 35203 8060 35204 8124
rect 35268 8060 35269 8124
rect 35203 8059 35269 8060
rect 24715 7580 24781 7581
rect 24715 7516 24716 7580
rect 24780 7516 24781 7580
rect 24715 7515 24781 7516
rect 26923 7580 26989 7581
rect 26923 7516 26924 7580
rect 26988 7516 26989 7580
rect 26923 7515 26989 7516
rect 28211 7580 28277 7581
rect 28211 7516 28212 7580
rect 28276 7516 28277 7580
rect 28211 7515 28277 7516
rect 33915 7580 33981 7581
rect 33915 7516 33916 7580
rect 33980 7516 33981 7580
rect 33915 7515 33981 7516
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 7104 35248 7880
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 7648 35908 8064
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 36310 7581 36370 9830
rect 37414 9830 37516 9890
rect 38624 9890 38684 10038
rect 38624 9830 38762 9890
rect 37414 7581 37474 9830
rect 38702 8125 38762 9830
rect 38699 8124 38765 8125
rect 38699 8060 38700 8124
rect 38764 8060 38765 8124
rect 38699 8059 38765 8060
rect 39806 7581 39866 10038
rect 40960 9890 41020 10038
rect 40910 9830 41020 9890
rect 42128 9890 42188 10038
rect 42128 9830 42258 9890
rect 40910 7581 40970 9830
rect 42198 7581 42258 9830
rect 43302 7581 43362 10038
rect 90403 9892 90469 9893
rect 90403 9828 90404 9892
rect 90468 9890 90469 9892
rect 90529 9890 90589 10038
rect 90468 9830 90589 9890
rect 90468 9828 90469 9830
rect 90403 9827 90469 9828
rect 36307 7580 36373 7581
rect 36307 7516 36308 7580
rect 36372 7516 36373 7580
rect 36307 7515 36373 7516
rect 37411 7580 37477 7581
rect 37411 7516 37412 7580
rect 37476 7516 37477 7580
rect 37411 7515 37477 7516
rect 39803 7580 39869 7581
rect 39803 7516 39804 7580
rect 39868 7516 39869 7580
rect 39803 7515 39869 7516
rect 40907 7580 40973 7581
rect 40907 7516 40908 7580
rect 40972 7516 40973 7580
rect 40907 7515 40973 7516
rect 42195 7580 42261 7581
rect 42195 7516 42196 7580
rect 42260 7516 42261 7580
rect 42195 7515 42261 7516
rect 43299 7580 43365 7581
rect 43299 7516 43300 7580
rect 43364 7516 43365 7580
rect 43299 7515 43365 7516
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
rect 65648 7104 65968 8064
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5624 65968 5952
rect 65648 5388 65690 5624
rect 65926 5388 65968 5624
rect 65648 4928 65968 5388
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 66308 7648 66628 8064
rect 66308 7584 66316 7648
rect 66380 7584 66396 7648
rect 66460 7584 66476 7648
rect 66540 7584 66556 7648
rect 66620 7584 66628 7648
rect 66308 6560 66628 7584
rect 90406 7581 90466 9827
rect 90682 9485 90742 10038
rect 90816 9890 90876 10038
rect 90955 9892 91021 9893
rect 90955 9890 90956 9892
rect 90816 9830 90956 9890
rect 90955 9828 90956 9830
rect 91020 9828 91021 9892
rect 90955 9827 91021 9828
rect 90679 9484 90745 9485
rect 90679 9420 90680 9484
rect 90744 9420 90745 9484
rect 90679 9419 90745 9420
rect 90958 7581 91018 9827
rect 107020 9280 107340 10304
rect 107020 9216 107028 9280
rect 107092 9216 107108 9280
rect 107172 9216 107188 9280
rect 107252 9216 107268 9280
rect 107332 9216 107340 9280
rect 107020 8192 107340 9216
rect 107020 8128 107028 8192
rect 107092 8128 107108 8192
rect 107172 8128 107188 8192
rect 107252 8128 107268 8192
rect 107332 8128 107340 8192
rect 90403 7580 90469 7581
rect 90403 7516 90404 7580
rect 90468 7516 90469 7580
rect 90403 7515 90469 7516
rect 90955 7580 91021 7581
rect 90955 7516 90956 7580
rect 91020 7516 91021 7580
rect 90955 7515 91021 7516
rect 66308 6496 66316 6560
rect 66380 6496 66396 6560
rect 66460 6496 66476 6560
rect 66540 6496 66556 6560
rect 66620 6496 66628 6560
rect 66308 6284 66628 6496
rect 66308 6048 66350 6284
rect 66586 6048 66628 6284
rect 66308 5472 66628 6048
rect 66308 5408 66316 5472
rect 66380 5408 66396 5472
rect 66460 5408 66476 5472
rect 66540 5408 66556 5472
rect 66620 5408 66628 5472
rect 66308 4384 66628 5408
rect 66308 4320 66316 4384
rect 66380 4320 66396 4384
rect 66460 4320 66476 4384
rect 66540 4320 66556 4384
rect 66620 4320 66628 4384
rect 66308 3296 66628 4320
rect 66308 3232 66316 3296
rect 66380 3232 66396 3296
rect 66460 3232 66476 3296
rect 66540 3232 66556 3296
rect 66620 3232 66628 3296
rect 66308 2208 66628 3232
rect 66308 2144 66316 2208
rect 66380 2144 66396 2208
rect 66460 2144 66476 2208
rect 66540 2144 66556 2208
rect 66620 2144 66628 2208
rect 66308 2128 66628 2144
rect 96368 7104 96688 8064
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 5624 96688 5952
rect 96368 5388 96410 5624
rect 96646 5388 96688 5624
rect 96368 4928 96688 5388
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2128 96688 2688
rect 97028 7648 97348 8064
rect 97028 7584 97036 7648
rect 97100 7584 97116 7648
rect 97180 7584 97196 7648
rect 97260 7584 97276 7648
rect 97340 7584 97348 7648
rect 97028 6560 97348 7584
rect 107020 7104 107340 8128
rect 107020 7040 107028 7104
rect 107092 7040 107108 7104
rect 107172 7040 107188 7104
rect 107252 7040 107268 7104
rect 107332 7040 107340 7104
rect 107020 7024 107340 7040
rect 107756 66400 108076 66416
rect 107756 66336 107764 66400
rect 107828 66336 107844 66400
rect 107908 66336 107924 66400
rect 107988 66336 108004 66400
rect 108068 66336 108076 66400
rect 107756 65312 108076 66336
rect 107756 65248 107764 65312
rect 107828 65248 107844 65312
rect 107908 65248 107924 65312
rect 107988 65248 108004 65312
rect 108068 65248 108076 65312
rect 107756 64224 108076 65248
rect 107756 64160 107764 64224
rect 107828 64160 107844 64224
rect 107908 64160 107924 64224
rect 107988 64160 108004 64224
rect 108068 64160 108076 64224
rect 107756 63136 108076 64160
rect 107756 63072 107764 63136
rect 107828 63072 107844 63136
rect 107908 63072 107924 63136
rect 107988 63072 108004 63136
rect 108068 63072 108076 63136
rect 107756 62048 108076 63072
rect 107756 61984 107764 62048
rect 107828 61984 107844 62048
rect 107908 61984 107924 62048
rect 107988 61984 108004 62048
rect 108068 61984 108076 62048
rect 107756 60960 108076 61984
rect 107756 60896 107764 60960
rect 107828 60896 107844 60960
rect 107908 60896 107924 60960
rect 107988 60896 108004 60960
rect 108068 60896 108076 60960
rect 107756 59872 108076 60896
rect 107756 59808 107764 59872
rect 107828 59808 107844 59872
rect 107908 59808 107924 59872
rect 107988 59808 108004 59872
rect 108068 59808 108076 59872
rect 107756 58784 108076 59808
rect 107756 58720 107764 58784
rect 107828 58720 107844 58784
rect 107908 58720 107924 58784
rect 107988 58720 108004 58784
rect 108068 58720 108076 58784
rect 107756 57696 108076 58720
rect 107756 57632 107764 57696
rect 107828 57632 107844 57696
rect 107908 57632 107924 57696
rect 107988 57632 108004 57696
rect 108068 57632 108076 57696
rect 107756 56608 108076 57632
rect 107756 56544 107764 56608
rect 107828 56544 107844 56608
rect 107908 56544 107924 56608
rect 107988 56544 108004 56608
rect 108068 56544 108076 56608
rect 107756 55520 108076 56544
rect 107756 55456 107764 55520
rect 107828 55456 107844 55520
rect 107908 55456 107924 55520
rect 107988 55456 108004 55520
rect 108068 55456 108076 55520
rect 107756 54432 108076 55456
rect 107756 54368 107764 54432
rect 107828 54368 107844 54432
rect 107908 54368 107924 54432
rect 107988 54368 108004 54432
rect 108068 54368 108076 54432
rect 107756 53344 108076 54368
rect 107756 53280 107764 53344
rect 107828 53280 107844 53344
rect 107908 53280 107924 53344
rect 107988 53280 108004 53344
rect 108068 53280 108076 53344
rect 107756 52256 108076 53280
rect 107756 52192 107764 52256
rect 107828 52192 107844 52256
rect 107908 52192 107924 52256
rect 107988 52192 108004 52256
rect 108068 52192 108076 52256
rect 107756 51168 108076 52192
rect 107756 51104 107764 51168
rect 107828 51104 107844 51168
rect 107908 51104 107924 51168
rect 107988 51104 108004 51168
rect 108068 51104 108076 51168
rect 107756 50080 108076 51104
rect 107756 50016 107764 50080
rect 107828 50016 107844 50080
rect 107908 50016 107924 50080
rect 107988 50016 108004 50080
rect 108068 50016 108076 50080
rect 107756 48992 108076 50016
rect 107756 48928 107764 48992
rect 107828 48928 107844 48992
rect 107908 48928 107924 48992
rect 107988 48928 108004 48992
rect 108068 48928 108076 48992
rect 107756 47904 108076 48928
rect 107756 47840 107764 47904
rect 107828 47840 107844 47904
rect 107908 47840 107924 47904
rect 107988 47840 108004 47904
rect 108068 47840 108076 47904
rect 107756 46816 108076 47840
rect 107756 46752 107764 46816
rect 107828 46752 107844 46816
rect 107908 46752 107924 46816
rect 107988 46752 108004 46816
rect 108068 46752 108076 46816
rect 107756 45728 108076 46752
rect 107756 45664 107764 45728
rect 107828 45664 107844 45728
rect 107908 45664 107924 45728
rect 107988 45664 108004 45728
rect 108068 45664 108076 45728
rect 107756 44640 108076 45664
rect 107756 44576 107764 44640
rect 107828 44576 107844 44640
rect 107908 44576 107924 44640
rect 107988 44576 108004 44640
rect 108068 44576 108076 44640
rect 107756 43552 108076 44576
rect 107756 43488 107764 43552
rect 107828 43488 107844 43552
rect 107908 43488 107924 43552
rect 107988 43488 108004 43552
rect 108068 43488 108076 43552
rect 107756 42464 108076 43488
rect 107756 42400 107764 42464
rect 107828 42400 107844 42464
rect 107908 42400 107924 42464
rect 107988 42400 108004 42464
rect 108068 42400 108076 42464
rect 107756 41376 108076 42400
rect 107756 41312 107764 41376
rect 107828 41312 107844 41376
rect 107908 41312 107924 41376
rect 107988 41312 108004 41376
rect 108068 41312 108076 41376
rect 107756 40288 108076 41312
rect 107756 40224 107764 40288
rect 107828 40224 107844 40288
rect 107908 40224 107924 40288
rect 107988 40224 108004 40288
rect 108068 40224 108076 40288
rect 107756 39200 108076 40224
rect 107756 39136 107764 39200
rect 107828 39136 107844 39200
rect 107908 39136 107924 39200
rect 107988 39136 108004 39200
rect 108068 39136 108076 39200
rect 107756 38112 108076 39136
rect 107756 38048 107764 38112
rect 107828 38048 107844 38112
rect 107908 38048 107924 38112
rect 107988 38048 108004 38112
rect 108068 38048 108076 38112
rect 107756 37024 108076 38048
rect 107756 36960 107764 37024
rect 107828 36960 107844 37024
rect 107908 36960 107924 37024
rect 107988 36960 108004 37024
rect 108068 36960 108076 37024
rect 107756 36920 108076 36960
rect 107756 36684 107798 36920
rect 108034 36684 108076 36920
rect 107756 35936 108076 36684
rect 107756 35872 107764 35936
rect 107828 35872 107844 35936
rect 107908 35872 107924 35936
rect 107988 35872 108004 35936
rect 108068 35872 108076 35936
rect 107756 34848 108076 35872
rect 107756 34784 107764 34848
rect 107828 34784 107844 34848
rect 107908 34784 107924 34848
rect 107988 34784 108004 34848
rect 108068 34784 108076 34848
rect 107756 33760 108076 34784
rect 107756 33696 107764 33760
rect 107828 33696 107844 33760
rect 107908 33696 107924 33760
rect 107988 33696 108004 33760
rect 108068 33696 108076 33760
rect 107756 32672 108076 33696
rect 107756 32608 107764 32672
rect 107828 32608 107844 32672
rect 107908 32608 107924 32672
rect 107988 32608 108004 32672
rect 108068 32608 108076 32672
rect 107756 31584 108076 32608
rect 107756 31520 107764 31584
rect 107828 31520 107844 31584
rect 107908 31520 107924 31584
rect 107988 31520 108004 31584
rect 108068 31520 108076 31584
rect 107756 30496 108076 31520
rect 107756 30432 107764 30496
rect 107828 30432 107844 30496
rect 107908 30432 107924 30496
rect 107988 30432 108004 30496
rect 108068 30432 108076 30496
rect 107756 29408 108076 30432
rect 107756 29344 107764 29408
rect 107828 29344 107844 29408
rect 107908 29344 107924 29408
rect 107988 29344 108004 29408
rect 108068 29344 108076 29408
rect 107756 28320 108076 29344
rect 107756 28256 107764 28320
rect 107828 28256 107844 28320
rect 107908 28256 107924 28320
rect 107988 28256 108004 28320
rect 108068 28256 108076 28320
rect 107756 27232 108076 28256
rect 107756 27168 107764 27232
rect 107828 27168 107844 27232
rect 107908 27168 107924 27232
rect 107988 27168 108004 27232
rect 108068 27168 108076 27232
rect 107756 26144 108076 27168
rect 107756 26080 107764 26144
rect 107828 26080 107844 26144
rect 107908 26080 107924 26144
rect 107988 26080 108004 26144
rect 108068 26080 108076 26144
rect 107756 25056 108076 26080
rect 107756 24992 107764 25056
rect 107828 24992 107844 25056
rect 107908 24992 107924 25056
rect 107988 24992 108004 25056
rect 108068 24992 108076 25056
rect 107756 23968 108076 24992
rect 107756 23904 107764 23968
rect 107828 23904 107844 23968
rect 107908 23904 107924 23968
rect 107988 23904 108004 23968
rect 108068 23904 108076 23968
rect 107756 22880 108076 23904
rect 107756 22816 107764 22880
rect 107828 22816 107844 22880
rect 107908 22816 107924 22880
rect 107988 22816 108004 22880
rect 108068 22816 108076 22880
rect 107756 21792 108076 22816
rect 107756 21728 107764 21792
rect 107828 21728 107844 21792
rect 107908 21728 107924 21792
rect 107988 21728 108004 21792
rect 108068 21728 108076 21792
rect 107756 20704 108076 21728
rect 107756 20640 107764 20704
rect 107828 20640 107844 20704
rect 107908 20640 107924 20704
rect 107988 20640 108004 20704
rect 108068 20640 108076 20704
rect 107756 19616 108076 20640
rect 107756 19552 107764 19616
rect 107828 19552 107844 19616
rect 107908 19552 107924 19616
rect 107988 19552 108004 19616
rect 108068 19552 108076 19616
rect 107756 18528 108076 19552
rect 107756 18464 107764 18528
rect 107828 18464 107844 18528
rect 107908 18464 107924 18528
rect 107988 18464 108004 18528
rect 108068 18464 108076 18528
rect 107756 17440 108076 18464
rect 107756 17376 107764 17440
rect 107828 17376 107844 17440
rect 107908 17376 107924 17440
rect 107988 17376 108004 17440
rect 108068 17376 108076 17440
rect 107756 16352 108076 17376
rect 107756 16288 107764 16352
rect 107828 16288 107844 16352
rect 107908 16288 107924 16352
rect 107988 16288 108004 16352
rect 108068 16288 108076 16352
rect 107756 15264 108076 16288
rect 107756 15200 107764 15264
rect 107828 15200 107844 15264
rect 107908 15200 107924 15264
rect 107988 15200 108004 15264
rect 108068 15200 108076 15264
rect 107756 14176 108076 15200
rect 107756 14112 107764 14176
rect 107828 14112 107844 14176
rect 107908 14112 107924 14176
rect 107988 14112 108004 14176
rect 108068 14112 108076 14176
rect 107756 13088 108076 14112
rect 107756 13024 107764 13088
rect 107828 13024 107844 13088
rect 107908 13024 107924 13088
rect 107988 13024 108004 13088
rect 108068 13024 108076 13088
rect 107756 12000 108076 13024
rect 107756 11936 107764 12000
rect 107828 11936 107844 12000
rect 107908 11936 107924 12000
rect 107988 11936 108004 12000
rect 108068 11936 108076 12000
rect 107756 10912 108076 11936
rect 107756 10848 107764 10912
rect 107828 10848 107844 10912
rect 107908 10848 107924 10912
rect 107988 10848 108004 10912
rect 108068 10848 108076 10912
rect 107756 9824 108076 10848
rect 107756 9760 107764 9824
rect 107828 9760 107844 9824
rect 107908 9760 107924 9824
rect 107988 9760 108004 9824
rect 108068 9760 108076 9824
rect 107756 8736 108076 9760
rect 107756 8672 107764 8736
rect 107828 8672 107844 8736
rect 107908 8672 107924 8736
rect 107988 8672 108004 8736
rect 108068 8672 108076 8736
rect 107756 7648 108076 8672
rect 107756 7584 107764 7648
rect 107828 7584 107844 7648
rect 107908 7584 107924 7648
rect 107988 7584 108004 7648
rect 108068 7584 108076 7648
rect 107756 7024 108076 7584
rect 97028 6496 97036 6560
rect 97100 6496 97116 6560
rect 97180 6496 97196 6560
rect 97260 6496 97276 6560
rect 97340 6496 97348 6560
rect 97028 6284 97348 6496
rect 97028 6048 97070 6284
rect 97306 6048 97348 6284
rect 97028 5472 97348 6048
rect 97028 5408 97036 5472
rect 97100 5408 97116 5472
rect 97180 5408 97196 5472
rect 97260 5408 97276 5472
rect 97340 5408 97348 5472
rect 97028 4384 97348 5408
rect 97028 4320 97036 4384
rect 97100 4320 97116 4384
rect 97180 4320 97196 4384
rect 97260 4320 97276 4384
rect 97340 4320 97348 4384
rect 97028 3296 97348 4320
rect 97028 3232 97036 3296
rect 97100 3232 97116 3296
rect 97180 3232 97196 3296
rect 97260 3232 97276 3296
rect 97340 3232 97348 3296
rect 97028 2208 97348 3232
rect 97028 2144 97036 2208
rect 97100 2144 97116 2208
rect 97180 2144 97196 2208
rect 97260 2144 97276 2208
rect 97340 2144 97348 2208
rect 97028 2128 97348 2144
<< via4 >>
rect 4250 66880 4280 66896
rect 4280 66880 4296 66896
rect 4296 66880 4360 66896
rect 4360 66880 4376 66896
rect 4376 66880 4440 66896
rect 4440 66880 4456 66896
rect 4456 66880 4486 66896
rect 4250 66660 4486 66880
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 67488 5146 67556
rect 4910 67424 4940 67488
rect 4940 67424 4956 67488
rect 4956 67424 5020 67488
rect 5020 67424 5036 67488
rect 5036 67424 5100 67488
rect 5100 67424 5116 67488
rect 5116 67424 5146 67488
rect 4910 67320 5146 67424
rect 34970 66880 35000 66896
rect 35000 66880 35016 66896
rect 35016 66880 35080 66896
rect 35080 66880 35096 66896
rect 35096 66880 35160 66896
rect 35160 66880 35176 66896
rect 35176 66880 35206 66896
rect 34970 66660 35206 66880
rect 35630 67488 35866 67556
rect 35630 67424 35660 67488
rect 35660 67424 35676 67488
rect 35676 67424 35740 67488
rect 35740 67424 35756 67488
rect 35756 67424 35820 67488
rect 35820 67424 35836 67488
rect 35836 67424 35866 67488
rect 35630 67320 35866 67424
rect 65690 66880 65720 66896
rect 65720 66880 65736 66896
rect 65736 66880 65800 66896
rect 65800 66880 65816 66896
rect 65816 66880 65880 66896
rect 65880 66880 65896 66896
rect 65896 66880 65926 66896
rect 65690 66660 65926 66880
rect 66350 67488 66586 67556
rect 66350 67424 66380 67488
rect 66380 67424 66396 67488
rect 66396 67424 66460 67488
rect 66460 67424 66476 67488
rect 66476 67424 66540 67488
rect 66540 67424 66556 67488
rect 66556 67424 66586 67488
rect 66350 67320 66586 67424
rect 96410 66880 96440 66896
rect 96440 66880 96456 66896
rect 96456 66880 96520 66896
rect 96520 66880 96536 66896
rect 96536 66880 96600 66896
rect 96600 66880 96616 66896
rect 96616 66880 96646 66896
rect 96410 66660 96646 66880
rect 97070 67488 97306 67556
rect 97070 67424 97100 67488
rect 97100 67424 97116 67488
rect 97116 67424 97180 67488
rect 97180 67424 97196 67488
rect 97196 67424 97260 67488
rect 97260 67424 97276 67488
rect 97276 67424 97306 67488
rect 97070 67320 97306 67424
rect 4910 36684 5146 36920
rect 10752 36684 10988 36920
rect 100992 36684 101228 36920
rect 10056 36024 10292 36260
rect 101688 36024 101924 36260
rect 107062 36024 107298 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 6048 35866 6284
rect 65690 5388 65926 5624
rect 66350 6048 66586 6284
rect 96410 5388 96646 5624
rect 107798 36684 108034 36920
rect 97070 6048 97306 6284
<< metal5 >>
rect 1056 67556 110908 67598
rect 1056 67320 4910 67556
rect 5146 67320 35630 67556
rect 35866 67320 66350 67556
rect 66586 67320 97070 67556
rect 97306 67320 110908 67556
rect 1056 67278 110908 67320
rect 1056 66896 110908 66938
rect 1056 66660 4250 66896
rect 4486 66660 34970 66896
rect 35206 66660 65690 66896
rect 65926 66660 96410 66896
rect 96646 66660 110908 66896
rect 1056 66618 110908 66660
rect 1056 36920 110908 36962
rect 1056 36684 4910 36920
rect 5146 36684 10752 36920
rect 10988 36684 100992 36920
rect 101228 36684 107798 36920
rect 108034 36684 110908 36920
rect 1056 36642 110908 36684
rect 1056 36260 110908 36302
rect 1056 36024 4250 36260
rect 4486 36024 10056 36260
rect 10292 36024 101688 36260
rect 101924 36024 107062 36260
rect 107298 36024 110908 36260
rect 1056 35982 110908 36024
rect 1056 6284 110908 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 66350 6284
rect 66586 6048 97070 6284
rect 97306 6048 110908 6284
rect 1056 6006 110908 6048
rect 1056 5624 110908 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 65690 5624
rect 65926 5388 96410 5624
rect 96646 5388 110908 5624
rect 1056 5346 110908 5388
use sky130_fd_sc_hd__inv_2  _040_
timestamp 1
transform -1 0 104604 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _041_
timestamp 1
transform -1 0 59156 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _042_
timestamp 1
transform -1 0 104972 0 1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _043_
timestamp 1
transform 1 0 104328 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _044_
timestamp 1
transform 1 0 104328 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _045_
timestamp 1
transform 1 0 104328 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _046_
timestamp 1
transform -1 0 105708 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _047_
timestamp 1
transform 1 0 105432 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _048_
timestamp 1
transform 1 0 104788 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _049_
timestamp 1
transform 1 0 104788 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _050_
timestamp 1
transform 1 0 104328 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _051_
timestamp 1
transform 1 0 104420 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _052_
timestamp 1
transform 1 0 104328 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _053_
timestamp 1
transform 1 0 104328 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _054_
timestamp 1
transform 1 0 104788 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _055_
timestamp 1
transform -1 0 104972 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 1
transform -1 0 60996 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1
transform -1 0 63296 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1
transform 1 0 64768 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 1
transform -1 0 66424 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1
transform -1 0 68080 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1
transform -1 0 69736 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1
transform -1 0 71576 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1
transform -1 0 73600 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1
transform 1 0 75900 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1
transform 1 0 91908 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _066_
timestamp 1
transform 1 0 104328 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _067_
timestamp 1
transform 1 0 104328 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1
transform 1 0 104328 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp 1
transform 1 0 104328 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1
transform 1 0 104328 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp 1
transform 1 0 104328 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp 1
transform 1 0 104788 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1
transform -1 0 48852 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1
transform -1 0 50692 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1
transform -1 0 52624 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 1
transform -1 0 54188 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1
transform -1 0 55844 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1
transform -1 0 58144 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _079_
timestamp 1
transform 1 0 55384 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _080_
timestamp 1
transform 1 0 57868 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _081_
timestamp 1
transform 1 0 59708 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _082_
timestamp 1
transform 1 0 61364 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _083_
timestamp 1
transform 1 0 63664 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _084_
timestamp 1
transform 1 0 65596 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _085_
timestamp 1
transform 1 0 68172 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _086_
timestamp 1
transform 1 0 70012 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _087_
timestamp 1
transform 1 0 71760 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _088_
timestamp 1
transform 1 0 74336 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _089_
timestamp 1
transform 1 0 104328 0 -1 57664
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _090_
timestamp 1
transform 1 0 104328 0 1 54400
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _091_
timestamp 1
transform 1 0 104328 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _092_
timestamp 1
transform -1 0 106168 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _093_
timestamp 1
transform -1 0 106168 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _094_
timestamp 1
transform 1 0 104328 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _095_
timestamp 1
transform 1 0 104328 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _096_
timestamp 1
transform 1 0 104328 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _097_
timestamp 1
transform 1 0 43332 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _098_
timestamp 1
transform 1 0 45540 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _099_
timestamp 1
transform 1 0 47748 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _100_
timestamp 1
transform 1 0 49680 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _101_
timestamp 1
transform 1 0 51612 0 1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _102_
timestamp 1
transform 1 0 53544 0 -1 67456
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform -1 0 43332 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform -1 0 45540 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform -1 0 47748 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 51704 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__042__A
timestamp 1
transform 1 0 104972 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__042__B
timestamp 1
transform 1 0 105156 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__043__A
timestamp 1
transform 1 0 105064 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__043__B
timestamp 1
transform -1 0 105432 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__043__C
timestamp 1
transform 1 0 105432 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__043__X
timestamp 1
transform -1 0 105064 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__044__A1
timestamp 1
transform 1 0 104696 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__044__A2
timestamp 1
transform 1 0 104880 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__044__B1
timestamp 1
transform -1 0 105248 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__045__A
timestamp 1
transform 1 0 104604 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__046__B
timestamp 1
transform 1 0 105708 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__047__B
timestamp 1
transform -1 0 106260 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__048__C
timestamp 1
transform 1 0 104604 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__050__C
timestamp 1
transform 1 0 105248 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__051__A1_N
timestamp 1
transform 1 0 105156 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__051__B2
timestamp 1
transform 1 0 105340 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__052__A
timestamp 1
transform 1 0 105248 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__052__B
timestamp 1
transform 1 0 105064 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__053__A1
timestamp 1
transform 1 0 104696 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__053__B1
timestamp 1
transform 1 0 104880 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1
transform 1 0 92368 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__Y
timestamp 1
transform 1 0 92184 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1
transform 1 0 104604 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1
transform 1 0 104604 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1
transform 1 0 104604 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1
transform 1 0 104604 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1
transform 1 0 104604 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1
transform 1 0 104604 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1
transform 1 0 105064 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__CLK
timestamp 1
transform 1 0 57224 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__CLK
timestamp 1
transform 1 0 57592 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__CLK
timestamp 1
transform 1 0 59524 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__CLK
timestamp 1
transform 1 0 61180 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__CLK
timestamp 1
transform 1 0 63480 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__CLK
timestamp 1
transform 1 0 65596 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__CLK
timestamp 1
transform 1 0 67896 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__CLK
timestamp 1
transform 1 0 69828 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__CLK
timestamp 1
transform 1 0 73600 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__CLK
timestamp 1
transform 1 0 76176 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__CLK
timestamp 1
transform 1 0 106628 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__Q
timestamp 1
transform -1 0 106628 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__RESET_B
timestamp 1
transform 1 0 104328 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__CLK
timestamp 1
transform -1 0 106904 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__Q
timestamp 1
transform -1 0 106628 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__CLK
timestamp 1
transform 1 0 106352 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__Q
timestamp 1
transform -1 0 106352 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__CLK
timestamp 1
transform 1 0 106168 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__CLK
timestamp 1
transform 1 0 106168 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__CLK
timestamp 1
transform 1 0 106444 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__Q
timestamp 1
transform -1 0 106444 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__CLK
timestamp 1
transform 1 0 106352 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__Q
timestamp 1
transform -1 0 106352 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__CLK
timestamp 1
transform 1 0 106352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__Q
timestamp 1
transform -1 0 106352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__CLK
timestamp 1
transform 1 0 45172 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__CLK
timestamp 1
transform 1 0 47564 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__CLK
timestamp 1
transform 1 0 49588 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__CLK
timestamp 1
transform 1 0 51704 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__CLK
timestamp 1
transform 1 0 53452 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__CLK
timestamp 1
transform 1 0 55384 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1
transform 1 0 63480 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 1
transform 1 0 63296 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 1
transform 1 0 58144 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_X
timestamp 1
transform 1 0 58328 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 1
transform -1 0 104972 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_X
timestamp 1
transform 1 0 106168 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 1
transform 1 0 106536 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout18_A
timestamp 1
transform 1 0 65044 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout19_A
timestamp 1
transform 1 0 76176 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout20_X
timestamp 1
transform -1 0 105524 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold1_A
timestamp 1
transform 1 0 105156 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1
transform 1 0 104328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1
transform -1 0 110308 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr0[0]
timestamp 1
transform -1 0 23644 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr0[1]
timestamp 1
transform -1 0 24840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr0[2]
timestamp 1
transform 1 0 7452 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr0[3]
timestamp 1
transform -1 0 7636 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr0[4]
timestamp 1
transform 1 0 7452 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr0[5]
timestamp 1
transform -1 0 7636 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr0[6]
timestamp 1
transform -1 0 7636 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr0[7]
timestamp 1
transform -1 0 7636 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[0]
timestamp 1
transform -1 0 87492 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[1]
timestamp 1
transform -1 0 86388 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[2]
timestamp 1
transform -1 0 104512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[5]
timestamp 1
transform -1 0 90712 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[6]
timestamp 1
transform -1 0 90896 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_addr1[7]
timestamp 1
transform -1 0 91080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_clk0
timestamp 1
transform -1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_clk1
timestamp 1
transform 1 0 95864 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_csb0
timestamp 1
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[0]
timestamp 1
transform -1 0 26036 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[1]
timestamp 1
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[2]
timestamp 1
transform 1 0 28152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[3]
timestamp 1
transform -1 0 29716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[4]
timestamp 1
transform -1 0 30636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[5]
timestamp 1
transform -1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[6]
timestamp 1
transform -1 0 33028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[7]
timestamp 1
transform 1 0 33948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[8]
timestamp 1
transform 1 0 35144 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[9]
timestamp 1
transform -1 0 36524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[10]
timestamp 1
transform -1 0 37628 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[11]
timestamp 1
transform -1 0 38824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[12]
timestamp 1
transform 1 0 39836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[13]
timestamp 1
transform 1 0 41032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[14]
timestamp 1
transform -1 0 42320 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_i_din0[15]
timestamp 1
transform -1 0 43516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 62928 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1
transform -1 0 57776 0 -1 66368
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1
transform 1 0 104328 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp 1
transform 1 0 104328 0 -1 42432
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_4  fanout18
timestamp 1
transform -1 0 64768 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1
transform -1 0 75808 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout20
timestamp 1
transform -1 0 105340 0 -1 32640
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636968456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636968456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636968456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636968456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636968456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636968456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636968456
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636968456
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1636968456
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636968456
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1636968456
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1636968456
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1636968456
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1636968456
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636968456
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636968456
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636968456
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1636968456
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1636968456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1636968456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1636968456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1636968456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1636968456
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1636968456
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_617
timestamp 1636968456
transform 1 0 57868 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_629
timestamp 1636968456
transform 1 0 58972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 1
transform 1 0 60076 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1636968456
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1636968456
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1636968456
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1636968456
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1636968456
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1636968456
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1636968456
transform 1 0 68172 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1636968456
transform 1 0 69276 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1636968456
transform 1 0 70748 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1636968456
transform 1 0 71852 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1
transform 1 0 72956 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1636968456
transform 1 0 73324 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1636968456
transform 1 0 74428 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1
transform 1 0 75532 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_813
timestamp 1636968456
transform 1 0 75900 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_825
timestamp 1636968456
transform 1 0 77004 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_837
timestamp 1
transform 1 0 78108 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_841
timestamp 1636968456
transform 1 0 78476 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_853
timestamp 1636968456
transform 1 0 79580 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_865
timestamp 1
transform 1 0 80684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1636968456
transform 1 0 81052 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1636968456
transform 1 0 82156 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 1
transform 1 0 83260 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1636968456
transform 1 0 83628 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_909
timestamp 1636968456
transform 1 0 84732 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_921
timestamp 1
transform 1 0 85836 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_925
timestamp 1636968456
transform 1 0 86204 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_937
timestamp 1636968456
transform 1 0 87308 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_949
timestamp 1
transform 1 0 88412 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_953
timestamp 1636968456
transform 1 0 88780 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_965
timestamp 1636968456
transform 1 0 89884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_977
timestamp 1
transform 1 0 90988 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_981
timestamp 1636968456
transform 1 0 91356 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_993
timestamp 1636968456
transform 1 0 92460 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1005
timestamp 1
transform 1 0 93564 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1009
timestamp 1636968456
transform 1 0 93932 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1021
timestamp 1636968456
transform 1 0 95036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1033
timestamp 1
transform 1 0 96140 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1037
timestamp 1636968456
transform 1 0 96508 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1049
timestamp 1636968456
transform 1 0 97612 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1061
timestamp 1
transform 1 0 98716 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1065
timestamp 1636968456
transform 1 0 99084 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1077
timestamp 1636968456
transform 1 0 100188 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1089
timestamp 1
transform 1 0 101292 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1093
timestamp 1636968456
transform 1 0 101660 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1105
timestamp 1636968456
transform 1 0 102764 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1121
timestamp 1636968456
transform 1 0 104236 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1133
timestamp 1636968456
transform 1 0 105340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1145
timestamp 1
transform 1 0 106444 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1149
timestamp 1636968456
transform 1 0 106812 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1161
timestamp 1636968456
transform 1 0 107916 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1173
timestamp 1
transform 1 0 109020 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1177
timestamp 1636968456
transform 1 0 109388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1189
timestamp 1
transform 1 0 110492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636968456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636968456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636968456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636968456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636968456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636968456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636968456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636968456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636968456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636968456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636968456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636968456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636968456
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636968456
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636968456
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636968456
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636968456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636968456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636968456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636968456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636968456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636968456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636968456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636968456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636968456
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636968456
transform 1 0 58972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636968456
transform 1 0 60076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636968456
transform 1 0 61180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1
transform 1 0 62284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636968456
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636968456
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636968456
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636968456
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636968456
transform 1 0 68172 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636968456
transform 1 0 69276 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636968456
transform 1 0 70380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636968456
transform 1 0 71484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1
transform 1 0 72588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636968456
transform 1 0 73324 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636968456
transform 1 0 74428 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636968456
transform 1 0 75532 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636968456
transform 1 0 76636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 1
transform 1 0 77740 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 1
transform 1 0 78292 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_841
timestamp 1636968456
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_853
timestamp 1636968456
transform 1 0 79580 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_865
timestamp 1636968456
transform 1 0 80684 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_877
timestamp 1636968456
transform 1 0 81788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_889
timestamp 1
transform 1 0 82892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 1
transform 1 0 83444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1636968456
transform 1 0 83628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_909
timestamp 1636968456
transform 1 0 84732 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_921
timestamp 1636968456
transform 1 0 85836 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_933
timestamp 1636968456
transform 1 0 86940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_945
timestamp 1
transform 1 0 88044 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_951
timestamp 1
transform 1 0 88596 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_953
timestamp 1636968456
transform 1 0 88780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_965
timestamp 1636968456
transform 1 0 89884 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_977
timestamp 1636968456
transform 1 0 90988 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_989
timestamp 1636968456
transform 1 0 92092 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1001
timestamp 1
transform 1 0 93196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1009
timestamp 1636968456
transform 1 0 93932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1021
timestamp 1636968456
transform 1 0 95036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1033
timestamp 1636968456
transform 1 0 96140 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1045
timestamp 1636968456
transform 1 0 97244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1057
timestamp 1
transform 1 0 98348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1065
timestamp 1636968456
transform 1 0 99084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1077
timestamp 1636968456
transform 1 0 100188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1089
timestamp 1636968456
transform 1 0 101292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1101
timestamp 1636968456
transform 1 0 102396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1113
timestamp 1
transform 1 0 103500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1119
timestamp 1
transform 1 0 104052 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1121
timestamp 1636968456
transform 1 0 104236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1133
timestamp 1636968456
transform 1 0 105340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1145
timestamp 1636968456
transform 1 0 106444 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1157
timestamp 1636968456
transform 1 0 107548 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1
transform 1 0 108652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1177
timestamp 1636968456
transform 1 0 109388 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1189
timestamp 1
transform 1 0 110492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636968456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636968456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636968456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636968456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636968456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636968456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636968456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636968456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636968456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636968456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636968456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636968456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636968456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636968456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636968456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636968456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636968456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636968456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636968456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636968456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636968456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636968456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636968456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636968456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636968456
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636968456
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636968456
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636968456
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636968456
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636968456
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636968456
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636968456
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636968456
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636968456
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636968456
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636968456
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636968456
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636968456
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636968456
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636968456
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636968456
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636968456
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636968456
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636968456
transform 1 0 83260 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_905
timestamp 1636968456
transform 1 0 84364 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_917
timestamp 1
transform 1 0 85468 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_923
timestamp 1
transform 1 0 86020 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_925
timestamp 1636968456
transform 1 0 86204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_937
timestamp 1636968456
transform 1 0 87308 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_949
timestamp 1636968456
transform 1 0 88412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_961
timestamp 1636968456
transform 1 0 89516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_973
timestamp 1
transform 1 0 90620 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_979
timestamp 1
transform 1 0 91172 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_981
timestamp 1636968456
transform 1 0 91356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_993
timestamp 1636968456
transform 1 0 92460 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1005
timestamp 1636968456
transform 1 0 93564 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1017
timestamp 1636968456
transform 1 0 94668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1029
timestamp 1
transform 1 0 95772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1037
timestamp 1636968456
transform 1 0 96508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1049
timestamp 1636968456
transform 1 0 97612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1061
timestamp 1636968456
transform 1 0 98716 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1073
timestamp 1636968456
transform 1 0 99820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1085
timestamp 1
transform 1 0 100924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1093
timestamp 1636968456
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1105
timestamp 1636968456
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1117
timestamp 1636968456
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1129
timestamp 1636968456
transform 1 0 104972 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1141
timestamp 1
transform 1 0 106076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1147
timestamp 1
transform 1 0 106628 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1149
timestamp 1636968456
transform 1 0 106812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1161
timestamp 1636968456
transform 1 0 107916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1173
timestamp 1636968456
transform 1 0 109020 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1185
timestamp 1
transform 1 0 110124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1189
timestamp 1
transform 1 0 110492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636968456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636968456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636968456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636968456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636968456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636968456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636968456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636968456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636968456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636968456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636968456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636968456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636968456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636968456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636968456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636968456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636968456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636968456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636968456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636968456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636968456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636968456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636968456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636968456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636968456
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636968456
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636968456
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636968456
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636968456
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636968456
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636968456
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636968456
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636968456
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636968456
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636968456
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636968456
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636968456
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636968456
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636968456
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636968456
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636968456
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636968456
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636968456
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636968456
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1636968456
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_909
timestamp 1636968456
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_921
timestamp 1636968456
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_933
timestamp 1636968456
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_953
timestamp 1636968456
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_965
timestamp 1636968456
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_977
timestamp 1636968456
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_989
timestamp 1636968456
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1009
timestamp 1636968456
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1021
timestamp 1636968456
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1033
timestamp 1636968456
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1045
timestamp 1636968456
transform 1 0 97244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1057
timestamp 1
transform 1 0 98348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1065
timestamp 1636968456
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1077
timestamp 1636968456
transform 1 0 100188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1089
timestamp 1636968456
transform 1 0 101292 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1101
timestamp 1636968456
transform 1 0 102396 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1113
timestamp 1
transform 1 0 103500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1121
timestamp 1636968456
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1133
timestamp 1636968456
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1145
timestamp 1636968456
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1157
timestamp 1636968456
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1177
timestamp 1636968456
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1189
timestamp 1
transform 1 0 110492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636968456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636968456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636968456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636968456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636968456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636968456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636968456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636968456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636968456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636968456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636968456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636968456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636968456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636968456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636968456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636968456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636968456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636968456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636968456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636968456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636968456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636968456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636968456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636968456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636968456
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636968456
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636968456
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636968456
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636968456
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636968456
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636968456
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636968456
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636968456
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636968456
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636968456
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636968456
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636968456
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636968456
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636968456
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_837
timestamp 1636968456
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_849
timestamp 1636968456
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636968456
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636968456
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_893
timestamp 1636968456
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_905
timestamp 1636968456
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_925
timestamp 1636968456
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_937
timestamp 1636968456
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_949
timestamp 1636968456
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_961
timestamp 1636968456
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_981
timestamp 1636968456
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_993
timestamp 1636968456
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1005
timestamp 1636968456
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1017
timestamp 1636968456
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1037
timestamp 1636968456
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1049
timestamp 1636968456
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1061
timestamp 1636968456
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1073
timestamp 1636968456
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1093
timestamp 1636968456
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1105
timestamp 1636968456
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1117
timestamp 1636968456
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1129
timestamp 1636968456
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1149
timestamp 1636968456
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1161
timestamp 1636968456
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1173
timestamp 1636968456
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1185
timestamp 1
transform 1 0 110124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1189
timestamp 1
transform 1 0 110492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636968456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636968456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636968456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636968456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636968456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636968456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636968456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636968456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636968456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636968456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636968456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636968456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636968456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636968456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636968456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636968456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636968456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636968456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636968456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636968456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636968456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636968456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636968456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636968456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636968456
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636968456
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636968456
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636968456
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636968456
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636968456
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636968456
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636968456
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636968456
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636968456
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636968456
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636968456
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636968456
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636968456
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1636968456
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_821
timestamp 1636968456
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_841
timestamp 1636968456
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_853
timestamp 1636968456
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_865
timestamp 1636968456
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_877
timestamp 1636968456
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1636968456
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_909
timestamp 1636968456
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_921
timestamp 1636968456
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_933
timestamp 1636968456
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_953
timestamp 1636968456
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_965
timestamp 1636968456
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_977
timestamp 1636968456
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_989
timestamp 1636968456
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1009
timestamp 1636968456
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1021
timestamp 1636968456
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1033
timestamp 1636968456
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1045
timestamp 1636968456
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1065
timestamp 1636968456
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1077
timestamp 1636968456
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1089
timestamp 1636968456
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1101
timestamp 1636968456
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1121
timestamp 1636968456
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1133
timestamp 1636968456
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1145
timestamp 1636968456
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1157
timestamp 1636968456
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1177
timestamp 1636968456
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1189
timestamp 1
transform 1 0 110492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636968456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636968456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636968456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636968456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636968456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636968456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636968456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636968456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636968456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636968456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636968456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636968456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636968456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636968456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636968456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636968456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636968456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1636968456
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1636968456
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636968456
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636968456
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1636968456
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1636968456
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636968456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636968456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1636968456
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1636968456
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636968456
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636968456
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1636968456
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1636968456
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636968456
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636968456
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1636968456
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1636968456
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636968456
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636968456
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1636968456
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1636968456
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1636968456
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_825
timestamp 1636968456
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_837
timestamp 1636968456
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_849
timestamp 1636968456
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_869
timestamp 1636968456
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_881
timestamp 1636968456
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_893
timestamp 1636968456
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_905
timestamp 1636968456
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_925
timestamp 1636968456
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_937
timestamp 1636968456
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_949
timestamp 1636968456
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_961
timestamp 1636968456
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_981
timestamp 1636968456
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_993
timestamp 1636968456
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1005
timestamp 1636968456
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1017
timestamp 1636968456
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1037
timestamp 1636968456
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1049
timestamp 1636968456
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1061
timestamp 1636968456
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1073
timestamp 1636968456
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1093
timestamp 1636968456
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1105
timestamp 1636968456
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1117
timestamp 1636968456
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1129
timestamp 1636968456
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1149
timestamp 1636968456
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1161
timestamp 1636968456
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1173
timestamp 1636968456
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1185
timestamp 1
transform 1 0 110124 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1189
timestamp 1
transform 1 0 110492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636968456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636968456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636968456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636968456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636968456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636968456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636968456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636968456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636968456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636968456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636968456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636968456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636968456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636968456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636968456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636968456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636968456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636968456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1636968456
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1636968456
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1636968456
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636968456
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636968456
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636968456
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636968456
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1636968456
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1636968456
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1636968456
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1636968456
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1636968456
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1636968456
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1636968456
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1636968456
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1636968456
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1636968456
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1636968456
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1636968456
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1636968456
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1636968456
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1636968456
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1636968456
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1636968456
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1636968456
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1636968456
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1636968456
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_841
timestamp 1636968456
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_853
timestamp 1636968456
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_865
timestamp 1636968456
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_877
timestamp 1636968456
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1636968456
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_909
timestamp 1636968456
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_921
timestamp 1636968456
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_933
timestamp 1636968456
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_953
timestamp 1636968456
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_965
timestamp 1636968456
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_977
timestamp 1636968456
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_989
timestamp 1636968456
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1009
timestamp 1636968456
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1021
timestamp 1636968456
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1033
timestamp 1636968456
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1045
timestamp 1636968456
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1065
timestamp 1636968456
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1077
timestamp 1636968456
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1089
timestamp 1636968456
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1101
timestamp 1636968456
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1121
timestamp 1636968456
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1133
timestamp 1636968456
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1145
timestamp 1636968456
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1157
timestamp 1636968456
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1177
timestamp 1636968456
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1189
timestamp 1
transform 1 0 110492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636968456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636968456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636968456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636968456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636968456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636968456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636968456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636968456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636968456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636968456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636968456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636968456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636968456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636968456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636968456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636968456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636968456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636968456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636968456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636968456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636968456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636968456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636968456
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636968456
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636968456
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636968456
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636968456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636968456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1636968456
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1636968456
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1636968456
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1636968456
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1636968456
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1636968456
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1636968456
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1636968456
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1636968456
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1636968456
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1636968456
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1636968456
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1636968456
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1636968456
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1636968456
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1636968456
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1636968456
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1636968456
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1636968456
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_825
timestamp 1636968456
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_837
timestamp 1636968456
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_849
timestamp 1636968456
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_869
timestamp 1636968456
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_881
timestamp 1636968456
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_893
timestamp 1636968456
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_905
timestamp 1636968456
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_925
timestamp 1636968456
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_937
timestamp 1636968456
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_949
timestamp 1636968456
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_961
timestamp 1636968456
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_981
timestamp 1636968456
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_993
timestamp 1636968456
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1005
timestamp 1636968456
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1017
timestamp 1636968456
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1037
timestamp 1636968456
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1049
timestamp 1636968456
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1061
timestamp 1636968456
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1073
timestamp 1636968456
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1093
timestamp 1636968456
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1105
timestamp 1636968456
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1117
timestamp 1636968456
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1129
timestamp 1636968456
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1149
timestamp 1636968456
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1161
timestamp 1636968456
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1173
timestamp 1636968456
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1185
timestamp 1
transform 1 0 110124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1189
timestamp 1
transform 1 0 110492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_29
timestamp 1636968456
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_41
timestamp 1636968456
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_81
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1636968456
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1636968456
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_141
timestamp 1636968456
transform 1 0 14076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_153
timestamp 1
transform 1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636968456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1636968456
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1636968456
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1
transform 1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_245
timestamp 1
transform 1 0 23644 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_251
timestamp 1
transform 1 0 24196 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_253
timestamp 1
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_258
timestamp 1
transform 1 0 24840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_266
timestamp 1
transform 1 0 25576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_283
timestamp 1
transform 1 0 27140 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_291
timestamp 1
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_296
timestamp 1636968456
transform 1 0 28336 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_311
timestamp 1
transform 1 0 29716 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_321
timestamp 1
transform 1 0 30636 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_329
timestamp 1
transform 1 0 31372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_337
timestamp 1
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_347
timestamp 1
transform 1 0 33028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_355
timestamp 1
transform 1 0 33764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_359
timestamp 1
transform 1 0 34132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_363
timestamp 1
transform 1 0 34500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_365
timestamp 1
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_369
timestamp 1
transform 1 0 35052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_372
timestamp 1
transform 1 0 35328 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_380
timestamp 1
transform 1 0 36064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_397
timestamp 1
transform 1 0 37628 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_405
timestamp 1
transform 1 0 38364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_410
timestamp 1
transform 1 0 38824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_418
timestamp 1
transform 1 0 39560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_423
timestamp 1
transform 1 0 40020 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_431
timestamp 1
transform 1 0 40756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_436
timestamp 1
transform 1 0 41216 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_444
timestamp 1
transform 1 0 41952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_449
timestamp 1
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_457
timestamp 1
transform 1 0 43148 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636968456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_473
timestamp 1
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_477
timestamp 1636968456
transform 1 0 44988 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_489
timestamp 1636968456
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636968456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636968456
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_529
timestamp 1
transform 1 0 49772 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_533
timestamp 1636968456
transform 1 0 50140 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_545
timestamp 1636968456
transform 1 0 51244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_557
timestamp 1
transform 1 0 52348 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1636968456
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1636968456
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_585
timestamp 1
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_589
timestamp 1636968456
transform 1 0 55292 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_601
timestamp 1636968456
transform 1 0 56396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_613
timestamp 1
transform 1 0 57500 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1636968456
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1636968456
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_641
timestamp 1
transform 1 0 60076 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_645
timestamp 1636968456
transform 1 0 60444 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_657
timestamp 1636968456
transform 1 0 61548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_669
timestamp 1
transform 1 0 62652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1636968456
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1636968456
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_697
timestamp 1
transform 1 0 65228 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_701
timestamp 1636968456
transform 1 0 65596 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_713
timestamp 1636968456
transform 1 0 66700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_725
timestamp 1
transform 1 0 67804 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1636968456
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1636968456
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_753
timestamp 1
transform 1 0 70380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_757
timestamp 1636968456
transform 1 0 70748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_769
timestamp 1636968456
transform 1 0 71852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_781
timestamp 1
transform 1 0 72956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1636968456
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1636968456
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_809
timestamp 1
transform 1 0 75532 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_813
timestamp 1636968456
transform 1 0 75900 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_825
timestamp 1636968456
transform 1 0 77004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_837
timestamp 1
transform 1 0 78108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_841
timestamp 1636968456
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_853
timestamp 1636968456
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_865
timestamp 1
transform 1 0 80684 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_869
timestamp 1636968456
transform 1 0 81052 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_881
timestamp 1636968456
transform 1 0 82156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_893
timestamp 1
transform 1 0 83260 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1636968456
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_909
timestamp 1636968456
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_921
timestamp 1
transform 1 0 85836 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_925
timestamp 1636968456
transform 1 0 86204 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_937
timestamp 1636968456
transform 1 0 87308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_949
timestamp 1
transform 1 0 88412 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_953
timestamp 1636968456
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_965
timestamp 1
transform 1 0 89884 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_971
timestamp 1
transform 1 0 90436 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_978
timestamp 1
transform 1 0 91080 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_981
timestamp 1636968456
transform 1 0 91356 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_993
timestamp 1636968456
transform 1 0 92460 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1005
timestamp 1
transform 1 0 93564 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1009
timestamp 1636968456
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1021
timestamp 1636968456
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1033
timestamp 1
transform 1 0 96140 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1037
timestamp 1636968456
transform 1 0 96508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1049
timestamp 1636968456
transform 1 0 97612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1061
timestamp 1
transform 1 0 98716 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1065
timestamp 1636968456
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1077
timestamp 1636968456
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1089
timestamp 1
transform 1 0 101292 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1093
timestamp 1636968456
transform 1 0 101660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1105
timestamp 1636968456
transform 1 0 102764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1117
timestamp 1
transform 1 0 103868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1121
timestamp 1636968456
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1133
timestamp 1636968456
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1145
timestamp 1
transform 1 0 106444 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1149
timestamp 1636968456
transform 1 0 106812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1161
timestamp 1636968456
transform 1 0 107916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_1173
timestamp 1
transform 1 0 109020 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1177
timestamp 1636968456
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1189
timestamp 1
transform 1 0 110492 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636968456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1122
timestamp 1636968456
transform 1 0 104328 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1134
timestamp 1636968456
transform 1 0 105432 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1146
timestamp 1
transform 1 0 106536 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1148
timestamp 1636968456
transform 1 0 106720 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1160
timestamp 1636968456
transform 1 0 107824 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1172
timestamp 1636968456
transform 1 0 108928 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1184
timestamp 1
transform 1 0 110032 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636968456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1122
timestamp 1636968456
transform 1 0 104328 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1134
timestamp 1636968456
transform 1 0 105432 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1146
timestamp 1636968456
transform 1 0 106536 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1158
timestamp 1636968456
transform 1 0 107640 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_1170
timestamp 1
transform 1 0 108744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1174
timestamp 1
transform 1 0 109112 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1176
timestamp 1636968456
transform 1 0 109296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_1188
timestamp 1
transform 1 0 110400 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636968456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_65
timestamp 1
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1122
timestamp 1636968456
transform 1 0 104328 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1134
timestamp 1636968456
transform 1 0 105432 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1146
timestamp 1
transform 1 0 106536 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1148
timestamp 1636968456
transform 1 0 106720 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1160
timestamp 1636968456
transform 1 0 107824 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1172
timestamp 1636968456
transform 1 0 108928 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1184
timestamp 1
transform 1 0 110032 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp 1
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1122
timestamp 1636968456
transform 1 0 104328 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1134
timestamp 1636968456
transform 1 0 105432 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1146
timestamp 1636968456
transform 1 0 106536 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1158
timestamp 1636968456
transform 1 0 107640 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_1170
timestamp 1
transform 1 0 108744 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1174
timestamp 1
transform 1 0 109112 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1176
timestamp 1636968456
transform 1 0 109296 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_1188
timestamp 1
transform 1 0 110400 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636968456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636968456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1122
timestamp 1636968456
transform 1 0 104328 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1134
timestamp 1636968456
transform 1 0 105432 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1146
timestamp 1
transform 1 0 106536 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1148
timestamp 1636968456
transform 1 0 106720 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1160
timestamp 1636968456
transform 1 0 107824 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1172
timestamp 1636968456
transform 1 0 108928 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1184
timestamp 1
transform 1 0 110032 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636968456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636968456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636968456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1122
timestamp 1636968456
transform 1 0 104328 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1134
timestamp 1636968456
transform 1 0 105432 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1146
timestamp 1636968456
transform 1 0 106536 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1158
timestamp 1636968456
transform 1 0 107640 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_1170
timestamp 1
transform 1 0 108744 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1174
timestamp 1
transform 1 0 109112 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1176
timestamp 1636968456
transform 1 0 109296 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_1188
timestamp 1
transform 1 0 110400 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636968456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636968456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_65
timestamp 1
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1122
timestamp 1636968456
transform 1 0 104328 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1134
timestamp 1636968456
transform 1 0 105432 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1146
timestamp 1
transform 1 0 106536 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1148
timestamp 1636968456
transform 1 0 106720 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1160
timestamp 1636968456
transform 1 0 107824 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1172
timestamp 1636968456
transform 1 0 108928 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1184
timestamp 1
transform 1 0 110032 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636968456
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636968456
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636968456
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1122
timestamp 1636968456
transform 1 0 104328 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1134
timestamp 1636968456
transform 1 0 105432 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1146
timestamp 1636968456
transform 1 0 106536 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1158
timestamp 1636968456
transform 1 0 107640 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1170
timestamp 1
transform 1 0 108744 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1174
timestamp 1
transform 1 0 109112 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1176
timestamp 1636968456
transform 1 0 109296 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1188
timestamp 1
transform 1 0 110400 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636968456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636968456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_65
timestamp 1
transform 1 0 7084 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1122
timestamp 1636968456
transform 1 0 104328 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1134
timestamp 1636968456
transform 1 0 105432 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1146
timestamp 1
transform 1 0 106536 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1148
timestamp 1636968456
transform 1 0 106720 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1160
timestamp 1636968456
transform 1 0 107824 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1172
timestamp 1636968456
transform 1 0 108928 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1184
timestamp 1
transform 1 0 110032 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636968456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636968456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636968456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636968456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1122
timestamp 1636968456
transform 1 0 104328 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1134
timestamp 1636968456
transform 1 0 105432 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1146
timestamp 1636968456
transform 1 0 106536 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1158
timestamp 1636968456
transform 1 0 107640 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1170
timestamp 1
transform 1 0 108744 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1174
timestamp 1
transform 1 0 109112 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1176
timestamp 1636968456
transform 1 0 109296 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1188
timestamp 1
transform 1 0 110400 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636968456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636968456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636968456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_65
timestamp 1
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1122
timestamp 1636968456
transform 1 0 104328 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1134
timestamp 1636968456
transform 1 0 105432 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1146
timestamp 1
transform 1 0 106536 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1148
timestamp 1636968456
transform 1 0 106720 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1160
timestamp 1636968456
transform 1 0 107824 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1172
timestamp 1636968456
transform 1 0 108928 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1184
timestamp 1
transform 1 0 110032 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636968456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636968456
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636968456
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636968456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1122
timestamp 1636968456
transform 1 0 104328 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1134
timestamp 1636968456
transform 1 0 105432 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1146
timestamp 1636968456
transform 1 0 106536 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1158
timestamp 1636968456
transform 1 0 107640 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_1170
timestamp 1
transform 1 0 108744 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1174
timestamp 1
transform 1 0 109112 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1176
timestamp 1636968456
transform 1 0 109296 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_1188
timestamp 1
transform 1 0 110400 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636968456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_65
timestamp 1
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1122
timestamp 1636968456
transform 1 0 104328 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1134
timestamp 1636968456
transform 1 0 105432 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1146
timestamp 1
transform 1 0 106536 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1148
timestamp 1636968456
transform 1 0 106720 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1160
timestamp 1636968456
transform 1 0 107824 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1172
timestamp 1636968456
transform 1 0 108928 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1184
timestamp 1
transform 1 0 110032 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636968456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636968456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1122
timestamp 1636968456
transform 1 0 104328 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1134
timestamp 1636968456
transform 1 0 105432 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1146
timestamp 1636968456
transform 1 0 106536 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1158
timestamp 1636968456
transform 1 0 107640 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_1170
timestamp 1
transform 1 0 108744 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1174
timestamp 1
transform 1 0 109112 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1176
timestamp 1636968456
transform 1 0 109296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_1188
timestamp 1
transform 1 0 110400 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636968456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1122
timestamp 1636968456
transform 1 0 104328 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1134
timestamp 1636968456
transform 1 0 105432 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1146
timestamp 1
transform 1 0 106536 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1148
timestamp 1636968456
transform 1 0 106720 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1160
timestamp 1636968456
transform 1 0 107824 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1172
timestamp 1636968456
transform 1 0 108928 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1184
timestamp 1
transform 1 0 110032 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636968456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636968456
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636968456
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1122
timestamp 1636968456
transform 1 0 104328 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1134
timestamp 1636968456
transform 1 0 105432 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1146
timestamp 1636968456
transform 1 0 106536 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1158
timestamp 1636968456
transform 1 0 107640 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_1170
timestamp 1
transform 1 0 108744 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1174
timestamp 1
transform 1 0 109112 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1176
timestamp 1636968456
transform 1 0 109296 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_1188
timestamp 1
transform 1 0 110400 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1122
timestamp 1636968456
transform 1 0 104328 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1134
timestamp 1636968456
transform 1 0 105432 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1146
timestamp 1
transform 1 0 106536 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1148
timestamp 1636968456
transform 1 0 106720 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1160
timestamp 1636968456
transform 1 0 107824 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1172
timestamp 1636968456
transform 1 0 108928 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1184
timestamp 1
transform 1 0 110032 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636968456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636968456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1122
timestamp 1636968456
transform 1 0 104328 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1134
timestamp 1636968456
transform 1 0 105432 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1146
timestamp 1636968456
transform 1 0 106536 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1158
timestamp 1636968456
transform 1 0 107640 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_1170
timestamp 1
transform 1 0 108744 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1174
timestamp 1
transform 1 0 109112 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1176
timestamp 1636968456
transform 1 0 109296 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_1188
timestamp 1
transform 1 0 110400 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636968456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_65
timestamp 1
transform 1 0 7084 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1122
timestamp 1636968456
transform 1 0 104328 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1134
timestamp 1636968456
transform 1 0 105432 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1146
timestamp 1
transform 1 0 106536 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1148
timestamp 1636968456
transform 1 0 106720 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1160
timestamp 1636968456
transform 1 0 107824 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1172
timestamp 1636968456
transform 1 0 108928 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1184
timestamp 1
transform 1 0 110032 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636968456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636968456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636968456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636968456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1122
timestamp 1636968456
transform 1 0 104328 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1134
timestamp 1636968456
transform 1 0 105432 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1146
timestamp 1636968456
transform 1 0 106536 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1158
timestamp 1636968456
transform 1 0 107640 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_1170
timestamp 1
transform 1 0 108744 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1174
timestamp 1
transform 1 0 109112 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1176
timestamp 1636968456
transform 1 0 109296 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_1188
timestamp 1
transform 1 0 110400 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636968456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636968456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636968456
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1122
timestamp 1636968456
transform 1 0 104328 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1134
timestamp 1636968456
transform 1 0 105432 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1146
timestamp 1
transform 1 0 106536 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1148
timestamp 1636968456
transform 1 0 106720 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1160
timestamp 1636968456
transform 1 0 107824 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1172
timestamp 1636968456
transform 1 0 108928 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1184
timestamp 1
transform 1 0 110032 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636968456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636968456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636968456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636968456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636968456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_69
timestamp 1
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1129
timestamp 1636968456
transform 1 0 104972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1141
timestamp 1636968456
transform 1 0 106076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1153
timestamp 1636968456
transform 1 0 107180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1165
timestamp 1
transform 1 0 108284 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1173
timestamp 1
transform 1 0 109020 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1176
timestamp 1636968456
transform 1 0 109296 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1188
timestamp 1
transform 1 0 110400 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636968456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636968456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636968456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636968456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636968456
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 1
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1124
timestamp 1636968456
transform 1 0 104512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_1136
timestamp 1
transform 1 0 105616 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_1144
timestamp 1
transform 1 0 106352 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1148
timestamp 1636968456
transform 1 0 106720 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1160
timestamp 1636968456
transform 1 0 107824 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_1172
timestamp 1636968456
transform 1 0 108928 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1184
timestamp 1
transform 1 0 110032 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636968456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636968456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636968456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636968456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1122
timestamp 1
transform 1 0 104328 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1131
timestamp 1636968456
transform 1 0 105156 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1143
timestamp 1636968456
transform 1 0 106260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1155
timestamp 1636968456
transform 1 0 107364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_1167
timestamp 1
transform 1 0 108468 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1176
timestamp 1636968456
transform 1 0 109296 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_1188
timestamp 1
transform 1 0 110400 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636968456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636968456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636968456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636968456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636968456
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_65
timestamp 1
transform 1 0 7084 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1146
timestamp 1
transform 1 0 106536 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1148
timestamp 1636968456
transform 1 0 106720 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1160
timestamp 1636968456
transform 1 0 107824 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1172
timestamp 1636968456
transform 1 0 108928 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1184
timestamp 1
transform 1 0 110032 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636968456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636968456
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636968456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636968456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1122
timestamp 1636968456
transform 1 0 104328 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1134
timestamp 1636968456
transform 1 0 105432 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1146
timestamp 1636968456
transform 1 0 106536 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1158
timestamp 1636968456
transform 1 0 107640 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_1170
timestamp 1
transform 1 0 108744 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1174
timestamp 1
transform 1 0 109112 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1176
timestamp 1636968456
transform 1 0 109296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_1188
timestamp 1
transform 1 0 110400 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636968456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636968456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636968456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636968456
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_65
timestamp 1
transform 1 0 7084 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1122
timestamp 1636968456
transform 1 0 104328 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1134
timestamp 1636968456
transform 1 0 105432 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1146
timestamp 1
transform 1 0 106536 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1148
timestamp 1636968456
transform 1 0 106720 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1160
timestamp 1636968456
transform 1 0 107824 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1172
timestamp 1636968456
transform 1 0 108928 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1184
timestamp 1
transform 1 0 110032 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636968456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636968456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636968456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636968456
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636968456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1122
timestamp 1636968456
transform 1 0 104328 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1134
timestamp 1636968456
transform 1 0 105432 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1146
timestamp 1636968456
transform 1 0 106536 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1158
timestamp 1636968456
transform 1 0 107640 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_1170
timestamp 1
transform 1 0 108744 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1174
timestamp 1
transform 1 0 109112 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_1176
timestamp 1636968456
transform 1 0 109296 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_1188
timestamp 1
transform 1 0 110400 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636968456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636968456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636968456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636968456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1122
timestamp 1636968456
transform 1 0 104328 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1134
timestamp 1636968456
transform 1 0 105432 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1146
timestamp 1
transform 1 0 106536 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1148
timestamp 1636968456
transform 1 0 106720 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1160
timestamp 1636968456
transform 1 0 107824 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1172
timestamp 1636968456
transform 1 0 108928 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1184
timestamp 1
transform 1 0 110032 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636968456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636968456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636968456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636968456
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636968456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_69
timestamp 1
transform 1 0 7452 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1134
timestamp 1636968456
transform 1 0 105432 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1146
timestamp 1636968456
transform 1 0 106536 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1158
timestamp 1636968456
transform 1 0 107640 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_1170
timestamp 1
transform 1 0 108744 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1174
timestamp 1
transform 1 0 109112 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1176
timestamp 1636968456
transform 1 0 109296 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_1188
timestamp 1
transform 1 0 110400 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636968456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636968456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636968456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636968456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_65
timestamp 1
transform 1 0 7084 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1130
timestamp 1636968456
transform 1 0 105064 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_1142
timestamp 1
transform 1 0 106168 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1146
timestamp 1
transform 1 0 106536 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1148
timestamp 1636968456
transform 1 0 106720 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1160
timestamp 1636968456
transform 1 0 107824 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1172
timestamp 1636968456
transform 1 0 108928 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1184
timestamp 1
transform 1 0 110032 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636968456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636968456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636968456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636968456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1124
timestamp 1636968456
transform 1 0 104512 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1136
timestamp 1636968456
transform 1 0 105616 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1148
timestamp 1636968456
transform 1 0 106720 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1160
timestamp 1636968456
transform 1 0 107824 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_1172
timestamp 1
transform 1 0 108928 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_1176
timestamp 1636968456
transform 1 0 109296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_1188
timestamp 1
transform 1 0 110400 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636968456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636968456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636968456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636968456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1134
timestamp 1636968456
transform 1 0 105432 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1146
timestamp 1
transform 1 0 106536 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1148
timestamp 1636968456
transform 1 0 106720 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1160
timestamp 1636968456
transform 1 0 107824 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_1172
timestamp 1636968456
transform 1 0 108928 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1184
timestamp 1
transform 1 0 110032 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636968456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636968456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1146
timestamp 1636968456
transform 1 0 106536 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1158
timestamp 1636968456
transform 1 0 107640 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_1170
timestamp 1
transform 1 0 108744 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1174
timestamp 1
transform 1 0 109112 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_1176
timestamp 1636968456
transform 1 0 109296 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_1188
timestamp 1
transform 1 0 110400 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636968456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636968456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636968456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636968456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636968456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_65
timestamp 1
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1122
timestamp 1636968456
transform 1 0 104328 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1134
timestamp 1636968456
transform 1 0 105432 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1146
timestamp 1
transform 1 0 106536 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1148
timestamp 1636968456
transform 1 0 106720 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1160
timestamp 1636968456
transform 1 0 107824 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1172
timestamp 1636968456
transform 1 0 108928 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1184
timestamp 1
transform 1 0 110032 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636968456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636968456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636968456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636968456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636968456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1122
timestamp 1
transform 1 0 104328 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1135
timestamp 1636968456
transform 1 0 105524 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1147
timestamp 1636968456
transform 1 0 106628 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1159
timestamp 1636968456
transform 1 0 107732 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1171
timestamp 1
transform 1 0 108836 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1176
timestamp 1636968456
transform 1 0 109296 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1188
timestamp 1
transform 1 0 110400 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636968456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636968456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_65
timestamp 1
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1122
timestamp 1636968456
transform 1 0 104328 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1134
timestamp 1636968456
transform 1 0 105432 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1146
timestamp 1
transform 1 0 106536 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1148
timestamp 1636968456
transform 1 0 106720 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1160
timestamp 1636968456
transform 1 0 107824 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_1172
timestamp 1636968456
transform 1 0 108928 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1184
timestamp 1
transform 1 0 110032 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_69
timestamp 1
transform 1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_1122
timestamp 1
transform 1 0 104328 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1132
timestamp 1636968456
transform 1 0 105248 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1144
timestamp 1636968456
transform 1 0 106352 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1156
timestamp 1636968456
transform 1 0 107456 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1168
timestamp 1
transform 1 0 108560 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1174
timestamp 1
transform 1 0 109112 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1176
timestamp 1636968456
transform 1 0 109296 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_1188
timestamp 1
transform 1 0 110400 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636968456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_65
timestamp 1
transform 1 0 7084 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1148
timestamp 1636968456
transform 1 0 106720 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1160
timestamp 1636968456
transform 1 0 107824 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1172
timestamp 1636968456
transform 1 0 108928 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1184
timestamp 1
transform 1 0 110032 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636968456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636968456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1636968456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1636968456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636968456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1
transform 1 0 7452 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1122
timestamp 1636968456
transform 1 0 104328 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1134
timestamp 1636968456
transform 1 0 105432 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1146
timestamp 1636968456
transform 1 0 106536 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1158
timestamp 1636968456
transform 1 0 107640 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_1170
timestamp 1
transform 1 0 108744 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1174
timestamp 1
transform 1 0 109112 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_1176
timestamp 1636968456
transform 1 0 109296 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_1188
timestamp 1
transform 1 0 110400 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636968456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636968456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636968456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636968456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636968456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_65
timestamp 1
transform 1 0 7084 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1127
timestamp 1636968456
transform 1 0 104788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1139
timestamp 1
transform 1 0 105892 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1148
timestamp 1636968456
transform 1 0 106720 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1160
timestamp 1636968456
transform 1 0 107824 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1172
timestamp 1636968456
transform 1 0 108928 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1184
timestamp 1
transform 1 0 110032 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636968456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636968456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636968456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636968456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636968456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_69
timestamp 1
transform 1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_1122
timestamp 1
transform 1 0 104328 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1126
timestamp 1
transform 1 0 104696 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1139
timestamp 1636968456
transform 1 0 105892 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1151
timestamp 1636968456
transform 1 0 106996 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1163
timestamp 1636968456
transform 1 0 108100 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1176
timestamp 1636968456
transform 1 0 109296 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_1188
timestamp 1
transform 1 0 110400 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636968456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636968456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636968456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636968456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1636968456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_65
timestamp 1
transform 1 0 7084 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1122
timestamp 1636968456
transform 1 0 104328 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1134
timestamp 1636968456
transform 1 0 105432 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1146
timestamp 1
transform 1 0 106536 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1148
timestamp 1636968456
transform 1 0 106720 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1160
timestamp 1636968456
transform 1 0 107824 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_1172
timestamp 1636968456
transform 1 0 108928 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1184
timestamp 1
transform 1 0 110032 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636968456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636968456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636968456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1636968456
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636968456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_69
timestamp 1
transform 1 0 7452 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_1122
timestamp 1
transform 1 0 104328 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1127
timestamp 1636968456
transform 1 0 104788 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1139
timestamp 1636968456
transform 1 0 105892 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1151
timestamp 1636968456
transform 1 0 106996 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1163
timestamp 1636968456
transform 1 0 108100 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1176
timestamp 1636968456
transform 1 0 109296 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_1188
timestamp 1
transform 1 0 110400 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636968456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636968456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636968456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1636968456
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1636968456
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_65
timestamp 1
transform 1 0 7084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1125
timestamp 1
transform 1 0 104604 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_1143
timestamp 1
transform 1 0 106260 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1148
timestamp 1636968456
transform 1 0 106720 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1160
timestamp 1636968456
transform 1 0 107824 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_1172
timestamp 1636968456
transform 1 0 108928 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1184
timestamp 1
transform 1 0 110032 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636968456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636968456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1636968456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1636968456
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1636968456
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_69
timestamp 1
transform 1 0 7452 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1135
timestamp 1636968456
transform 1 0 105524 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1147
timestamp 1636968456
transform 1 0 106628 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1159
timestamp 1636968456
transform 1 0 107732 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_1171
timestamp 1
transform 1 0 108836 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1176
timestamp 1636968456
transform 1 0 109296 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_1188
timestamp 1
transform 1 0 110400 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636968456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636968456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636968456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636968456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1636968456
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_65
timestamp 1
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_56_1144
timestamp 1
transform 1 0 106352 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1148
timestamp 1636968456
transform 1 0 106720 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1160
timestamp 1636968456
transform 1 0 107824 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1172
timestamp 1636968456
transform 1 0 108928 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1184
timestamp 1
transform 1 0 110032 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636968456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636968456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636968456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636968456
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636968456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_69
timestamp 1
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_1122
timestamp 1
transform 1 0 104328 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1134
timestamp 1636968456
transform 1 0 105432 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1146
timestamp 1636968456
transform 1 0 106536 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1158
timestamp 1636968456
transform 1 0 107640 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_1170
timestamp 1
transform 1 0 108744 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1174
timestamp 1
transform 1 0 109112 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1176
timestamp 1636968456
transform 1 0 109296 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_1188
timestamp 1
transform 1 0 110400 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636968456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636968456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636968456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636968456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636968456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_65
timestamp 1
transform 1 0 7084 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_1144
timestamp 1
transform 1 0 106352 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1148
timestamp 1636968456
transform 1 0 106720 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1160
timestamp 1636968456
transform 1 0 107824 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1172
timestamp 1636968456
transform 1 0 108928 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1184
timestamp 1
transform 1 0 110032 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636968456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636968456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636968456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636968456
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636968456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_69
timestamp 1
transform 1 0 7452 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1122
timestamp 1636968456
transform 1 0 104328 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1134
timestamp 1636968456
transform 1 0 105432 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1146
timestamp 1636968456
transform 1 0 106536 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1158
timestamp 1636968456
transform 1 0 107640 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_1170
timestamp 1
transform 1 0 108744 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1174
timestamp 1
transform 1 0 109112 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1176
timestamp 1636968456
transform 1 0 109296 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1188
timestamp 1
transform 1 0 110400 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636968456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636968456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636968456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636968456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636968456
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_65
timestamp 1
transform 1 0 7084 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1122
timestamp 1636968456
transform 1 0 104328 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1134
timestamp 1636968456
transform 1 0 105432 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1146
timestamp 1
transform 1 0 106536 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1148
timestamp 1636968456
transform 1 0 106720 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1160
timestamp 1636968456
transform 1 0 107824 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1172
timestamp 1636968456
transform 1 0 108928 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1184
timestamp 1
transform 1 0 110032 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636968456
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636968456
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1636968456
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1636968456
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636968456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1127
timestamp 1636968456
transform 1 0 104788 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1139
timestamp 1636968456
transform 1 0 105892 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1151
timestamp 1636968456
transform 1 0 106996 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1163
timestamp 1636968456
transform 1 0 108100 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1176
timestamp 1636968456
transform 1 0 109296 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1188
timestamp 1
transform 1 0 110400 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636968456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636968456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636968456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636968456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1636968456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_65
timestamp 1
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1122
timestamp 1636968456
transform 1 0 104328 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1134
timestamp 1636968456
transform 1 0 105432 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1146
timestamp 1
transform 1 0 106536 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1148
timestamp 1636968456
transform 1 0 106720 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1160
timestamp 1636968456
transform 1 0 107824 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1172
timestamp 1636968456
transform 1 0 108928 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1184
timestamp 1
transform 1 0 110032 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636968456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636968456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1636968456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1636968456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1636968456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1127
timestamp 1636968456
transform 1 0 104788 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1139
timestamp 1636968456
transform 1 0 105892 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1151
timestamp 1636968456
transform 1 0 106996 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1163
timestamp 1636968456
transform 1 0 108100 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1176
timestamp 1636968456
transform 1 0 109296 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1188
timestamp 1
transform 1 0 110400 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636968456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636968456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636968456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1636968456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1636968456
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_65
timestamp 1
transform 1 0 7084 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1122
timestamp 1636968456
transform 1 0 104328 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1134
timestamp 1636968456
transform 1 0 105432 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1146
timestamp 1
transform 1 0 106536 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1148
timestamp 1636968456
transform 1 0 106720 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1160
timestamp 1636968456
transform 1 0 107824 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1172
timestamp 1636968456
transform 1 0 108928 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1184
timestamp 1
transform 1 0 110032 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1636968456
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1636968456
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1636968456
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1636968456
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1636968456
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_69
timestamp 1
transform 1 0 7452 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1122
timestamp 1636968456
transform 1 0 104328 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1134
timestamp 1636968456
transform 1 0 105432 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1146
timestamp 1636968456
transform 1 0 106536 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1158
timestamp 1636968456
transform 1 0 107640 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_1170
timestamp 1
transform 1 0 108744 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1174
timestamp 1
transform 1 0 109112 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1176
timestamp 1636968456
transform 1 0 109296 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_1188
timestamp 1
transform 1 0 110400 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636968456
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636968456
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636968456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1636968456
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1636968456
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_65
timestamp 1
transform 1 0 7084 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1122
timestamp 1636968456
transform 1 0 104328 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1134
timestamp 1636968456
transform 1 0 105432 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1146
timestamp 1
transform 1 0 106536 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1148
timestamp 1636968456
transform 1 0 106720 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1160
timestamp 1636968456
transform 1 0 107824 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1172
timestamp 1636968456
transform 1 0 108928 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_1184
timestamp 1
transform 1 0 110032 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636968456
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636968456
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1636968456
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1636968456
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636968456
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1122
timestamp 1636968456
transform 1 0 104328 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1134
timestamp 1636968456
transform 1 0 105432 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1146
timestamp 1636968456
transform 1 0 106536 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1158
timestamp 1636968456
transform 1 0 107640 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_1170
timestamp 1
transform 1 0 108744 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_1174
timestamp 1
transform 1 0 109112 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1176
timestamp 1636968456
transform 1 0 109296 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_1188
timestamp 1
transform 1 0 110400 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636968456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636968456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636968456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636968456
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636968456
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_65
timestamp 1
transform 1 0 7084 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1122
timestamp 1636968456
transform 1 0 104328 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1134
timestamp 1636968456
transform 1 0 105432 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1146
timestamp 1
transform 1 0 106536 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1148
timestamp 1636968456
transform 1 0 106720 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1160
timestamp 1636968456
transform 1 0 107824 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1172
timestamp 1636968456
transform 1 0 108928 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_1184
timestamp 1
transform 1 0 110032 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636968456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636968456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636968456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636968456
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636968456
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1122
timestamp 1636968456
transform 1 0 104328 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1134
timestamp 1636968456
transform 1 0 105432 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1146
timestamp 1636968456
transform 1 0 106536 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1158
timestamp 1636968456
transform 1 0 107640 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_1170
timestamp 1
transform 1 0 108744 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_1174
timestamp 1
transform 1 0 109112 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1176
timestamp 1636968456
transform 1 0 109296 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_1188
timestamp 1
transform 1 0 110400 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636968456
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636968456
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636968456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636968456
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636968456
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_65
timestamp 1
transform 1 0 7084 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1122
timestamp 1636968456
transform 1 0 104328 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1134
timestamp 1636968456
transform 1 0 105432 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1146
timestamp 1
transform 1 0 106536 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1148
timestamp 1636968456
transform 1 0 106720 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1160
timestamp 1636968456
transform 1 0 107824 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1172
timestamp 1636968456
transform 1 0 108928 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_1184
timestamp 1
transform 1 0 110032 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636968456
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636968456
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636968456
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636968456
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636968456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_69
timestamp 1
transform 1 0 7452 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1129
timestamp 1636968456
transform 1 0 104972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1141
timestamp 1636968456
transform 1 0 106076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1153
timestamp 1636968456
transform 1 0 107180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_1165
timestamp 1
transform 1 0 108284 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1173
timestamp 1
transform 1 0 109020 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_1176
timestamp 1636968456
transform 1 0 109296 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1188
timestamp 1
transform 1 0 110400 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636968456
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636968456
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636968456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636968456
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636968456
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_65
timestamp 1
transform 1 0 7084 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_1144
timestamp 1
transform 1 0 106352 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1148
timestamp 1636968456
transform 1 0 106720 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1160
timestamp 1636968456
transform 1 0 107824 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1172
timestamp 1636968456
transform 1 0 108928 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_1184
timestamp 1
transform 1 0 110032 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636968456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636968456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636968456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636968456
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636968456
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_69
timestamp 1
transform 1 0 7452 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1148
timestamp 1636968456
transform 1 0 106720 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1160
timestamp 1636968456
transform 1 0 107824 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_1172
timestamp 1
transform 1 0 108928 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1176
timestamp 1636968456
transform 1 0 109296 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_1188
timestamp 1
transform 1 0 110400 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636968456
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636968456
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636968456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636968456
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636968456
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_65
timestamp 1
transform 1 0 7084 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1146
timestamp 1
transform 1 0 106536 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1148
timestamp 1636968456
transform 1 0 106720 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1160
timestamp 1636968456
transform 1 0 107824 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1172
timestamp 1636968456
transform 1 0 108928 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_1184
timestamp 1
transform 1 0 110032 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636968456
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636968456
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1636968456
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1636968456
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636968456
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_69
timestamp 1
transform 1 0 7452 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1122
timestamp 1636968456
transform 1 0 104328 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1134
timestamp 1636968456
transform 1 0 105432 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1146
timestamp 1636968456
transform 1 0 106536 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1158
timestamp 1636968456
transform 1 0 107640 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_1170
timestamp 1
transform 1 0 108744 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_1174
timestamp 1
transform 1 0 109112 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1176
timestamp 1636968456
transform 1 0 109296 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_1188
timestamp 1
transform 1 0 110400 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636968456
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636968456
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636968456
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1636968456
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1636968456
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_65
timestamp 1
transform 1 0 7084 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1127
timestamp 1636968456
transform 1 0 104788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_1139
timestamp 1
transform 1 0 105892 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1148
timestamp 1636968456
transform 1 0 106720 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1160
timestamp 1636968456
transform 1 0 107824 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1172
timestamp 1636968456
transform 1 0 108928 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1184
timestamp 1
transform 1 0 110032 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636968456
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636968456
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1636968456
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1636968456
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1636968456
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_69
timestamp 1
transform 1 0 7452 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1122
timestamp 1636968456
transform 1 0 104328 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1134
timestamp 1636968456
transform 1 0 105432 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1146
timestamp 1636968456
transform 1 0 106536 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1158
timestamp 1636968456
transform 1 0 107640 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_1170
timestamp 1
transform 1 0 108744 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_1174
timestamp 1
transform 1 0 109112 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1176
timestamp 1636968456
transform 1 0 109296 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_1188
timestamp 1
transform 1 0 110400 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636968456
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636968456
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636968456
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1636968456
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1636968456
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_65
timestamp 1
transform 1 0 7084 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_78_1136
timestamp 1
transform 1 0 105616 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_1144
timestamp 1
transform 1 0 106352 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1148
timestamp 1636968456
transform 1 0 106720 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1160
timestamp 1636968456
transform 1 0 107824 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1172
timestamp 1636968456
transform 1 0 108928 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_1184
timestamp 1
transform 1 0 110032 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636968456
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636968456
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636968456
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1636968456
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1636968456
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_69
timestamp 1
transform 1 0 7452 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1122
timestamp 1636968456
transform 1 0 104328 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1134
timestamp 1636968456
transform 1 0 105432 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1146
timestamp 1636968456
transform 1 0 106536 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1158
timestamp 1636968456
transform 1 0 107640 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_1170
timestamp 1
transform 1 0 108744 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_1174
timestamp 1
transform 1 0 109112 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1176
timestamp 1636968456
transform 1 0 109296 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_1188
timestamp 1
transform 1 0 110400 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636968456
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636968456
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636968456
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1636968456
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1636968456
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_65
timestamp 1
transform 1 0 7084 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1132
timestamp 1636968456
transform 1 0 105248 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_1144
timestamp 1
transform 1 0 106352 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1148
timestamp 1636968456
transform 1 0 106720 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1160
timestamp 1636968456
transform 1 0 107824 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1172
timestamp 1636968456
transform 1 0 108928 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_1184
timestamp 1
transform 1 0 110032 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636968456
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636968456
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1636968456
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1636968456
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1636968456
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_69
timestamp 1
transform 1 0 7452 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1122
timestamp 1636968456
transform 1 0 104328 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1134
timestamp 1636968456
transform 1 0 105432 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1146
timestamp 1636968456
transform 1 0 106536 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1158
timestamp 1636968456
transform 1 0 107640 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_1170
timestamp 1
transform 1 0 108744 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_1174
timestamp 1
transform 1 0 109112 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1176
timestamp 1636968456
transform 1 0 109296 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_1188
timestamp 1
transform 1 0 110400 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636968456
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636968456
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636968456
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1636968456
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1636968456
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_65
timestamp 1
transform 1 0 7084 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1122
timestamp 1636968456
transform 1 0 104328 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1134
timestamp 1636968456
transform 1 0 105432 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1146
timestamp 1
transform 1 0 106536 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1148
timestamp 1636968456
transform 1 0 106720 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1160
timestamp 1636968456
transform 1 0 107824 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1172
timestamp 1636968456
transform 1 0 108928 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_1184
timestamp 1
transform 1 0 110032 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636968456
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636968456
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636968456
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1636968456
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1636968456
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_69
timestamp 1
transform 1 0 7452 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1122
timestamp 1636968456
transform 1 0 104328 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1134
timestamp 1636968456
transform 1 0 105432 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1146
timestamp 1636968456
transform 1 0 106536 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1158
timestamp 1636968456
transform 1 0 107640 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_1170
timestamp 1
transform 1 0 108744 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_1174
timestamp 1
transform 1 0 109112 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1176
timestamp 1636968456
transform 1 0 109296 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_1188
timestamp 1
transform 1 0 110400 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636968456
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636968456
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636968456
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1636968456
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1636968456
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_65
timestamp 1
transform 1 0 7084 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1122
timestamp 1636968456
transform 1 0 104328 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1134
timestamp 1636968456
transform 1 0 105432 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_1146
timestamp 1
transform 1 0 106536 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1148
timestamp 1636968456
transform 1 0 106720 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1160
timestamp 1636968456
transform 1 0 107824 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1172
timestamp 1636968456
transform 1 0 108928 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_1184
timestamp 1
transform 1 0 110032 0 1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1636968456
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1636968456
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1636968456
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1636968456
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1636968456
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_69
timestamp 1
transform 1 0 7452 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1122
timestamp 1636968456
transform 1 0 104328 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1134
timestamp 1636968456
transform 1 0 105432 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1146
timestamp 1636968456
transform 1 0 106536 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1158
timestamp 1636968456
transform 1 0 107640 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_1170
timestamp 1
transform 1 0 108744 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_1174
timestamp 1
transform 1 0 109112 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1176
timestamp 1636968456
transform 1 0 109296 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_1188
timestamp 1
transform 1 0 110400 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636968456
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636968456
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636968456
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1636968456
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1636968456
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_65
timestamp 1
transform 1 0 7084 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1122
timestamp 1636968456
transform 1 0 104328 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1134
timestamp 1636968456
transform 1 0 105432 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_1146
timestamp 1
transform 1 0 106536 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1148
timestamp 1636968456
transform 1 0 106720 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1160
timestamp 1636968456
transform 1 0 107824 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1172
timestamp 1636968456
transform 1 0 108928 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_1184
timestamp 1
transform 1 0 110032 0 1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636968456
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636968456
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1636968456
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1636968456
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1636968456
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_69
timestamp 1
transform 1 0 7452 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1122
timestamp 1636968456
transform 1 0 104328 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1134
timestamp 1636968456
transform 1 0 105432 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1146
timestamp 1636968456
transform 1 0 106536 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1158
timestamp 1636968456
transform 1 0 107640 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_1170
timestamp 1
transform 1 0 108744 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_1174
timestamp 1
transform 1 0 109112 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1176
timestamp 1636968456
transform 1 0 109296 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_1188
timestamp 1
transform 1 0 110400 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636968456
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636968456
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636968456
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1636968456
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1636968456
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_65
timestamp 1
transform 1 0 7084 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1122
timestamp 1636968456
transform 1 0 104328 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1134
timestamp 1636968456
transform 1 0 105432 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_1146
timestamp 1
transform 1 0 106536 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1148
timestamp 1636968456
transform 1 0 106720 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1160
timestamp 1636968456
transform 1 0 107824 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1172
timestamp 1636968456
transform 1 0 108928 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_1184
timestamp 1
transform 1 0 110032 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636968456
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636968456
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1636968456
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1636968456
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1636968456
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_69
timestamp 1
transform 1 0 7452 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1122
timestamp 1636968456
transform 1 0 104328 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1134
timestamp 1636968456
transform 1 0 105432 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1146
timestamp 1636968456
transform 1 0 106536 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1158
timestamp 1636968456
transform 1 0 107640 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_1170
timestamp 1
transform 1 0 108744 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_1174
timestamp 1
transform 1 0 109112 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1176
timestamp 1636968456
transform 1 0 109296 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_1188
timestamp 1
transform 1 0 110400 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1636968456
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1636968456
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636968456
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1636968456
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1636968456
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_65
timestamp 1
transform 1 0 7084 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1122
timestamp 1636968456
transform 1 0 104328 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1134
timestamp 1636968456
transform 1 0 105432 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_1146
timestamp 1
transform 1 0 106536 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1148
timestamp 1636968456
transform 1 0 106720 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1160
timestamp 1636968456
transform 1 0 107824 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1172
timestamp 1636968456
transform 1 0 108928 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_1184
timestamp 1
transform 1 0 110032 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636968456
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636968456
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1636968456
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1636968456
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1636968456
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_69
timestamp 1
transform 1 0 7452 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1122
timestamp 1636968456
transform 1 0 104328 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1134
timestamp 1636968456
transform 1 0 105432 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1146
timestamp 1636968456
transform 1 0 106536 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1158
timestamp 1636968456
transform 1 0 107640 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_1170
timestamp 1
transform 1 0 108744 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_1174
timestamp 1
transform 1 0 109112 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1176
timestamp 1636968456
transform 1 0 109296 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_1188
timestamp 1
transform 1 0 110400 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1636968456
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1636968456
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636968456
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1636968456
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1636968456
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_65
timestamp 1
transform 1 0 7084 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1122
timestamp 1636968456
transform 1 0 104328 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1134
timestamp 1636968456
transform 1 0 105432 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_1146
timestamp 1
transform 1 0 106536 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1148
timestamp 1636968456
transform 1 0 106720 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1160
timestamp 1636968456
transform 1 0 107824 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1172
timestamp 1636968456
transform 1 0 108928 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_1184
timestamp 1
transform 1 0 110032 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636968456
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636968456
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636968456
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1636968456
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1636968456
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_69
timestamp 1
transform 1 0 7452 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1122
timestamp 1636968456
transform 1 0 104328 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1134
timestamp 1636968456
transform 1 0 105432 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1146
timestamp 1636968456
transform 1 0 106536 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1158
timestamp 1636968456
transform 1 0 107640 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_1170
timestamp 1
transform 1 0 108744 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_1174
timestamp 1
transform 1 0 109112 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1176
timestamp 1636968456
transform 1 0 109296 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_1188
timestamp 1
transform 1 0 110400 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636968456
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636968456
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636968456
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1636968456
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1636968456
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_65
timestamp 1
transform 1 0 7084 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1133
timestamp 1636968456
transform 1 0 105340 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_1145
timestamp 1
transform 1 0 106444 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1148
timestamp 1636968456
transform 1 0 106720 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1160
timestamp 1636968456
transform 1 0 107824 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1172
timestamp 1636968456
transform 1 0 108928 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_1184
timestamp 1
transform 1 0 110032 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1636968456
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1636968456
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1636968456
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1636968456
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1636968456
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_69
timestamp 1
transform 1 0 7452 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1127
timestamp 1636968456
transform 1 0 104788 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1139
timestamp 1636968456
transform 1 0 105892 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1151
timestamp 1636968456
transform 1 0 106996 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1163
timestamp 1636968456
transform 1 0 108100 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1176
timestamp 1636968456
transform 1 0 109296 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_1188
timestamp 1
transform 1 0 110400 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636968456
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636968456
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636968456
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1636968456
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1636968456
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_65
timestamp 1
transform 1 0 7084 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1150
timestamp 1636968456
transform 1 0 106904 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1162
timestamp 1636968456
transform 1 0 108008 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1174
timestamp 1636968456
transform 1 0 109112 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_1186
timestamp 1
transform 1 0 110216 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636968456
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636968456
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1636968456
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1636968456
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1636968456
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_69
timestamp 1
transform 1 0 7452 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1122
timestamp 1636968456
transform 1 0 104328 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1134
timestamp 1636968456
transform 1 0 105432 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1146
timestamp 1636968456
transform 1 0 106536 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1158
timestamp 1636968456
transform 1 0 107640 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_1170
timestamp 1
transform 1 0 108744 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_1174
timestamp 1
transform 1 0 109112 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1176
timestamp 1636968456
transform 1 0 109296 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_1188
timestamp 1
transform 1 0 110400 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636968456
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636968456
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636968456
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1636968456
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1636968456
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_65
timestamp 1
transform 1 0 7084 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1125
timestamp 1636968456
transform 1 0 104604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_1137
timestamp 1
transform 1 0 105708 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_1145
timestamp 1
transform 1 0 106444 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1148
timestamp 1636968456
transform 1 0 106720 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1160
timestamp 1636968456
transform 1 0 107824 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1172
timestamp 1636968456
transform 1 0 108928 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_1184
timestamp 1
transform 1 0 110032 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636968456
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636968456
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1636968456
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1636968456
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1636968456
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_69
timestamp 1
transform 1 0 7452 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1122
timestamp 1636968456
transform 1 0 104328 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1134
timestamp 1636968456
transform 1 0 105432 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1146
timestamp 1636968456
transform 1 0 106536 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1158
timestamp 1636968456
transform 1 0 107640 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_1170
timestamp 1
transform 1 0 108744 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_1174
timestamp 1
transform 1 0 109112 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1176
timestamp 1636968456
transform 1 0 109296 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_1188
timestamp 1
transform 1 0 110400 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1636968456
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1636968456
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1636968456
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1636968456
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1636968456
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_65
timestamp 1
transform 1 0 7084 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_1122
timestamp 1
transform 1 0 104328 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1133
timestamp 1636968456
transform 1 0 105340 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_1145
timestamp 1
transform 1 0 106444 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1148
timestamp 1636968456
transform 1 0 106720 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1160
timestamp 1636968456
transform 1 0 107824 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1172
timestamp 1636968456
transform 1 0 108928 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_1184
timestamp 1
transform 1 0 110032 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636968456
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636968456
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_27
timestamp 1636968456
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1636968456
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1636968456
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_69
timestamp 1
transform 1 0 7452 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1149
timestamp 1636968456
transform 1 0 106812 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1161
timestamp 1636968456
transform 1 0 107916 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_1173
timestamp 1
transform 1 0 109020 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1176
timestamp 1636968456
transform 1 0 109296 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_1188
timestamp 1
transform 1 0 110400 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1636968456
transform 1 0 1380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1636968456
transform 1 0 2484 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1636968456
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1636968456
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1636968456
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_65
timestamp 1
transform 1 0 7084 0 1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1124
timestamp 1636968456
transform 1 0 104512 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_1136
timestamp 1
transform 1 0 105616 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_102_1144
timestamp 1
transform 1 0 106352 0 1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1148
timestamp 1636968456
transform 1 0 106720 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1160
timestamp 1636968456
transform 1 0 107824 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1172
timestamp 1636968456
transform 1 0 108928 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_1184
timestamp 1
transform 1 0 110032 0 1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636968456
transform 1 0 1380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636968456
transform 1 0 2484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1636968456
transform 1 0 3588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_39
timestamp 1636968456
transform 1 0 4692 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1
transform 1 0 5796 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1636968456
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_69
timestamp 1
transform 1 0 7452 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1122
timestamp 1636968456
transform 1 0 104328 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1134
timestamp 1636968456
transform 1 0 105432 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1146
timestamp 1636968456
transform 1 0 106536 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1158
timestamp 1636968456
transform 1 0 107640 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_1170
timestamp 1
transform 1 0 108744 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_1174
timestamp 1
transform 1 0 109112 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1176
timestamp 1636968456
transform 1 0 109296 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_1188
timestamp 1
transform 1 0 110400 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1636968456
transform 1 0 1380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1636968456
transform 1 0 2484 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1636968456
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1636968456
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1636968456
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_65
timestamp 1
transform 1 0 7084 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1122
timestamp 1636968456
transform 1 0 104328 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1134
timestamp 1636968456
transform 1 0 105432 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_1146
timestamp 1
transform 1 0 106536 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1148
timestamp 1636968456
transform 1 0 106720 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1160
timestamp 1636968456
transform 1 0 107824 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1172
timestamp 1636968456
transform 1 0 108928 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_1184
timestamp 1
transform 1 0 110032 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_105_3
timestamp 1636968456
transform 1 0 1380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_15
timestamp 1636968456
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_27
timestamp 1636968456
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_39
timestamp 1636968456
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1636968456
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_69
timestamp 1
transform 1 0 7452 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1122
timestamp 1636968456
transform 1 0 104328 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1134
timestamp 1636968456
transform 1 0 105432 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1146
timestamp 1636968456
transform 1 0 106536 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1158
timestamp 1636968456
transform 1 0 107640 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_1170
timestamp 1
transform 1 0 108744 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_1174
timestamp 1
transform 1 0 109112 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1176
timestamp 1636968456
transform 1 0 109296 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_105_1188
timestamp 1
transform 1 0 110400 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636968456
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636968456
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636968456
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1636968456
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1636968456
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_65
timestamp 1
transform 1 0 7084 0 1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1125
timestamp 1636968456
transform 1 0 104604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_1137
timestamp 1
transform 1 0 105708 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_1145
timestamp 1
transform 1 0 106444 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1148
timestamp 1636968456
transform 1 0 106720 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1160
timestamp 1636968456
transform 1 0 107824 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1172
timestamp 1636968456
transform 1 0 108928 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_1184
timestamp 1
transform 1 0 110032 0 1 59840
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636968456
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636968456
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1636968456
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_39
timestamp 1636968456
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1636968456
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_69
timestamp 1
transform 1 0 7452 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1122
timestamp 1636968456
transform 1 0 104328 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1134
timestamp 1636968456
transform 1 0 105432 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1146
timestamp 1636968456
transform 1 0 106536 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1158
timestamp 1636968456
transform 1 0 107640 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_1170
timestamp 1
transform 1 0 108744 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_1174
timestamp 1
transform 1 0 109112 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1176
timestamp 1636968456
transform 1 0 109296 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_1188
timestamp 1
transform 1 0 110400 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636968456
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636968456
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636968456
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1636968456
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1636968456
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_65
timestamp 1
transform 1 0 7084 0 1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1122
timestamp 1636968456
transform 1 0 104328 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1134
timestamp 1636968456
transform 1 0 105432 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_1146
timestamp 1
transform 1 0 106536 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1148
timestamp 1636968456
transform 1 0 106720 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1160
timestamp 1636968456
transform 1 0 107824 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1172
timestamp 1636968456
transform 1 0 108928 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_1184
timestamp 1
transform 1 0 110032 0 1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1636968456
transform 1 0 1380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1636968456
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_27
timestamp 1636968456
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_39
timestamp 1636968456
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1636968456
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_69
timestamp 1
transform 1 0 7452 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1122
timestamp 1636968456
transform 1 0 104328 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1134
timestamp 1636968456
transform 1 0 105432 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1146
timestamp 1636968456
transform 1 0 106536 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1158
timestamp 1636968456
transform 1 0 107640 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_1170
timestamp 1
transform 1 0 108744 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_1174
timestamp 1
transform 1 0 109112 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1176
timestamp 1636968456
transform 1 0 109296 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_1188
timestamp 1
transform 1 0 110400 0 -1 62016
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_110_3
timestamp 1636968456
transform 1 0 1380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_15
timestamp 1636968456
transform 1 0 2484 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636968456
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1636968456
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1636968456
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_65
timestamp 1
transform 1 0 7084 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1122
timestamp 1636968456
transform 1 0 104328 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1134
timestamp 1636968456
transform 1 0 105432 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_1146
timestamp 1
transform 1 0 106536 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1148
timestamp 1636968456
transform 1 0 106720 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1160
timestamp 1636968456
transform 1 0 107824 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1172
timestamp 1636968456
transform 1 0 108928 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_1184
timestamp 1
transform 1 0 110032 0 1 62016
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636968456
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636968456
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1636968456
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_39
timestamp 1636968456
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1636968456
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_69
timestamp 1
transform 1 0 7452 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1122
timestamp 1636968456
transform 1 0 104328 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1134
timestamp 1636968456
transform 1 0 105432 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1146
timestamp 1636968456
transform 1 0 106536 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1158
timestamp 1636968456
transform 1 0 107640 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_1170
timestamp 1
transform 1 0 108744 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_1174
timestamp 1
transform 1 0 109112 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1176
timestamp 1636968456
transform 1 0 109296 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_1188
timestamp 1
transform 1 0 110400 0 -1 63104
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1636968456
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1636968456
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636968456
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1636968456
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1636968456
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_65
timestamp 1
transform 1 0 7084 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1122
timestamp 1636968456
transform 1 0 104328 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1134
timestamp 1636968456
transform 1 0 105432 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_1146
timestamp 1
transform 1 0 106536 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1148
timestamp 1636968456
transform 1 0 106720 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1160
timestamp 1636968456
transform 1 0 107824 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1172
timestamp 1636968456
transform 1 0 108928 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_1184
timestamp 1
transform 1 0 110032 0 1 63104
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636968456
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636968456
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636968456
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1636968456
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1636968456
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_69
timestamp 1
transform 1 0 7452 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1122
timestamp 1636968456
transform 1 0 104328 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1134
timestamp 1636968456
transform 1 0 105432 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1146
timestamp 1636968456
transform 1 0 106536 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1158
timestamp 1636968456
transform 1 0 107640 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_1170
timestamp 1
transform 1 0 108744 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_1174
timestamp 1
transform 1 0 109112 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1176
timestamp 1636968456
transform 1 0 109296 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_1188
timestamp 1
transform 1 0 110400 0 -1 64192
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636968456
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636968456
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636968456
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1636968456
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1636968456
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_65
timestamp 1
transform 1 0 7084 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1122
timestamp 1636968456
transform 1 0 104328 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1134
timestamp 1636968456
transform 1 0 105432 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_1146
timestamp 1
transform 1 0 106536 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1148
timestamp 1636968456
transform 1 0 106720 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1160
timestamp 1636968456
transform 1 0 107824 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1172
timestamp 1636968456
transform 1 0 108928 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_1184
timestamp 1
transform 1 0 110032 0 1 64192
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_115_3
timestamp 1636968456
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_15
timestamp 1636968456
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_27
timestamp 1636968456
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_39
timestamp 1636968456
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1636968456
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_115_69
timestamp 1
transform 1 0 7452 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1122
timestamp 1636968456
transform 1 0 104328 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1134
timestamp 1636968456
transform 1 0 105432 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1146
timestamp 1636968456
transform 1 0 106536 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1158
timestamp 1636968456
transform 1 0 107640 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_1170
timestamp 1
transform 1 0 108744 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_1174
timestamp 1
transform 1 0 109112 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1176
timestamp 1636968456
transform 1 0 109296 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_115_1188
timestamp 1
transform 1 0 110400 0 -1 65280
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636968456
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636968456
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636968456
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1636968456
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_53
timestamp 1636968456
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_65
timestamp 1
transform 1 0 7084 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1122
timestamp 1636968456
transform 1 0 104328 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1134
timestamp 1636968456
transform 1 0 105432 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_1146
timestamp 1
transform 1 0 106536 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1148
timestamp 1636968456
transform 1 0 106720 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1160
timestamp 1636968456
transform 1 0 107824 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1172
timestamp 1636968456
transform 1 0 108928 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_1184
timestamp 1
transform 1 0 110032 0 1 65280
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636968456
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636968456
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_27
timestamp 1
transform 1 0 3588 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_29
timestamp 1636968456
transform 1 0 3772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_41
timestamp 1636968456
transform 1 0 4876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_53
timestamp 1
transform 1 0 5980 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1636968456
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1636968456
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_81
timestamp 1
transform 1 0 8556 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_85
timestamp 1636968456
transform 1 0 8924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_97
timestamp 1636968456
transform 1 0 10028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_109
timestamp 1
transform 1 0 11132 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1636968456
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_125
timestamp 1636968456
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_137
timestamp 1
transform 1 0 13708 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_141
timestamp 1636968456
transform 1 0 14076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_153
timestamp 1636968456
transform 1 0 15180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_165
timestamp 1
transform 1 0 16284 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_169
timestamp 1636968456
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_181
timestamp 1636968456
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_193
timestamp 1
transform 1 0 18860 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_197
timestamp 1636968456
transform 1 0 19228 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_209
timestamp 1636968456
transform 1 0 20332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_221
timestamp 1
transform 1 0 21436 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_225
timestamp 1636968456
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_237
timestamp 1636968456
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_249
timestamp 1
transform 1 0 24012 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_253
timestamp 1636968456
transform 1 0 24380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_265
timestamp 1636968456
transform 1 0 25484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_277
timestamp 1
transform 1 0 26588 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_281
timestamp 1636968456
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_293
timestamp 1636968456
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_305
timestamp 1
transform 1 0 29164 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_309
timestamp 1636968456
transform 1 0 29532 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_321
timestamp 1636968456
transform 1 0 30636 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_333
timestamp 1
transform 1 0 31740 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_337
timestamp 1636968456
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_349
timestamp 1636968456
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_361
timestamp 1
transform 1 0 34316 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_365
timestamp 1636968456
transform 1 0 34684 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_377
timestamp 1636968456
transform 1 0 35788 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_389
timestamp 1
transform 1 0 36892 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_393
timestamp 1636968456
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_405
timestamp 1636968456
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_417
timestamp 1
transform 1 0 39468 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_421
timestamp 1636968456
transform 1 0 39836 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_433
timestamp 1636968456
transform 1 0 40940 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_445
timestamp 1
transform 1 0 42044 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_449
timestamp 1636968456
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_461
timestamp 1636968456
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_473
timestamp 1
transform 1 0 44620 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_477
timestamp 1636968456
transform 1 0 44988 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_489
timestamp 1636968456
transform 1 0 46092 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_501
timestamp 1
transform 1 0 47196 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_117_505
timestamp 1
transform 1 0 47564 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_513
timestamp 1
transform 1 0 48300 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_519
timestamp 1636968456
transform 1 0 48852 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_531
timestamp 1
transform 1 0 49956 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_117_533
timestamp 1
transform 1 0 50140 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_539
timestamp 1636968456
transform 1 0 50692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_551
timestamp 1
transform 1 0 51796 0 -1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_561
timestamp 1636968456
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_573
timestamp 1
transform 1 0 53820 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_577
timestamp 1
transform 1 0 54188 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_585
timestamp 1
transform 1 0 54924 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_117_589
timestamp 1
transform 1 0 55292 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_117_595
timestamp 1
transform 1 0 55844 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_624
timestamp 1
transform 1 0 58512 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_631
timestamp 1636968456
transform 1 0 59156 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_643
timestamp 1
transform 1 0 60260 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_117_645
timestamp 1
transform 1 0 60444 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_117_651
timestamp 1
transform 1 0 60996 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_117_680
timestamp 1
transform 1 0 63664 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_117_697
timestamp 1
transform 1 0 65228 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_117_701
timestamp 1
transform 1 0 65596 0 -1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_710
timestamp 1636968456
transform 1 0 66424 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_722
timestamp 1
transform 1 0 67528 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_729
timestamp 1636968456
transform 1 0 68172 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_741
timestamp 1
transform 1 0 69276 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_117_746
timestamp 1
transform 1 0 69736 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_754
timestamp 1
transform 1 0 70472 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_117_757
timestamp 1
transform 1 0 70748 0 -1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_766
timestamp 1636968456
transform 1 0 71576 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_778
timestamp 1
transform 1 0 72680 0 -1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_788
timestamp 1636968456
transform 1 0 73600 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_800
timestamp 1
transform 1 0 74704 0 -1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_818
timestamp 1636968456
transform 1 0 76360 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_830
timestamp 1
transform 1 0 77464 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_838
timestamp 1
transform 1 0 78200 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_841
timestamp 1636968456
transform 1 0 78476 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_853
timestamp 1636968456
transform 1 0 79580 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_865
timestamp 1
transform 1 0 80684 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_869
timestamp 1636968456
transform 1 0 81052 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_881
timestamp 1636968456
transform 1 0 82156 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_893
timestamp 1
transform 1 0 83260 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_897
timestamp 1636968456
transform 1 0 83628 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_909
timestamp 1636968456
transform 1 0 84732 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_921
timestamp 1
transform 1 0 85836 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_117_927
timestamp 1
transform 1 0 86388 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_935
timestamp 1
transform 1 0 87124 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_939
timestamp 1636968456
transform 1 0 87492 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_951
timestamp 1
transform 1 0 88596 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_953
timestamp 1636968456
transform 1 0 88780 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_965
timestamp 1636968456
transform 1 0 89884 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_977
timestamp 1
transform 1 0 90988 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_117_981
timestamp 1
transform 1 0 91356 0 -1 66368
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_117_994
timestamp 1636968456
transform 1 0 92552 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_117_1006
timestamp 1
transform 1 0 93656 0 -1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1009
timestamp 1636968456
transform 1 0 93932 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_1021
timestamp 1
transform 1 0 95036 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1029
timestamp 1
transform 1 0 95772 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_117_1032
timestamp 1
transform 1 0 96048 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1037
timestamp 1636968456
transform 1 0 96508 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1049
timestamp 1636968456
transform 1 0 97612 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1061
timestamp 1
transform 1 0 98716 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1065
timestamp 1636968456
transform 1 0 99084 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1077
timestamp 1636968456
transform 1 0 100188 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1089
timestamp 1
transform 1 0 101292 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1093
timestamp 1636968456
transform 1 0 101660 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1105
timestamp 1636968456
transform 1 0 102764 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1117
timestamp 1
transform 1 0 103868 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1121
timestamp 1636968456
transform 1 0 104236 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1133
timestamp 1636968456
transform 1 0 105340 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1145
timestamp 1
transform 1 0 106444 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1149
timestamp 1636968456
transform 1 0 106812 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1161
timestamp 1636968456
transform 1 0 107916 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_1173
timestamp 1
transform 1 0 109020 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1177
timestamp 1636968456
transform 1 0 109388 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1189
timestamp 1
transform 1 0 110492 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636968456
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636968456
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636968456
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1636968456
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1636968456
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1636968456
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1636968456
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1636968456
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1636968456
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1636968456
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1636968456
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1636968456
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_165
timestamp 1636968456
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_177
timestamp 1636968456
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_197
timestamp 1636968456
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_209
timestamp 1636968456
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_221
timestamp 1636968456
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_233
timestamp 1636968456
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_253
timestamp 1636968456
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_265
timestamp 1636968456
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_277
timestamp 1636968456
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_289
timestamp 1636968456
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_309
timestamp 1636968456
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_321
timestamp 1636968456
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_333
timestamp 1636968456
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_345
timestamp 1636968456
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_365
timestamp 1636968456
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_377
timestamp 1636968456
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_389
timestamp 1636968456
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_401
timestamp 1636968456
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_421
timestamp 1636968456
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_433
timestamp 1636968456
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_445
timestamp 1636968456
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_457
timestamp 1636968456
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_477
timestamp 1636968456
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_489
timestamp 1636968456
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_501
timestamp 1
transform 1 0 47196 0 1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_507
timestamp 1636968456
transform 1 0 47748 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_519
timestamp 1
transform 1 0 48852 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_529
timestamp 1
transform 1 0 49772 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_533
timestamp 1636968456
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_545
timestamp 1
transform 1 0 51244 0 1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_571
timestamp 1636968456
transform 1 0 53636 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_583
timestamp 1
transform 1 0 54740 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_118_589
timestamp 1
transform 1 0 55292 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_592
timestamp 1636968456
transform 1 0 55568 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_604
timestamp 1636968456
transform 1 0 56672 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_616
timestamp 1636968456
transform 1 0 57776 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_628
timestamp 1
transform 1 0 58880 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_634
timestamp 1
transform 1 0 59432 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_645
timestamp 1
transform 1 0 60444 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_118_675
timestamp 1636968456
transform 1 0 63204 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_687
timestamp 1636968456
transform 1 0 64308 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_703
timestamp 1636968456
transform 1 0 65780 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_715
timestamp 1636968456
transform 1 0 66884 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_727
timestamp 1636968456
transform 1 0 67988 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_739
timestamp 1
transform 1 0 69092 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_118_749
timestamp 1
transform 1 0 70012 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_755
timestamp 1
transform 1 0 70564 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_757
timestamp 1
transform 1 0 70748 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_118_765
timestamp 1
transform 1 0 71484 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_790
timestamp 1636968456
transform 1 0 73784 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_802
timestamp 1
transform 1 0 74888 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_118_810
timestamp 1
transform 1 0 75624 0 1 66368
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_118_813
timestamp 1636968456
transform 1 0 75900 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_825
timestamp 1636968456
transform 1 0 77004 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_837
timestamp 1636968456
transform 1 0 78108 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_849
timestamp 1636968456
transform 1 0 79212 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_861
timestamp 1
transform 1 0 80316 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_867
timestamp 1
transform 1 0 80868 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_869
timestamp 1636968456
transform 1 0 81052 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_881
timestamp 1636968456
transform 1 0 82156 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_893
timestamp 1636968456
transform 1 0 83260 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_905
timestamp 1636968456
transform 1 0 84364 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_917
timestamp 1
transform 1 0 85468 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_923
timestamp 1
transform 1 0 86020 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_925
timestamp 1636968456
transform 1 0 86204 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_937
timestamp 1636968456
transform 1 0 87308 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_949
timestamp 1636968456
transform 1 0 88412 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_961
timestamp 1636968456
transform 1 0 89516 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_973
timestamp 1
transform 1 0 90620 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_979
timestamp 1
transform 1 0 91172 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_981
timestamp 1636968456
transform 1 0 91356 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_993
timestamp 1636968456
transform 1 0 92460 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1005
timestamp 1636968456
transform 1 0 93564 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1017
timestamp 1636968456
transform 1 0 94668 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1029
timestamp 1
transform 1 0 95772 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1035
timestamp 1
transform 1 0 96324 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1037
timestamp 1636968456
transform 1 0 96508 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1049
timestamp 1636968456
transform 1 0 97612 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1061
timestamp 1636968456
transform 1 0 98716 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1073
timestamp 1636968456
transform 1 0 99820 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1085
timestamp 1
transform 1 0 100924 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1091
timestamp 1
transform 1 0 101476 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1093
timestamp 1636968456
transform 1 0 101660 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1105
timestamp 1636968456
transform 1 0 102764 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1117
timestamp 1636968456
transform 1 0 103868 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1129
timestamp 1636968456
transform 1 0 104972 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1141
timestamp 1
transform 1 0 106076 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1147
timestamp 1
transform 1 0 106628 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1149
timestamp 1636968456
transform 1 0 106812 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1161
timestamp 1636968456
transform 1 0 107916 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1173
timestamp 1636968456
transform 1 0 109020 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_1185
timestamp 1
transform 1 0 110124 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1189
timestamp 1
transform 1 0 110492 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636968456
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636968456
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1636968456
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_39
timestamp 1636968456
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1636968456
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_69
timestamp 1636968456
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_81
timestamp 1636968456
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_93
timestamp 1636968456
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1636968456
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1636968456
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1636968456
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1636968456
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_169
timestamp 1636968456
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_181
timestamp 1636968456
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_193
timestamp 1636968456
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_205
timestamp 1636968456
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_225
timestamp 1636968456
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_237
timestamp 1636968456
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_249
timestamp 1636968456
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_261
timestamp 1636968456
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_281
timestamp 1636968456
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_293
timestamp 1636968456
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_305
timestamp 1636968456
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_317
timestamp 1636968456
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_337
timestamp 1636968456
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_349
timestamp 1636968456
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_361
timestamp 1636968456
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_373
timestamp 1636968456
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_393
timestamp 1636968456
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_405
timestamp 1636968456
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_417
timestamp 1636968456
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_429
timestamp 1636968456
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_449
timestamp 1
transform 1 0 42412 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_119_527
timestamp 1
transform 1 0 49588 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_119_552
timestamp 1
transform 1 0 51888 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_119_561
timestamp 1
transform 1 0 52716 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_569
timestamp 1
transform 1 0 53452 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_119_612
timestamp 1
transform 1 0 57408 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_657
timestamp 1636968456
transform 1 0 61548 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_669
timestamp 1
transform 1 0 62652 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_673
timestamp 1
transform 1 0 63020 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_677
timestamp 1
transform 1 0 63388 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_119_700
timestamp 1
transform 1 0 65504 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_721
timestamp 1
transform 1 0 67436 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_725
timestamp 1
transform 1 0 67804 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_769
timestamp 1636968456
transform 1 0 71852 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_781
timestamp 1
transform 1 0 72956 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_119_785
timestamp 1
transform 1 0 73324 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_793
timestamp 1
transform 1 0 74060 0 -1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_818
timestamp 1636968456
transform 1 0 76360 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_830
timestamp 1
transform 1 0 77464 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_119_838
timestamp 1
transform 1 0 78200 0 -1 67456
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_841
timestamp 1636968456
transform 1 0 78476 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_853
timestamp 1636968456
transform 1 0 79580 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_865
timestamp 1636968456
transform 1 0 80684 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_877
timestamp 1636968456
transform 1 0 81788 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_889
timestamp 1
transform 1 0 82892 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_895
timestamp 1
transform 1 0 83444 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_897
timestamp 1636968456
transform 1 0 83628 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_909
timestamp 1636968456
transform 1 0 84732 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_921
timestamp 1636968456
transform 1 0 85836 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_933
timestamp 1636968456
transform 1 0 86940 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_945
timestamp 1
transform 1 0 88044 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_951
timestamp 1
transform 1 0 88596 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_953
timestamp 1636968456
transform 1 0 88780 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_965
timestamp 1636968456
transform 1 0 89884 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_977
timestamp 1636968456
transform 1 0 90988 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_989
timestamp 1636968456
transform 1 0 92092 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1001
timestamp 1
transform 1 0 93196 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1007
timestamp 1
transform 1 0 93748 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1009
timestamp 1636968456
transform 1 0 93932 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1021
timestamp 1636968456
transform 1 0 95036 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1033
timestamp 1636968456
transform 1 0 96140 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1045
timestamp 1636968456
transform 1 0 97244 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1057
timestamp 1
transform 1 0 98348 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1063
timestamp 1
transform 1 0 98900 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1065
timestamp 1636968456
transform 1 0 99084 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1077
timestamp 1636968456
transform 1 0 100188 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1089
timestamp 1636968456
transform 1 0 101292 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1101
timestamp 1636968456
transform 1 0 102396 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1113
timestamp 1
transform 1 0 103500 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1119
timestamp 1
transform 1 0 104052 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1121
timestamp 1636968456
transform 1 0 104236 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1133
timestamp 1636968456
transform 1 0 105340 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1145
timestamp 1636968456
transform 1 0 106444 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1157
timestamp 1636968456
transform 1 0 107548 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1169
timestamp 1
transform 1 0 108652 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1175
timestamp 1
transform 1 0 109204 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1177
timestamp 1636968456
transform 1 0 109388 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1189
timestamp 1
transform 1 0 110492 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1636968456
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1636968456
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636968456
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1636968456
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1636968456
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_65
timestamp 1636968456
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1636968456
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1636968456
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_109
timestamp 1636968456
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_121
timestamp 1636968456
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1636968456
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_153
timestamp 1636968456
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_165
timestamp 1636968456
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_177
timestamp 1636968456
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_197
timestamp 1636968456
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_209
timestamp 1636968456
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_221
timestamp 1636968456
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_233
timestamp 1636968456
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_253
timestamp 1636968456
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_265
timestamp 1636968456
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_277
timestamp 1636968456
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_289
timestamp 1636968456
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_309
timestamp 1636968456
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_321
timestamp 1636968456
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_333
timestamp 1636968456
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_345
timestamp 1636968456
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_365
timestamp 1636968456
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_377
timestamp 1636968456
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_389
timestamp 1636968456
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_401
timestamp 1636968456
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_421
timestamp 1636968456
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_433
timestamp 1636968456
transform 1 0 40940 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_445
timestamp 1636968456
transform 1 0 42044 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_457
timestamp 1636968456
transform 1 0 43148 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1
transform 1 0 44252 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1
transform 1 0 44804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_477
timestamp 1636968456
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_489
timestamp 1636968456
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_501
timestamp 1636968456
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_513
timestamp 1636968456
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_533
timestamp 1636968456
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_545
timestamp 1636968456
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_557
timestamp 1636968456
transform 1 0 52348 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_569
timestamp 1636968456
transform 1 0 53452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1
transform 1 0 54556 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1
transform 1 0 55108 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_589
timestamp 1636968456
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_601
timestamp 1636968456
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_613
timestamp 1636968456
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_625
timestamp 1636968456
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_645
timestamp 1636968456
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_657
timestamp 1636968456
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_669
timestamp 1636968456
transform 1 0 62652 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_681
timestamp 1636968456
transform 1 0 63756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1
transform 1 0 64860 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_701
timestamp 1636968456
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_713
timestamp 1636968456
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_725
timestamp 1636968456
transform 1 0 67804 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_737
timestamp 1636968456
transform 1 0 68908 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_749
timestamp 1
transform 1 0 70012 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_755
timestamp 1
transform 1 0 70564 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_757
timestamp 1636968456
transform 1 0 70748 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_769
timestamp 1636968456
transform 1 0 71852 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_781
timestamp 1636968456
transform 1 0 72956 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_793
timestamp 1636968456
transform 1 0 74060 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_805
timestamp 1
transform 1 0 75164 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_811
timestamp 1
transform 1 0 75716 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_813
timestamp 1636968456
transform 1 0 75900 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_825
timestamp 1636968456
transform 1 0 77004 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_837
timestamp 1636968456
transform 1 0 78108 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_849
timestamp 1636968456
transform 1 0 79212 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_861
timestamp 1
transform 1 0 80316 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_867
timestamp 1
transform 1 0 80868 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_869
timestamp 1636968456
transform 1 0 81052 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_881
timestamp 1636968456
transform 1 0 82156 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_893
timestamp 1636968456
transform 1 0 83260 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_905
timestamp 1636968456
transform 1 0 84364 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_917
timestamp 1
transform 1 0 85468 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_923
timestamp 1
transform 1 0 86020 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_925
timestamp 1636968456
transform 1 0 86204 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_937
timestamp 1636968456
transform 1 0 87308 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_949
timestamp 1636968456
transform 1 0 88412 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_961
timestamp 1636968456
transform 1 0 89516 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_973
timestamp 1
transform 1 0 90620 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_979
timestamp 1
transform 1 0 91172 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_981
timestamp 1636968456
transform 1 0 91356 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_993
timestamp 1636968456
transform 1 0 92460 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1005
timestamp 1636968456
transform 1 0 93564 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1017
timestamp 1636968456
transform 1 0 94668 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1029
timestamp 1
transform 1 0 95772 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1035
timestamp 1
transform 1 0 96324 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1037
timestamp 1636968456
transform 1 0 96508 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1049
timestamp 1636968456
transform 1 0 97612 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1061
timestamp 1636968456
transform 1 0 98716 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1073
timestamp 1636968456
transform 1 0 99820 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1085
timestamp 1
transform 1 0 100924 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1091
timestamp 1
transform 1 0 101476 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1093
timestamp 1636968456
transform 1 0 101660 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1105
timestamp 1636968456
transform 1 0 102764 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1117
timestamp 1636968456
transform 1 0 103868 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1129
timestamp 1636968456
transform 1 0 104972 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1141
timestamp 1
transform 1 0 106076 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1147
timestamp 1
transform 1 0 106628 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1149
timestamp 1636968456
transform 1 0 106812 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1161
timestamp 1636968456
transform 1 0 107916 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1173
timestamp 1636968456
transform 1 0 109020 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_1185
timestamp 1
transform 1 0 110124 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1189
timestamp 1
transform 1 0 110492 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636968456
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636968456
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1636968456
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_39
timestamp 1636968456
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1636968456
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_69
timestamp 1636968456
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_81
timestamp 1636968456
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_93
timestamp 1636968456
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_113
timestamp 1636968456
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_125
timestamp 1636968456
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_137
timestamp 1636968456
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_149
timestamp 1636968456
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_169
timestamp 1636968456
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_181
timestamp 1636968456
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_193
timestamp 1636968456
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_205
timestamp 1636968456
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_225
timestamp 1636968456
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_237
timestamp 1636968456
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_249
timestamp 1636968456
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_261
timestamp 1636968456
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_281
timestamp 1636968456
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_293
timestamp 1636968456
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_305
timestamp 1636968456
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_317
timestamp 1636968456
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_337
timestamp 1636968456
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_349
timestamp 1636968456
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_361
timestamp 1636968456
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_373
timestamp 1636968456
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_393
timestamp 1636968456
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_405
timestamp 1636968456
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_417
timestamp 1636968456
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_429
timestamp 1636968456
transform 1 0 40572 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_441
timestamp 1
transform 1 0 41676 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1
transform 1 0 42228 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_449
timestamp 1636968456
transform 1 0 42412 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_461
timestamp 1636968456
transform 1 0 43516 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_473
timestamp 1636968456
transform 1 0 44620 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_485
timestamp 1636968456
transform 1 0 45724 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1
transform 1 0 46828 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1
transform 1 0 47380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_505
timestamp 1636968456
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_517
timestamp 1636968456
transform 1 0 48668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_529
timestamp 1636968456
transform 1 0 49772 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_541
timestamp 1636968456
transform 1 0 50876 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_553
timestamp 1
transform 1 0 51980 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_559
timestamp 1
transform 1 0 52532 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_561
timestamp 1636968456
transform 1 0 52716 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_573
timestamp 1636968456
transform 1 0 53820 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_585
timestamp 1636968456
transform 1 0 54924 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_597
timestamp 1636968456
transform 1 0 56028 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_609
timestamp 1
transform 1 0 57132 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1
transform 1 0 57684 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_617
timestamp 1636968456
transform 1 0 57868 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_629
timestamp 1636968456
transform 1 0 58972 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_641
timestamp 1636968456
transform 1 0 60076 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_653
timestamp 1636968456
transform 1 0 61180 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_665
timestamp 1
transform 1 0 62284 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_671
timestamp 1
transform 1 0 62836 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_673
timestamp 1636968456
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_685
timestamp 1636968456
transform 1 0 64124 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_697
timestamp 1636968456
transform 1 0 65228 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_709
timestamp 1636968456
transform 1 0 66332 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_729
timestamp 1636968456
transform 1 0 68172 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_741
timestamp 1636968456
transform 1 0 69276 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_753
timestamp 1636968456
transform 1 0 70380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_765
timestamp 1636968456
transform 1 0 71484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_777
timestamp 1
transform 1 0 72588 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_783
timestamp 1
transform 1 0 73140 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_785
timestamp 1636968456
transform 1 0 73324 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_797
timestamp 1636968456
transform 1 0 74428 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_809
timestamp 1636968456
transform 1 0 75532 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_821
timestamp 1636968456
transform 1 0 76636 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_833
timestamp 1
transform 1 0 77740 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_839
timestamp 1
transform 1 0 78292 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_841
timestamp 1636968456
transform 1 0 78476 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_853
timestamp 1636968456
transform 1 0 79580 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_865
timestamp 1636968456
transform 1 0 80684 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_877
timestamp 1636968456
transform 1 0 81788 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_889
timestamp 1
transform 1 0 82892 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_895
timestamp 1
transform 1 0 83444 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_897
timestamp 1636968456
transform 1 0 83628 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_909
timestamp 1636968456
transform 1 0 84732 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_921
timestamp 1636968456
transform 1 0 85836 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_933
timestamp 1636968456
transform 1 0 86940 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_945
timestamp 1
transform 1 0 88044 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_951
timestamp 1
transform 1 0 88596 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_953
timestamp 1636968456
transform 1 0 88780 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_965
timestamp 1636968456
transform 1 0 89884 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_977
timestamp 1636968456
transform 1 0 90988 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_989
timestamp 1636968456
transform 1 0 92092 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1001
timestamp 1
transform 1 0 93196 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1007
timestamp 1
transform 1 0 93748 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1009
timestamp 1636968456
transform 1 0 93932 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1021
timestamp 1636968456
transform 1 0 95036 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1033
timestamp 1636968456
transform 1 0 96140 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1045
timestamp 1636968456
transform 1 0 97244 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1057
timestamp 1
transform 1 0 98348 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1063
timestamp 1
transform 1 0 98900 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1065
timestamp 1636968456
transform 1 0 99084 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1077
timestamp 1636968456
transform 1 0 100188 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1089
timestamp 1636968456
transform 1 0 101292 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1101
timestamp 1636968456
transform 1 0 102396 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1113
timestamp 1
transform 1 0 103500 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1119
timestamp 1
transform 1 0 104052 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1121
timestamp 1636968456
transform 1 0 104236 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1133
timestamp 1636968456
transform 1 0 105340 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1145
timestamp 1636968456
transform 1 0 106444 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1157
timestamp 1636968456
transform 1 0 107548 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1169
timestamp 1
transform 1 0 108652 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1175
timestamp 1
transform 1 0 109204 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1177
timestamp 1636968456
transform 1 0 109388 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1189
timestamp 1
transform 1 0 110492 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1636968456
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1636968456
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636968456
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1636968456
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1636968456
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_65
timestamp 1636968456
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_85
timestamp 1636968456
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_97
timestamp 1636968456
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_109
timestamp 1636968456
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_121
timestamp 1636968456
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_141
timestamp 1636968456
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_153
timestamp 1636968456
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_165
timestamp 1636968456
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_177
timestamp 1636968456
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_197
timestamp 1636968456
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_209
timestamp 1636968456
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_221
timestamp 1636968456
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_233
timestamp 1636968456
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_253
timestamp 1636968456
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_265
timestamp 1636968456
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_277
timestamp 1636968456
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_289
timestamp 1636968456
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_309
timestamp 1636968456
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_321
timestamp 1636968456
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_333
timestamp 1636968456
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_345
timestamp 1636968456
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_365
timestamp 1636968456
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_377
timestamp 1636968456
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_389
timestamp 1636968456
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_401
timestamp 1636968456
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_421
timestamp 1636968456
transform 1 0 39836 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_433
timestamp 1636968456
transform 1 0 40940 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_445
timestamp 1636968456
transform 1 0 42044 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_457
timestamp 1636968456
transform 1 0 43148 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_469
timestamp 1
transform 1 0 44252 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_475
timestamp 1
transform 1 0 44804 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_477
timestamp 1636968456
transform 1 0 44988 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_489
timestamp 1636968456
transform 1 0 46092 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_501
timestamp 1636968456
transform 1 0 47196 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_513
timestamp 1636968456
transform 1 0 48300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_525
timestamp 1
transform 1 0 49404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_531
timestamp 1
transform 1 0 49956 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_533
timestamp 1636968456
transform 1 0 50140 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_545
timestamp 1636968456
transform 1 0 51244 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_557
timestamp 1636968456
transform 1 0 52348 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_569
timestamp 1636968456
transform 1 0 53452 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_581
timestamp 1
transform 1 0 54556 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1
transform 1 0 55108 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_589
timestamp 1636968456
transform 1 0 55292 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_601
timestamp 1636968456
transform 1 0 56396 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_613
timestamp 1636968456
transform 1 0 57500 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_625
timestamp 1636968456
transform 1 0 58604 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_637
timestamp 1
transform 1 0 59708 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_643
timestamp 1
transform 1 0 60260 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_645
timestamp 1636968456
transform 1 0 60444 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_657
timestamp 1636968456
transform 1 0 61548 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_669
timestamp 1636968456
transform 1 0 62652 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_681
timestamp 1636968456
transform 1 0 63756 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_693
timestamp 1
transform 1 0 64860 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1
transform 1 0 65412 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_701
timestamp 1636968456
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_713
timestamp 1636968456
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_725
timestamp 1636968456
transform 1 0 67804 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_737
timestamp 1636968456
transform 1 0 68908 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_749
timestamp 1
transform 1 0 70012 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_755
timestamp 1
transform 1 0 70564 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_757
timestamp 1636968456
transform 1 0 70748 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_769
timestamp 1636968456
transform 1 0 71852 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_781
timestamp 1636968456
transform 1 0 72956 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_793
timestamp 1636968456
transform 1 0 74060 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_805
timestamp 1
transform 1 0 75164 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_811
timestamp 1
transform 1 0 75716 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_813
timestamp 1636968456
transform 1 0 75900 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_825
timestamp 1636968456
transform 1 0 77004 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_837
timestamp 1636968456
transform 1 0 78108 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_849
timestamp 1636968456
transform 1 0 79212 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_861
timestamp 1
transform 1 0 80316 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_867
timestamp 1
transform 1 0 80868 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_869
timestamp 1636968456
transform 1 0 81052 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_881
timestamp 1636968456
transform 1 0 82156 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_893
timestamp 1636968456
transform 1 0 83260 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_905
timestamp 1636968456
transform 1 0 84364 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_917
timestamp 1
transform 1 0 85468 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_923
timestamp 1
transform 1 0 86020 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_925
timestamp 1636968456
transform 1 0 86204 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_937
timestamp 1636968456
transform 1 0 87308 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_949
timestamp 1636968456
transform 1 0 88412 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_961
timestamp 1636968456
transform 1 0 89516 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_973
timestamp 1
transform 1 0 90620 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_979
timestamp 1
transform 1 0 91172 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_981
timestamp 1636968456
transform 1 0 91356 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_993
timestamp 1636968456
transform 1 0 92460 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1005
timestamp 1636968456
transform 1 0 93564 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1017
timestamp 1636968456
transform 1 0 94668 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1029
timestamp 1
transform 1 0 95772 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1035
timestamp 1
transform 1 0 96324 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1037
timestamp 1636968456
transform 1 0 96508 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1049
timestamp 1636968456
transform 1 0 97612 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1061
timestamp 1636968456
transform 1 0 98716 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1073
timestamp 1636968456
transform 1 0 99820 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1085
timestamp 1
transform 1 0 100924 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1091
timestamp 1
transform 1 0 101476 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1093
timestamp 1636968456
transform 1 0 101660 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1105
timestamp 1636968456
transform 1 0 102764 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1117
timestamp 1636968456
transform 1 0 103868 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1129
timestamp 1636968456
transform 1 0 104972 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1141
timestamp 1
transform 1 0 106076 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1147
timestamp 1
transform 1 0 106628 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1149
timestamp 1636968456
transform 1 0 106812 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1161
timestamp 1636968456
transform 1 0 107916 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1173
timestamp 1636968456
transform 1 0 109020 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_1185
timestamp 1
transform 1 0 110124 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1189
timestamp 1
transform 1 0 110492 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636968456
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636968456
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636968456
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_39
timestamp 1636968456
transform 1 0 4692 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1
transform 1 0 5796 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1636968456
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_69
timestamp 1636968456
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_81
timestamp 1636968456
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_93
timestamp 1636968456
transform 1 0 9660 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_105
timestamp 1
transform 1 0 10764 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_111
timestamp 1
transform 1 0 11316 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_113
timestamp 1636968456
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_125
timestamp 1636968456
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_137
timestamp 1636968456
transform 1 0 13708 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_149
timestamp 1636968456
transform 1 0 14812 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1
transform 1 0 15916 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_169
timestamp 1636968456
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_181
timestamp 1636968456
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_193
timestamp 1636968456
transform 1 0 18860 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_205
timestamp 1636968456
transform 1 0 19964 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_217
timestamp 1
transform 1 0 21068 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_223
timestamp 1
transform 1 0 21620 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_225
timestamp 1636968456
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_237
timestamp 1636968456
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_249
timestamp 1636968456
transform 1 0 24012 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_261
timestamp 1636968456
transform 1 0 25116 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_273
timestamp 1
transform 1 0 26220 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_279
timestamp 1
transform 1 0 26772 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_281
timestamp 1636968456
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_293
timestamp 1636968456
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_305
timestamp 1636968456
transform 1 0 29164 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_317
timestamp 1636968456
transform 1 0 30268 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_329
timestamp 1
transform 1 0 31372 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_335
timestamp 1
transform 1 0 31924 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_337
timestamp 1636968456
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_349
timestamp 1636968456
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_361
timestamp 1636968456
transform 1 0 34316 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_373
timestamp 1636968456
transform 1 0 35420 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_385
timestamp 1
transform 1 0 36524 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_391
timestamp 1
transform 1 0 37076 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_393
timestamp 1636968456
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_405
timestamp 1636968456
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_417
timestamp 1636968456
transform 1 0 39468 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_429
timestamp 1636968456
transform 1 0 40572 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_441
timestamp 1
transform 1 0 41676 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_447
timestamp 1
transform 1 0 42228 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_449
timestamp 1636968456
transform 1 0 42412 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_461
timestamp 1636968456
transform 1 0 43516 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_473
timestamp 1636968456
transform 1 0 44620 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_485
timestamp 1636968456
transform 1 0 45724 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_497
timestamp 1
transform 1 0 46828 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_503
timestamp 1
transform 1 0 47380 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_505
timestamp 1636968456
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_517
timestamp 1636968456
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_529
timestamp 1636968456
transform 1 0 49772 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_541
timestamp 1636968456
transform 1 0 50876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_553
timestamp 1
transform 1 0 51980 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_559
timestamp 1
transform 1 0 52532 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_561
timestamp 1636968456
transform 1 0 52716 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_573
timestamp 1636968456
transform 1 0 53820 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_585
timestamp 1636968456
transform 1 0 54924 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_597
timestamp 1636968456
transform 1 0 56028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_609
timestamp 1
transform 1 0 57132 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_615
timestamp 1
transform 1 0 57684 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_617
timestamp 1636968456
transform 1 0 57868 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_629
timestamp 1636968456
transform 1 0 58972 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_641
timestamp 1636968456
transform 1 0 60076 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_653
timestamp 1636968456
transform 1 0 61180 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_665
timestamp 1
transform 1 0 62284 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_671
timestamp 1
transform 1 0 62836 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_673
timestamp 1636968456
transform 1 0 63020 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_685
timestamp 1636968456
transform 1 0 64124 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_697
timestamp 1636968456
transform 1 0 65228 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_709
timestamp 1636968456
transform 1 0 66332 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_721
timestamp 1
transform 1 0 67436 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_727
timestamp 1
transform 1 0 67988 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_729
timestamp 1636968456
transform 1 0 68172 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_741
timestamp 1636968456
transform 1 0 69276 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_753
timestamp 1636968456
transform 1 0 70380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_765
timestamp 1636968456
transform 1 0 71484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_777
timestamp 1
transform 1 0 72588 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_783
timestamp 1
transform 1 0 73140 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_785
timestamp 1636968456
transform 1 0 73324 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_797
timestamp 1636968456
transform 1 0 74428 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_809
timestamp 1636968456
transform 1 0 75532 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_821
timestamp 1636968456
transform 1 0 76636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_833
timestamp 1
transform 1 0 77740 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_839
timestamp 1
transform 1 0 78292 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_841
timestamp 1636968456
transform 1 0 78476 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_853
timestamp 1636968456
transform 1 0 79580 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_865
timestamp 1636968456
transform 1 0 80684 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_877
timestamp 1636968456
transform 1 0 81788 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_889
timestamp 1
transform 1 0 82892 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_895
timestamp 1
transform 1 0 83444 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_897
timestamp 1636968456
transform 1 0 83628 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_909
timestamp 1636968456
transform 1 0 84732 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_921
timestamp 1636968456
transform 1 0 85836 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_933
timestamp 1636968456
transform 1 0 86940 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_945
timestamp 1
transform 1 0 88044 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_951
timestamp 1
transform 1 0 88596 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_953
timestamp 1636968456
transform 1 0 88780 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_965
timestamp 1636968456
transform 1 0 89884 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_977
timestamp 1636968456
transform 1 0 90988 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_989
timestamp 1636968456
transform 1 0 92092 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1001
timestamp 1
transform 1 0 93196 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1007
timestamp 1
transform 1 0 93748 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1009
timestamp 1636968456
transform 1 0 93932 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1021
timestamp 1636968456
transform 1 0 95036 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1033
timestamp 1636968456
transform 1 0 96140 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1045
timestamp 1636968456
transform 1 0 97244 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1057
timestamp 1
transform 1 0 98348 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1063
timestamp 1
transform 1 0 98900 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1065
timestamp 1636968456
transform 1 0 99084 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1077
timestamp 1636968456
transform 1 0 100188 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1089
timestamp 1636968456
transform 1 0 101292 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1101
timestamp 1636968456
transform 1 0 102396 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1113
timestamp 1
transform 1 0 103500 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1119
timestamp 1
transform 1 0 104052 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1121
timestamp 1636968456
transform 1 0 104236 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1133
timestamp 1636968456
transform 1 0 105340 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1145
timestamp 1636968456
transform 1 0 106444 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1157
timestamp 1636968456
transform 1 0 107548 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1169
timestamp 1
transform 1 0 108652 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1175
timestamp 1
transform 1 0 109204 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1177
timestamp 1636968456
transform 1 0 109388 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1189
timestamp 1
transform 1 0 110492 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636968456
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636968456
transform 1 0 2484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 1
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1636968456
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_41
timestamp 1636968456
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_53
timestamp 1636968456
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_65
timestamp 1636968456
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_85
timestamp 1636968456
transform 1 0 8924 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_97
timestamp 1636968456
transform 1 0 10028 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_109
timestamp 1636968456
transform 1 0 11132 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_121
timestamp 1636968456
transform 1 0 12236 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_133
timestamp 1
transform 1 0 13340 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_139
timestamp 1
transform 1 0 13892 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_141
timestamp 1636968456
transform 1 0 14076 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_153
timestamp 1636968456
transform 1 0 15180 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_165
timestamp 1636968456
transform 1 0 16284 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_177
timestamp 1636968456
transform 1 0 17388 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_189
timestamp 1
transform 1 0 18492 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_195
timestamp 1
transform 1 0 19044 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_197
timestamp 1636968456
transform 1 0 19228 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_209
timestamp 1636968456
transform 1 0 20332 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_221
timestamp 1636968456
transform 1 0 21436 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_233
timestamp 1636968456
transform 1 0 22540 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_245
timestamp 1
transform 1 0 23644 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_251
timestamp 1
transform 1 0 24196 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_253
timestamp 1636968456
transform 1 0 24380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_265
timestamp 1636968456
transform 1 0 25484 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_277
timestamp 1636968456
transform 1 0 26588 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_289
timestamp 1636968456
transform 1 0 27692 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_301
timestamp 1
transform 1 0 28796 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_307
timestamp 1
transform 1 0 29348 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_309
timestamp 1636968456
transform 1 0 29532 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_321
timestamp 1636968456
transform 1 0 30636 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_333
timestamp 1636968456
transform 1 0 31740 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_345
timestamp 1636968456
transform 1 0 32844 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_357
timestamp 1
transform 1 0 33948 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_363
timestamp 1
transform 1 0 34500 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_365
timestamp 1636968456
transform 1 0 34684 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_377
timestamp 1636968456
transform 1 0 35788 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_389
timestamp 1636968456
transform 1 0 36892 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_401
timestamp 1636968456
transform 1 0 37996 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_413
timestamp 1
transform 1 0 39100 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_419
timestamp 1
transform 1 0 39652 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_421
timestamp 1636968456
transform 1 0 39836 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_433
timestamp 1636968456
transform 1 0 40940 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_445
timestamp 1636968456
transform 1 0 42044 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_457
timestamp 1636968456
transform 1 0 43148 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_469
timestamp 1
transform 1 0 44252 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_475
timestamp 1
transform 1 0 44804 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_477
timestamp 1636968456
transform 1 0 44988 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_489
timestamp 1636968456
transform 1 0 46092 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_501
timestamp 1636968456
transform 1 0 47196 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_513
timestamp 1636968456
transform 1 0 48300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_525
timestamp 1
transform 1 0 49404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_531
timestamp 1
transform 1 0 49956 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_533
timestamp 1636968456
transform 1 0 50140 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_545
timestamp 1636968456
transform 1 0 51244 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_557
timestamp 1636968456
transform 1 0 52348 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_569
timestamp 1636968456
transform 1 0 53452 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_581
timestamp 1
transform 1 0 54556 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_587
timestamp 1
transform 1 0 55108 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_589
timestamp 1636968456
transform 1 0 55292 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_601
timestamp 1636968456
transform 1 0 56396 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_613
timestamp 1636968456
transform 1 0 57500 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_625
timestamp 1636968456
transform 1 0 58604 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_637
timestamp 1
transform 1 0 59708 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_643
timestamp 1
transform 1 0 60260 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_645
timestamp 1636968456
transform 1 0 60444 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_657
timestamp 1636968456
transform 1 0 61548 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_669
timestamp 1636968456
transform 1 0 62652 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_681
timestamp 1636968456
transform 1 0 63756 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_693
timestamp 1
transform 1 0 64860 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_699
timestamp 1
transform 1 0 65412 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_701
timestamp 1636968456
transform 1 0 65596 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_713
timestamp 1636968456
transform 1 0 66700 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_725
timestamp 1636968456
transform 1 0 67804 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_737
timestamp 1636968456
transform 1 0 68908 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_749
timestamp 1
transform 1 0 70012 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_755
timestamp 1
transform 1 0 70564 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_757
timestamp 1636968456
transform 1 0 70748 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_769
timestamp 1636968456
transform 1 0 71852 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_781
timestamp 1636968456
transform 1 0 72956 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_793
timestamp 1636968456
transform 1 0 74060 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_805
timestamp 1
transform 1 0 75164 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_811
timestamp 1
transform 1 0 75716 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_813
timestamp 1636968456
transform 1 0 75900 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_825
timestamp 1636968456
transform 1 0 77004 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_837
timestamp 1636968456
transform 1 0 78108 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_849
timestamp 1636968456
transform 1 0 79212 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_861
timestamp 1
transform 1 0 80316 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_867
timestamp 1
transform 1 0 80868 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_869
timestamp 1636968456
transform 1 0 81052 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_881
timestamp 1636968456
transform 1 0 82156 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_893
timestamp 1636968456
transform 1 0 83260 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_905
timestamp 1636968456
transform 1 0 84364 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_917
timestamp 1
transform 1 0 85468 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_923
timestamp 1
transform 1 0 86020 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_925
timestamp 1636968456
transform 1 0 86204 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_937
timestamp 1636968456
transform 1 0 87308 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_949
timestamp 1636968456
transform 1 0 88412 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_961
timestamp 1636968456
transform 1 0 89516 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_973
timestamp 1
transform 1 0 90620 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_979
timestamp 1
transform 1 0 91172 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_981
timestamp 1636968456
transform 1 0 91356 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_993
timestamp 1636968456
transform 1 0 92460 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1005
timestamp 1636968456
transform 1 0 93564 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1017
timestamp 1636968456
transform 1 0 94668 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1029
timestamp 1
transform 1 0 95772 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1035
timestamp 1
transform 1 0 96324 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1037
timestamp 1636968456
transform 1 0 96508 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1049
timestamp 1636968456
transform 1 0 97612 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1061
timestamp 1636968456
transform 1 0 98716 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1073
timestamp 1636968456
transform 1 0 99820 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1085
timestamp 1
transform 1 0 100924 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1091
timestamp 1
transform 1 0 101476 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1093
timestamp 1636968456
transform 1 0 101660 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1105
timestamp 1636968456
transform 1 0 102764 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1117
timestamp 1636968456
transform 1 0 103868 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1129
timestamp 1636968456
transform 1 0 104972 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1141
timestamp 1
transform 1 0 106076 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1147
timestamp 1
transform 1 0 106628 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1149
timestamp 1636968456
transform 1 0 106812 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1161
timestamp 1636968456
transform 1 0 107916 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1173
timestamp 1636968456
transform 1 0 109020 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_1185
timestamp 1
transform 1 0 110124 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1189
timestamp 1
transform 1 0 110492 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_3
timestamp 1636968456
transform 1 0 1380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_15
timestamp 1636968456
transform 1 0 2484 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_27
timestamp 1636968456
transform 1 0 3588 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_39
timestamp 1636968456
transform 1 0 4692 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1
transform 1 0 5796 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1636968456
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_69
timestamp 1636968456
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_81
timestamp 1636968456
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_93
timestamp 1636968456
transform 1 0 9660 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1
transform 1 0 10764 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1
transform 1 0 11316 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_113
timestamp 1636968456
transform 1 0 11500 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_125
timestamp 1636968456
transform 1 0 12604 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_137
timestamp 1636968456
transform 1 0 13708 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_149
timestamp 1636968456
transform 1 0 14812 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_161
timestamp 1
transform 1 0 15916 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_167
timestamp 1
transform 1 0 16468 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_169
timestamp 1636968456
transform 1 0 16652 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_181
timestamp 1636968456
transform 1 0 17756 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_193
timestamp 1636968456
transform 1 0 18860 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_205
timestamp 1636968456
transform 1 0 19964 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_217
timestamp 1
transform 1 0 21068 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_223
timestamp 1
transform 1 0 21620 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_225
timestamp 1636968456
transform 1 0 21804 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_237
timestamp 1636968456
transform 1 0 22908 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_249
timestamp 1636968456
transform 1 0 24012 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_261
timestamp 1636968456
transform 1 0 25116 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_273
timestamp 1
transform 1 0 26220 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_279
timestamp 1
transform 1 0 26772 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_281
timestamp 1636968456
transform 1 0 26956 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_293
timestamp 1636968456
transform 1 0 28060 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_305
timestamp 1636968456
transform 1 0 29164 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_317
timestamp 1636968456
transform 1 0 30268 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_329
timestamp 1
transform 1 0 31372 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_335
timestamp 1
transform 1 0 31924 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_337
timestamp 1636968456
transform 1 0 32108 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_349
timestamp 1636968456
transform 1 0 33212 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_361
timestamp 1636968456
transform 1 0 34316 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_373
timestamp 1636968456
transform 1 0 35420 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_385
timestamp 1
transform 1 0 36524 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_391
timestamp 1
transform 1 0 37076 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_393
timestamp 1636968456
transform 1 0 37260 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_405
timestamp 1636968456
transform 1 0 38364 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_417
timestamp 1636968456
transform 1 0 39468 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_429
timestamp 1636968456
transform 1 0 40572 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_441
timestamp 1
transform 1 0 41676 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_447
timestamp 1
transform 1 0 42228 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_449
timestamp 1636968456
transform 1 0 42412 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_461
timestamp 1636968456
transform 1 0 43516 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_473
timestamp 1636968456
transform 1 0 44620 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_485
timestamp 1636968456
transform 1 0 45724 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_497
timestamp 1
transform 1 0 46828 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_503
timestamp 1
transform 1 0 47380 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_505
timestamp 1636968456
transform 1 0 47564 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_517
timestamp 1636968456
transform 1 0 48668 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_529
timestamp 1636968456
transform 1 0 49772 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_541
timestamp 1636968456
transform 1 0 50876 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_553
timestamp 1
transform 1 0 51980 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_559
timestamp 1
transform 1 0 52532 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_561
timestamp 1636968456
transform 1 0 52716 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_573
timestamp 1636968456
transform 1 0 53820 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_585
timestamp 1636968456
transform 1 0 54924 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_597
timestamp 1636968456
transform 1 0 56028 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_609
timestamp 1
transform 1 0 57132 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_615
timestamp 1
transform 1 0 57684 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_617
timestamp 1636968456
transform 1 0 57868 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_629
timestamp 1636968456
transform 1 0 58972 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_641
timestamp 1636968456
transform 1 0 60076 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_653
timestamp 1636968456
transform 1 0 61180 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_665
timestamp 1
transform 1 0 62284 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_671
timestamp 1
transform 1 0 62836 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_673
timestamp 1636968456
transform 1 0 63020 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_685
timestamp 1636968456
transform 1 0 64124 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_697
timestamp 1636968456
transform 1 0 65228 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_709
timestamp 1636968456
transform 1 0 66332 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_721
timestamp 1
transform 1 0 67436 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_727
timestamp 1
transform 1 0 67988 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_729
timestamp 1636968456
transform 1 0 68172 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_741
timestamp 1636968456
transform 1 0 69276 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_753
timestamp 1636968456
transform 1 0 70380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_765
timestamp 1636968456
transform 1 0 71484 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_777
timestamp 1
transform 1 0 72588 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_783
timestamp 1
transform 1 0 73140 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_785
timestamp 1636968456
transform 1 0 73324 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_797
timestamp 1636968456
transform 1 0 74428 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_809
timestamp 1636968456
transform 1 0 75532 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_821
timestamp 1636968456
transform 1 0 76636 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_833
timestamp 1
transform 1 0 77740 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_839
timestamp 1
transform 1 0 78292 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_841
timestamp 1636968456
transform 1 0 78476 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_853
timestamp 1636968456
transform 1 0 79580 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_865
timestamp 1636968456
transform 1 0 80684 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_877
timestamp 1636968456
transform 1 0 81788 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_889
timestamp 1
transform 1 0 82892 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_895
timestamp 1
transform 1 0 83444 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_897
timestamp 1636968456
transform 1 0 83628 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_909
timestamp 1636968456
transform 1 0 84732 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_921
timestamp 1636968456
transform 1 0 85836 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_933
timestamp 1636968456
transform 1 0 86940 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_945
timestamp 1
transform 1 0 88044 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_951
timestamp 1
transform 1 0 88596 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_953
timestamp 1636968456
transform 1 0 88780 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_965
timestamp 1636968456
transform 1 0 89884 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_977
timestamp 1636968456
transform 1 0 90988 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_989
timestamp 1636968456
transform 1 0 92092 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1001
timestamp 1
transform 1 0 93196 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1007
timestamp 1
transform 1 0 93748 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1009
timestamp 1636968456
transform 1 0 93932 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1021
timestamp 1636968456
transform 1 0 95036 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1033
timestamp 1636968456
transform 1 0 96140 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1045
timestamp 1636968456
transform 1 0 97244 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1057
timestamp 1
transform 1 0 98348 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1063
timestamp 1
transform 1 0 98900 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1065
timestamp 1636968456
transform 1 0 99084 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1077
timestamp 1636968456
transform 1 0 100188 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1089
timestamp 1636968456
transform 1 0 101292 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1101
timestamp 1636968456
transform 1 0 102396 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1113
timestamp 1
transform 1 0 103500 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1119
timestamp 1
transform 1 0 104052 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1121
timestamp 1636968456
transform 1 0 104236 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1133
timestamp 1636968456
transform 1 0 105340 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1145
timestamp 1636968456
transform 1 0 106444 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1157
timestamp 1636968456
transform 1 0 107548 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1169
timestamp 1
transform 1 0 108652 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1175
timestamp 1
transform 1 0 109204 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1177
timestamp 1636968456
transform 1 0 109388 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1189
timestamp 1
transform 1 0 110492 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636968456
transform 1 0 1380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636968456
transform 1 0 2484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 1
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636968456
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1636968456
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_53
timestamp 1636968456
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_65
timestamp 1636968456
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_85
timestamp 1636968456
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_97
timestamp 1636968456
transform 1 0 10028 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_109
timestamp 1636968456
transform 1 0 11132 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_121
timestamp 1636968456
transform 1 0 12236 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_133
timestamp 1
transform 1 0 13340 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_139
timestamp 1
transform 1 0 13892 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_141
timestamp 1636968456
transform 1 0 14076 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_153
timestamp 1636968456
transform 1 0 15180 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_165
timestamp 1636968456
transform 1 0 16284 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_177
timestamp 1636968456
transform 1 0 17388 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_189
timestamp 1
transform 1 0 18492 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_195
timestamp 1
transform 1 0 19044 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_197
timestamp 1636968456
transform 1 0 19228 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_209
timestamp 1636968456
transform 1 0 20332 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_221
timestamp 1636968456
transform 1 0 21436 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_233
timestamp 1636968456
transform 1 0 22540 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_245
timestamp 1
transform 1 0 23644 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_251
timestamp 1
transform 1 0 24196 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_253
timestamp 1636968456
transform 1 0 24380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_265
timestamp 1636968456
transform 1 0 25484 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_277
timestamp 1636968456
transform 1 0 26588 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_289
timestamp 1636968456
transform 1 0 27692 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_301
timestamp 1
transform 1 0 28796 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_307
timestamp 1
transform 1 0 29348 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_309
timestamp 1636968456
transform 1 0 29532 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_321
timestamp 1636968456
transform 1 0 30636 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_333
timestamp 1636968456
transform 1 0 31740 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_345
timestamp 1636968456
transform 1 0 32844 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_357
timestamp 1
transform 1 0 33948 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_363
timestamp 1
transform 1 0 34500 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_365
timestamp 1636968456
transform 1 0 34684 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_377
timestamp 1636968456
transform 1 0 35788 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_389
timestamp 1636968456
transform 1 0 36892 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_401
timestamp 1636968456
transform 1 0 37996 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_413
timestamp 1
transform 1 0 39100 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_419
timestamp 1
transform 1 0 39652 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_421
timestamp 1636968456
transform 1 0 39836 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_433
timestamp 1636968456
transform 1 0 40940 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_445
timestamp 1636968456
transform 1 0 42044 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_457
timestamp 1636968456
transform 1 0 43148 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_469
timestamp 1
transform 1 0 44252 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_475
timestamp 1
transform 1 0 44804 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_477
timestamp 1636968456
transform 1 0 44988 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_489
timestamp 1636968456
transform 1 0 46092 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_501
timestamp 1636968456
transform 1 0 47196 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_513
timestamp 1636968456
transform 1 0 48300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_525
timestamp 1
transform 1 0 49404 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_531
timestamp 1
transform 1 0 49956 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_533
timestamp 1636968456
transform 1 0 50140 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_545
timestamp 1636968456
transform 1 0 51244 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_557
timestamp 1636968456
transform 1 0 52348 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_569
timestamp 1636968456
transform 1 0 53452 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_581
timestamp 1
transform 1 0 54556 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_587
timestamp 1
transform 1 0 55108 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_589
timestamp 1636968456
transform 1 0 55292 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_601
timestamp 1636968456
transform 1 0 56396 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_613
timestamp 1636968456
transform 1 0 57500 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_625
timestamp 1636968456
transform 1 0 58604 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_637
timestamp 1
transform 1 0 59708 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_643
timestamp 1
transform 1 0 60260 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_645
timestamp 1636968456
transform 1 0 60444 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_657
timestamp 1636968456
transform 1 0 61548 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_669
timestamp 1636968456
transform 1 0 62652 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_681
timestamp 1636968456
transform 1 0 63756 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_693
timestamp 1
transform 1 0 64860 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_699
timestamp 1
transform 1 0 65412 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_701
timestamp 1636968456
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_713
timestamp 1636968456
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_725
timestamp 1636968456
transform 1 0 67804 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_737
timestamp 1636968456
transform 1 0 68908 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_749
timestamp 1
transform 1 0 70012 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_755
timestamp 1
transform 1 0 70564 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_757
timestamp 1636968456
transform 1 0 70748 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_769
timestamp 1636968456
transform 1 0 71852 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_781
timestamp 1636968456
transform 1 0 72956 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_793
timestamp 1636968456
transform 1 0 74060 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_805
timestamp 1
transform 1 0 75164 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_811
timestamp 1
transform 1 0 75716 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_813
timestamp 1636968456
transform 1 0 75900 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_825
timestamp 1636968456
transform 1 0 77004 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_837
timestamp 1636968456
transform 1 0 78108 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_849
timestamp 1636968456
transform 1 0 79212 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_861
timestamp 1
transform 1 0 80316 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_867
timestamp 1
transform 1 0 80868 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_869
timestamp 1636968456
transform 1 0 81052 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_881
timestamp 1636968456
transform 1 0 82156 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_893
timestamp 1636968456
transform 1 0 83260 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_905
timestamp 1636968456
transform 1 0 84364 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_917
timestamp 1
transform 1 0 85468 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_923
timestamp 1
transform 1 0 86020 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_925
timestamp 1636968456
transform 1 0 86204 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_937
timestamp 1636968456
transform 1 0 87308 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_949
timestamp 1636968456
transform 1 0 88412 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_961
timestamp 1636968456
transform 1 0 89516 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_973
timestamp 1
transform 1 0 90620 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_979
timestamp 1
transform 1 0 91172 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_981
timestamp 1636968456
transform 1 0 91356 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_993
timestamp 1636968456
transform 1 0 92460 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1005
timestamp 1636968456
transform 1 0 93564 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1017
timestamp 1636968456
transform 1 0 94668 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1029
timestamp 1
transform 1 0 95772 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1035
timestamp 1
transform 1 0 96324 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1037
timestamp 1636968456
transform 1 0 96508 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1049
timestamp 1636968456
transform 1 0 97612 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1061
timestamp 1636968456
transform 1 0 98716 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1073
timestamp 1636968456
transform 1 0 99820 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1085
timestamp 1
transform 1 0 100924 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1091
timestamp 1
transform 1 0 101476 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1093
timestamp 1636968456
transform 1 0 101660 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1105
timestamp 1636968456
transform 1 0 102764 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1117
timestamp 1636968456
transform 1 0 103868 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1129
timestamp 1636968456
transform 1 0 104972 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1141
timestamp 1
transform 1 0 106076 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1147
timestamp 1
transform 1 0 106628 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1149
timestamp 1636968456
transform 1 0 106812 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1161
timestamp 1636968456
transform 1 0 107916 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1173
timestamp 1636968456
transform 1 0 109020 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_1185
timestamp 1
transform 1 0 110124 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1189
timestamp 1
transform 1 0 110492 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1636968456
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1636968456
transform 1 0 2484 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_127_27
timestamp 1
transform 1 0 3588 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_29
timestamp 1636968456
transform 1 0 3772 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_41
timestamp 1636968456
transform 1 0 4876 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_53
timestamp 1
transform 1 0 5980 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1636968456
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_69
timestamp 1636968456
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_81
timestamp 1
transform 1 0 8556 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_85
timestamp 1636968456
transform 1 0 8924 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_97
timestamp 1636968456
transform 1 0 10028 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_109
timestamp 1
transform 1 0 11132 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_113
timestamp 1636968456
transform 1 0 11500 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_125
timestamp 1636968456
transform 1 0 12604 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_137
timestamp 1
transform 1 0 13708 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_141
timestamp 1636968456
transform 1 0 14076 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_153
timestamp 1636968456
transform 1 0 15180 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_165
timestamp 1
transform 1 0 16284 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_169
timestamp 1636968456
transform 1 0 16652 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_181
timestamp 1636968456
transform 1 0 17756 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_193
timestamp 1
transform 1 0 18860 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_197
timestamp 1636968456
transform 1 0 19228 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_209
timestamp 1636968456
transform 1 0 20332 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_221
timestamp 1
transform 1 0 21436 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_225
timestamp 1636968456
transform 1 0 21804 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_237
timestamp 1636968456
transform 1 0 22908 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_249
timestamp 1
transform 1 0 24012 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_253
timestamp 1636968456
transform 1 0 24380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_265
timestamp 1636968456
transform 1 0 25484 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_277
timestamp 1
transform 1 0 26588 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_281
timestamp 1636968456
transform 1 0 26956 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_293
timestamp 1636968456
transform 1 0 28060 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_305
timestamp 1
transform 1 0 29164 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_309
timestamp 1636968456
transform 1 0 29532 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_321
timestamp 1636968456
transform 1 0 30636 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_333
timestamp 1
transform 1 0 31740 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_337
timestamp 1636968456
transform 1 0 32108 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_349
timestamp 1636968456
transform 1 0 33212 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_361
timestamp 1
transform 1 0 34316 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_365
timestamp 1636968456
transform 1 0 34684 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_377
timestamp 1636968456
transform 1 0 35788 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_389
timestamp 1
transform 1 0 36892 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_393
timestamp 1636968456
transform 1 0 37260 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_405
timestamp 1636968456
transform 1 0 38364 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_417
timestamp 1
transform 1 0 39468 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_421
timestamp 1636968456
transform 1 0 39836 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_433
timestamp 1636968456
transform 1 0 40940 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_445
timestamp 1
transform 1 0 42044 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_449
timestamp 1636968456
transform 1 0 42412 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_461
timestamp 1
transform 1 0 43516 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_127_469
timestamp 1
transform 1 0 44252 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_477
timestamp 1636968456
transform 1 0 44988 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_489
timestamp 1
transform 1 0 46092 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_127_497
timestamp 1
transform 1 0 46828 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_505
timestamp 1636968456
transform 1 0 47564 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_517
timestamp 1
transform 1 0 48668 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_127_525
timestamp 1
transform 1 0 49404 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_533
timestamp 1636968456
transform 1 0 50140 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_545
timestamp 1
transform 1 0 51244 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_127_553
timestamp 1
transform 1 0 51980 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_559
timestamp 1
transform 1 0 52532 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_561
timestamp 1
transform 1 0 52716 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_569
timestamp 1
transform 1 0 53452 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_574
timestamp 1636968456
transform 1 0 53912 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_586
timestamp 1
transform 1 0 55016 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_127_589
timestamp 1
transform 1 0 55292 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_127_595
timestamp 1636968456
transform 1 0 55844 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_607
timestamp 1
transform 1 0 56948 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_611
timestamp 1
transform 1 0 57316 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_617
timestamp 1636968456
transform 1 0 57868 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_629
timestamp 1
transform 1 0 58972 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_127_637
timestamp 1
transform 1 0 59708 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_643
timestamp 1
transform 1 0 60260 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_645
timestamp 1
transform 1 0 60444 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_653
timestamp 1
transform 1 0 61180 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_658
timestamp 1636968456
transform 1 0 61640 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_670
timestamp 1
transform 1 0 62744 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_127_673
timestamp 1
transform 1 0 63020 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_127_679
timestamp 1636968456
transform 1 0 63572 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_691
timestamp 1
transform 1 0 64676 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_699
timestamp 1
transform 1 0 65412 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_127_701
timestamp 1
transform 1 0 65596 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_127_707
timestamp 1636968456
transform 1 0 66148 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_719
timestamp 1
transform 1 0 67252 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_723
timestamp 1
transform 1 0 67620 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_729
timestamp 1636968456
transform 1 0 68172 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_741
timestamp 1
transform 1 0 69276 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_127_749
timestamp 1
transform 1 0 70012 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_755
timestamp 1
transform 1 0 70564 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_757
timestamp 1
transform 1 0 70748 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_765
timestamp 1
transform 1 0 71484 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_770
timestamp 1636968456
transform 1 0 71944 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_782
timestamp 1
transform 1 0 73048 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_127_785
timestamp 1
transform 1 0 73324 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_793
timestamp 1
transform 1 0 74060 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_798
timestamp 1636968456
transform 1 0 74520 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_127_810
timestamp 1
transform 1 0 75624 0 -1 71808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_127_813
timestamp 1636968456
transform 1 0 75900 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_825
timestamp 1
transform 1 0 77004 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_127_833
timestamp 1
transform 1 0 77740 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_839
timestamp 1
transform 1 0 78292 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_841
timestamp 1636968456
transform 1 0 78476 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_853
timestamp 1636968456
transform 1 0 79580 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_865
timestamp 1
transform 1 0 80684 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_869
timestamp 1636968456
transform 1 0 81052 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_881
timestamp 1636968456
transform 1 0 82156 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_893
timestamp 1
transform 1 0 83260 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_897
timestamp 1636968456
transform 1 0 83628 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_909
timestamp 1636968456
transform 1 0 84732 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_921
timestamp 1
transform 1 0 85836 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_925
timestamp 1636968456
transform 1 0 86204 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_937
timestamp 1636968456
transform 1 0 87308 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_949
timestamp 1
transform 1 0 88412 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_953
timestamp 1636968456
transform 1 0 88780 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_965
timestamp 1636968456
transform 1 0 89884 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_977
timestamp 1
transform 1 0 90988 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_981
timestamp 1636968456
transform 1 0 91356 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_993
timestamp 1636968456
transform 1 0 92460 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1005
timestamp 1
transform 1 0 93564 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1009
timestamp 1636968456
transform 1 0 93932 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1021
timestamp 1636968456
transform 1 0 95036 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1033
timestamp 1
transform 1 0 96140 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1037
timestamp 1636968456
transform 1 0 96508 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1049
timestamp 1636968456
transform 1 0 97612 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1061
timestamp 1
transform 1 0 98716 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1065
timestamp 1636968456
transform 1 0 99084 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1077
timestamp 1636968456
transform 1 0 100188 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1089
timestamp 1
transform 1 0 101292 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1093
timestamp 1636968456
transform 1 0 101660 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1105
timestamp 1636968456
transform 1 0 102764 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1117
timestamp 1
transform 1 0 103868 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1121
timestamp 1636968456
transform 1 0 104236 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1133
timestamp 1636968456
transform 1 0 105340 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1145
timestamp 1
transform 1 0 106444 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1149
timestamp 1636968456
transform 1 0 106812 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1161
timestamp 1636968456
transform 1 0 107916 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_1173
timestamp 1
transform 1 0 109020 0 -1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1177
timestamp 1636968456
transform 1 0 109388 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1189
timestamp 1
transform 1 0 110492 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 105156 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 104696 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 105156 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform 1 0 104696 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1
transform -1 0 110584 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i_21
timestamp 1
transform -1 0 104604 0 1 59840
box -38 -48 314 592
use ram256x16  mem_i
timestamp 0
transform 1 0 10000 0 1 10000
box 0 0 1 1
use sky130_fd_sc_hd__buf_2  output2
timestamp 1
transform -1 0 44896 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1
transform 1 0 65780 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1
transform 1 0 67712 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1
transform -1 0 70012 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1
transform -1 0 71944 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1
transform 1 0 74152 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1
transform 1 0 77372 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1
transform -1 0 47472 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform 1 0 49680 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform 1 0 51612 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 53544 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform 1 0 55476 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform 1 0 57408 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform -1 0 59708 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1
transform -1 0 61640 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform 1 0 63204 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_128
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 110860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_129
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 110860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_130
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 110860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_131
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 110860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_132
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 110860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_133
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 110860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_134
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 110860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_135
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 110860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_136
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 110860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_137
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 110860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_255
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_469
timestamp 1
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_256
timestamp 1
transform 1 0 104052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_21
timestamp 1
transform -1 0 110860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_138
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_363
timestamp 1
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_257
timestamp 1
transform 1 0 104052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_22
timestamp 1
transform -1 0 110860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_139
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_364
timestamp 1
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_258
timestamp 1
transform 1 0 104052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_23
timestamp 1
transform -1 0 110860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_140
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_365
timestamp 1
transform -1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_259
timestamp 1
transform 1 0 104052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_24
timestamp 1
transform -1 0 110860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_141
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_366
timestamp 1
transform -1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_260
timestamp 1
transform 1 0 104052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_25
timestamp 1
transform -1 0 110860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_142
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_367
timestamp 1
transform -1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_261
timestamp 1
transform 1 0 104052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_26
timestamp 1
transform -1 0 110860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_143
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_368
timestamp 1
transform -1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_262
timestamp 1
transform 1 0 104052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_27
timestamp 1
transform -1 0 110860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_144
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_369
timestamp 1
transform -1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_263
timestamp 1
transform 1 0 104052 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_28
timestamp 1
transform -1 0 110860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_145
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_370
timestamp 1
transform -1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_264
timestamp 1
transform 1 0 104052 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_29
timestamp 1
transform -1 0 110860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_146
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_371
timestamp 1
transform -1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_265
timestamp 1
transform 1 0 104052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_30
timestamp 1
transform -1 0 110860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_147
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_372
timestamp 1
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_266
timestamp 1
transform 1 0 104052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_31
timestamp 1
transform -1 0 110860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_148
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_373
timestamp 1
transform -1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_267
timestamp 1
transform 1 0 104052 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_32
timestamp 1
transform -1 0 110860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_149
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_374
timestamp 1
transform -1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_268
timestamp 1
transform 1 0 104052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_33
timestamp 1
transform -1 0 110860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_150
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_375
timestamp 1
transform -1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_269
timestamp 1
transform 1 0 104052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_34
timestamp 1
transform -1 0 110860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_151
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_376
timestamp 1
transform -1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_270
timestamp 1
transform 1 0 104052 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_35
timestamp 1
transform -1 0 110860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_152
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_377
timestamp 1
transform -1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_271
timestamp 1
transform 1 0 104052 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_36
timestamp 1
transform -1 0 110860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_153
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_378
timestamp 1
transform -1 0 7912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_272
timestamp 1
transform 1 0 104052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_37
timestamp 1
transform -1 0 110860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_154
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_379
timestamp 1
transform -1 0 7912 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_273
timestamp 1
transform 1 0 104052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_38
timestamp 1
transform -1 0 110860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_155
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_380
timestamp 1
transform -1 0 7912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_274
timestamp 1
transform 1 0 104052 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_39
timestamp 1
transform -1 0 110860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_156
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_381
timestamp 1
transform -1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_275
timestamp 1
transform 1 0 104052 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_40
timestamp 1
transform -1 0 110860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_157
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_382
timestamp 1
transform -1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_276
timestamp 1
transform 1 0 104052 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_41
timestamp 1
transform -1 0 110860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_158
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_383
timestamp 1
transform -1 0 7912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_277
timestamp 1
transform 1 0 104052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_42
timestamp 1
transform -1 0 110860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_159
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_384
timestamp 1
transform -1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_278
timestamp 1
transform 1 0 104052 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_43
timestamp 1
transform -1 0 110860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_160
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_385
timestamp 1
transform -1 0 7912 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_279
timestamp 1
transform 1 0 104052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_44
timestamp 1
transform -1 0 110860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_161
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_386
timestamp 1
transform -1 0 7912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_280
timestamp 1
transform 1 0 104052 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_45
timestamp 1
transform -1 0 110860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_162
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_387
timestamp 1
transform -1 0 7912 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_281
timestamp 1
transform 1 0 104052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_46
timestamp 1
transform -1 0 110860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_163
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_388
timestamp 1
transform -1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_282
timestamp 1
transform 1 0 104052 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_47
timestamp 1
transform -1 0 110860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_164
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_389
timestamp 1
transform -1 0 7912 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_283
timestamp 1
transform 1 0 104052 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_48
timestamp 1
transform -1 0 110860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_165
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_390
timestamp 1
transform -1 0 7912 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_284
timestamp 1
transform 1 0 104052 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_49
timestamp 1
transform -1 0 110860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_166
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_391
timestamp 1
transform -1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_285
timestamp 1
transform 1 0 104052 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_50
timestamp 1
transform -1 0 110860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_167
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_392
timestamp 1
transform -1 0 7912 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_286
timestamp 1
transform 1 0 104052 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_51
timestamp 1
transform -1 0 110860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_168
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_393
timestamp 1
transform -1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_287
timestamp 1
transform 1 0 104052 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_52
timestamp 1
transform -1 0 110860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_169
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_394
timestamp 1
transform -1 0 7912 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_288
timestamp 1
transform 1 0 104052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_53
timestamp 1
transform -1 0 110860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_170
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_395
timestamp 1
transform -1 0 7912 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_289
timestamp 1
transform 1 0 104052 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_54
timestamp 1
transform -1 0 110860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_171
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_396
timestamp 1
transform -1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_290
timestamp 1
transform 1 0 104052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_55
timestamp 1
transform -1 0 110860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_172
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_397
timestamp 1
transform -1 0 7912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_291
timestamp 1
transform 1 0 104052 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_56
timestamp 1
transform -1 0 110860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_173
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_398
timestamp 1
transform -1 0 7912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_292
timestamp 1
transform 1 0 104052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_57
timestamp 1
transform -1 0 110860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_174
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_399
timestamp 1
transform -1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_293
timestamp 1
transform 1 0 104052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_58
timestamp 1
transform -1 0 110860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_175
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_400
timestamp 1
transform -1 0 7912 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_294
timestamp 1
transform 1 0 104052 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_59
timestamp 1
transform -1 0 110860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_176
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_401
timestamp 1
transform -1 0 7912 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_295
timestamp 1
transform 1 0 104052 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_60
timestamp 1
transform -1 0 110860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_177
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_402
timestamp 1
transform -1 0 7912 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_296
timestamp 1
transform 1 0 104052 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_61
timestamp 1
transform -1 0 110860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_178
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_403
timestamp 1
transform -1 0 7912 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_297
timestamp 1
transform 1 0 104052 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_62
timestamp 1
transform -1 0 110860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_179
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_404
timestamp 1
transform -1 0 7912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_298
timestamp 1
transform 1 0 104052 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_63
timestamp 1
transform -1 0 110860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_180
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_405
timestamp 1
transform -1 0 7912 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_299
timestamp 1
transform 1 0 104052 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_64
timestamp 1
transform -1 0 110860 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_181
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_406
timestamp 1
transform -1 0 7912 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_300
timestamp 1
transform 1 0 104052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_65
timestamp 1
transform -1 0 110860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_182
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_407
timestamp 1
transform -1 0 7912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_301
timestamp 1
transform 1 0 104052 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_66
timestamp 1
transform -1 0 110860 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_183
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_408
timestamp 1
transform -1 0 7912 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_302
timestamp 1
transform 1 0 104052 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_67
timestamp 1
transform -1 0 110860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_184
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_409
timestamp 1
transform -1 0 7912 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_303
timestamp 1
transform 1 0 104052 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_68
timestamp 1
transform -1 0 110860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_185
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_410
timestamp 1
transform -1 0 7912 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_304
timestamp 1
transform 1 0 104052 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_69
timestamp 1
transform -1 0 110860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_186
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_411
timestamp 1
transform -1 0 7912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_305
timestamp 1
transform 1 0 104052 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_70
timestamp 1
transform -1 0 110860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_187
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_412
timestamp 1
transform -1 0 7912 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_306
timestamp 1
transform 1 0 104052 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_71
timestamp 1
transform -1 0 110860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_188
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_413
timestamp 1
transform -1 0 7912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_307
timestamp 1
transform 1 0 104052 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_72
timestamp 1
transform -1 0 110860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_189
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_414
timestamp 1
transform -1 0 7912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_308
timestamp 1
transform 1 0 104052 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_73
timestamp 1
transform -1 0 110860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_190
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_415
timestamp 1
transform -1 0 7912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_309
timestamp 1
transform 1 0 104052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_74
timestamp 1
transform -1 0 110860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_191
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_416
timestamp 1
transform -1 0 7912 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_310
timestamp 1
transform 1 0 104052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_75
timestamp 1
transform -1 0 110860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_192
timestamp 1
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_417
timestamp 1
transform -1 0 7912 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_311
timestamp 1
transform 1 0 104052 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_76
timestamp 1
transform -1 0 110860 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_193
timestamp 1
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_418
timestamp 1
transform -1 0 7912 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_312
timestamp 1
transform 1 0 104052 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_77
timestamp 1
transform -1 0 110860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_194
timestamp 1
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_419
timestamp 1
transform -1 0 7912 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_313
timestamp 1
transform 1 0 104052 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_78
timestamp 1
transform -1 0 110860 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_195
timestamp 1
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_420
timestamp 1
transform -1 0 7912 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_314
timestamp 1
transform 1 0 104052 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_79
timestamp 1
transform -1 0 110860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_196
timestamp 1
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_421
timestamp 1
transform -1 0 7912 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_315
timestamp 1
transform 1 0 104052 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_80
timestamp 1
transform -1 0 110860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_197
timestamp 1
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_422
timestamp 1
transform -1 0 7912 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_316
timestamp 1
transform 1 0 104052 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_81
timestamp 1
transform -1 0 110860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_198
timestamp 1
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_423
timestamp 1
transform -1 0 7912 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_317
timestamp 1
transform 1 0 104052 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_82
timestamp 1
transform -1 0 110860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_199
timestamp 1
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_424
timestamp 1
transform -1 0 7912 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_318
timestamp 1
transform 1 0 104052 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_83
timestamp 1
transform -1 0 110860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_200
timestamp 1
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_425
timestamp 1
transform -1 0 7912 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_319
timestamp 1
transform 1 0 104052 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_84
timestamp 1
transform -1 0 110860 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_201
timestamp 1
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_426
timestamp 1
transform -1 0 7912 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_320
timestamp 1
transform 1 0 104052 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_85
timestamp 1
transform -1 0 110860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_202
timestamp 1
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_427
timestamp 1
transform -1 0 7912 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_321
timestamp 1
transform 1 0 104052 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_86
timestamp 1
transform -1 0 110860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_203
timestamp 1
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_428
timestamp 1
transform -1 0 7912 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_322
timestamp 1
transform 1 0 104052 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_87
timestamp 1
transform -1 0 110860 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_204
timestamp 1
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_429
timestamp 1
transform -1 0 7912 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_323
timestamp 1
transform 1 0 104052 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_88
timestamp 1
transform -1 0 110860 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_205
timestamp 1
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_430
timestamp 1
transform -1 0 7912 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_324
timestamp 1
transform 1 0 104052 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_89
timestamp 1
transform -1 0 110860 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_206
timestamp 1
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_431
timestamp 1
transform -1 0 7912 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_325
timestamp 1
transform 1 0 104052 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_90
timestamp 1
transform -1 0 110860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_207
timestamp 1
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_432
timestamp 1
transform -1 0 7912 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_326
timestamp 1
transform 1 0 104052 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_91
timestamp 1
transform -1 0 110860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_208
timestamp 1
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_433
timestamp 1
transform -1 0 7912 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_327
timestamp 1
transform 1 0 104052 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_92
timestamp 1
transform -1 0 110860 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_209
timestamp 1
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_434
timestamp 1
transform -1 0 7912 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_328
timestamp 1
transform 1 0 104052 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_93
timestamp 1
transform -1 0 110860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_210
timestamp 1
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_435
timestamp 1
transform -1 0 7912 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_329
timestamp 1
transform 1 0 104052 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_94
timestamp 1
transform -1 0 110860 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_211
timestamp 1
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_436
timestamp 1
transform -1 0 7912 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_330
timestamp 1
transform 1 0 104052 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_95
timestamp 1
transform -1 0 110860 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_212
timestamp 1
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_437
timestamp 1
transform -1 0 7912 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_331
timestamp 1
transform 1 0 104052 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_96
timestamp 1
transform -1 0 110860 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_213
timestamp 1
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_438
timestamp 1
transform -1 0 7912 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_332
timestamp 1
transform 1 0 104052 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_97
timestamp 1
transform -1 0 110860 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_214
timestamp 1
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_439
timestamp 1
transform -1 0 7912 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_333
timestamp 1
transform 1 0 104052 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_98
timestamp 1
transform -1 0 110860 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_215
timestamp 1
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_440
timestamp 1
transform -1 0 7912 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_334
timestamp 1
transform 1 0 104052 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_99
timestamp 1
transform -1 0 110860 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_216
timestamp 1
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_441
timestamp 1
transform -1 0 7912 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_335
timestamp 1
transform 1 0 104052 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_100
timestamp 1
transform -1 0 110860 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_217
timestamp 1
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_442
timestamp 1
transform -1 0 7912 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_336
timestamp 1
transform 1 0 104052 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_101
timestamp 1
transform -1 0 110860 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_218
timestamp 1
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_443
timestamp 1
transform -1 0 7912 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_337
timestamp 1
transform 1 0 104052 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_102
timestamp 1
transform -1 0 110860 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_219
timestamp 1
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_444
timestamp 1
transform -1 0 7912 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_338
timestamp 1
transform 1 0 104052 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_103
timestamp 1
transform -1 0 110860 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_220
timestamp 1
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_445
timestamp 1
transform -1 0 7912 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_339
timestamp 1
transform 1 0 104052 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_104
timestamp 1
transform -1 0 110860 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_221
timestamp 1
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_446
timestamp 1
transform -1 0 7912 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_340
timestamp 1
transform 1 0 104052 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_105
timestamp 1
transform -1 0 110860 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_222
timestamp 1
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_447
timestamp 1
transform -1 0 7912 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_341
timestamp 1
transform 1 0 104052 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_106
timestamp 1
transform -1 0 110860 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_223
timestamp 1
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_448
timestamp 1
transform -1 0 7912 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_342
timestamp 1
transform 1 0 104052 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_107
timestamp 1
transform -1 0 110860 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_224
timestamp 1
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_449
timestamp 1
transform -1 0 7912 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_343
timestamp 1
transform 1 0 104052 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_108
timestamp 1
transform -1 0 110860 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_225
timestamp 1
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_450
timestamp 1
transform -1 0 7912 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_344
timestamp 1
transform 1 0 104052 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_109
timestamp 1
transform -1 0 110860 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_226
timestamp 1
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_451
timestamp 1
transform -1 0 7912 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_345
timestamp 1
transform 1 0 104052 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_110
timestamp 1
transform -1 0 110860 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_227
timestamp 1
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_452
timestamp 1
transform -1 0 7912 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_346
timestamp 1
transform 1 0 104052 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_111
timestamp 1
transform -1 0 110860 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_228
timestamp 1
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_453
timestamp 1
transform -1 0 7912 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_347
timestamp 1
transform 1 0 104052 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_112
timestamp 1
transform -1 0 110860 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_229
timestamp 1
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_454
timestamp 1
transform -1 0 7912 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_348
timestamp 1
transform 1 0 104052 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_113
timestamp 1
transform -1 0 110860 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_230
timestamp 1
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_455
timestamp 1
transform -1 0 7912 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_349
timestamp 1
transform 1 0 104052 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_114
timestamp 1
transform -1 0 110860 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_231
timestamp 1
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_456
timestamp 1
transform -1 0 7912 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_350
timestamp 1
transform 1 0 104052 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_115
timestamp 1
transform -1 0 110860 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_232
timestamp 1
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_457
timestamp 1
transform -1 0 7912 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_351
timestamp 1
transform 1 0 104052 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_116
timestamp 1
transform -1 0 110860 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_233
timestamp 1
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_458
timestamp 1
transform -1 0 7912 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_352
timestamp 1
transform 1 0 104052 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_117
timestamp 1
transform -1 0 110860 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_234
timestamp 1
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_459
timestamp 1
transform -1 0 7912 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_353
timestamp 1
transform 1 0 104052 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_118
timestamp 1
transform -1 0 110860 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_235
timestamp 1
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_460
timestamp 1
transform -1 0 7912 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_354
timestamp 1
transform 1 0 104052 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_119
timestamp 1
transform -1 0 110860 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_236
timestamp 1
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_461
timestamp 1
transform -1 0 7912 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_355
timestamp 1
transform 1 0 104052 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_120
timestamp 1
transform -1 0 110860 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_237
timestamp 1
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_462
timestamp 1
transform -1 0 7912 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_356
timestamp 1
transform 1 0 104052 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_121
timestamp 1
transform -1 0 110860 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_238
timestamp 1
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_463
timestamp 1
transform -1 0 7912 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_357
timestamp 1
transform 1 0 104052 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_122
timestamp 1
transform -1 0 110860 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_239
timestamp 1
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_464
timestamp 1
transform -1 0 7912 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_358
timestamp 1
transform 1 0 104052 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_123
timestamp 1
transform -1 0 110860 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_240
timestamp 1
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_465
timestamp 1
transform -1 0 7912 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_359
timestamp 1
transform 1 0 104052 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_124
timestamp 1
transform -1 0 110860 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_241
timestamp 1
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_466
timestamp 1
transform -1 0 7912 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_360
timestamp 1
transform 1 0 104052 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_125
timestamp 1
transform -1 0 110860 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_242
timestamp 1
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_467
timestamp 1
transform -1 0 7912 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_361
timestamp 1
transform 1 0 104052 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_126
timestamp 1
transform -1 0 110860 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_243
timestamp 1
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_468
timestamp 1
transform -1 0 7912 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_362
timestamp 1
transform 1 0 104052 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_127
timestamp 1
transform -1 0 110860 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_244
timestamp 1
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_10
timestamp 1
transform -1 0 110860 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_245
timestamp 1
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_11
timestamp 1
transform -1 0 110860 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_246
timestamp 1
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_12
timestamp 1
transform -1 0 110860 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_247
timestamp 1
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_13
timestamp 1
transform -1 0 110860 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_248
timestamp 1
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_14
timestamp 1
transform -1 0 110860 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_249
timestamp 1
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_15
timestamp 1
transform -1 0 110860 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_250
timestamp 1
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_16
timestamp 1
transform -1 0 110860 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Left_251
timestamp 1
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Right_17
timestamp 1
transform -1 0 110860 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Left_252
timestamp 1
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Right_18
timestamp 1
transform -1 0 110860 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Left_253
timestamp 1
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Right_19
timestamp 1
transform -1 0 110860 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Left_254
timestamp 1
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Right_20
timestamp 1
transform -1 0 110860 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_470
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_471
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_472
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_473
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_474
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_475
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_476
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_477
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_478
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_479
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_480
timestamp 1
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_481
timestamp 1
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_482
timestamp 1
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_483
timestamp 1
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_484
timestamp 1
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_485
timestamp 1
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_486
timestamp 1
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_487
timestamp 1
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_488
timestamp 1
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_489
timestamp 1
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_490
timestamp 1
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_491
timestamp 1
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_492
timestamp 1
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_493
timestamp 1
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_494
timestamp 1
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_495
timestamp 1
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_496
timestamp 1
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_497
timestamp 1
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_498
timestamp 1
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_499
timestamp 1
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_500
timestamp 1
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_501
timestamp 1
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_502
timestamp 1
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_503
timestamp 1
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_504
timestamp 1
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_505
timestamp 1
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_506
timestamp 1
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_507
timestamp 1
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_508
timestamp 1
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_509
timestamp 1
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_510
timestamp 1
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_511
timestamp 1
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_512
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_513
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_514
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_515
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_516
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_517
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_518
timestamp 1
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_519
timestamp 1
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_520
timestamp 1
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_521
timestamp 1
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_522
timestamp 1
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_523
timestamp 1
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_524
timestamp 1
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_525
timestamp 1
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_526
timestamp 1
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_527
timestamp 1
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_528
timestamp 1
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_529
timestamp 1
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_530
timestamp 1
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_531
timestamp 1
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_532
timestamp 1
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_533
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_534
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_535
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_536
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_537
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_538
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_539
timestamp 1
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_540
timestamp 1
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_541
timestamp 1
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_542
timestamp 1
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_543
timestamp 1
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_544
timestamp 1
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_545
timestamp 1
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_546
timestamp 1
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_547
timestamp 1
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_548
timestamp 1
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_549
timestamp 1
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_550
timestamp 1
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_551
timestamp 1
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_552
timestamp 1
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_553
timestamp 1
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_554
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_555
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_556
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_557
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_558
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_559
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_560
timestamp 1
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_561
timestamp 1
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_562
timestamp 1
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_563
timestamp 1
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_564
timestamp 1
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_565
timestamp 1
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_566
timestamp 1
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_567
timestamp 1
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_568
timestamp 1
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_569
timestamp 1
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_570
timestamp 1
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_571
timestamp 1
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_572
timestamp 1
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_573
timestamp 1
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_574
timestamp 1
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_575
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_576
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_577
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_578
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_579
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_580
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_581
timestamp 1
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_582
timestamp 1
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_583
timestamp 1
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_584
timestamp 1
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_585
timestamp 1
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_586
timestamp 1
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_587
timestamp 1
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_588
timestamp 1
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_589
timestamp 1
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_590
timestamp 1
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_591
timestamp 1
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_592
timestamp 1
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_593
timestamp 1
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_594
timestamp 1
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_595
timestamp 1
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_596
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_597
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_598
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_599
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_600
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_601
timestamp 1
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_602
timestamp 1
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_603
timestamp 1
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_604
timestamp 1
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_605
timestamp 1
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_606
timestamp 1
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_607
timestamp 1
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_608
timestamp 1
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_609
timestamp 1
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_610
timestamp 1
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_611
timestamp 1
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_612
timestamp 1
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_613
timestamp 1
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_614
timestamp 1
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_615
timestamp 1
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_616
timestamp 1
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_617
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_618
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_619
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_620
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_621
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_622
timestamp 1
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_623
timestamp 1
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_624
timestamp 1
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_625
timestamp 1
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_626
timestamp 1
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_627
timestamp 1
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_628
timestamp 1
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_629
timestamp 1
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_630
timestamp 1
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_631
timestamp 1
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_632
timestamp 1
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_633
timestamp 1
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_634
timestamp 1
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_635
timestamp 1
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_636
timestamp 1
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_637
timestamp 1
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_638
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_639
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_640
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_641
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_642
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_643
timestamp 1
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_644
timestamp 1
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_645
timestamp 1
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_646
timestamp 1
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_647
timestamp 1
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_648
timestamp 1
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_649
timestamp 1
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_650
timestamp 1
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_651
timestamp 1
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_652
timestamp 1
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_653
timestamp 1
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_654
timestamp 1
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_655
timestamp 1
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_656
timestamp 1
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_657
timestamp 1
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_658
timestamp 1
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_659
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_660
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_661
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_662
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_663
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_664
timestamp 1
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_665
timestamp 1
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_666
timestamp 1
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_667
timestamp 1
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_668
timestamp 1
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_669
timestamp 1
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_670
timestamp 1
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_671
timestamp 1
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_672
timestamp 1
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_673
timestamp 1
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_674
timestamp 1
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_675
timestamp 1
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_676
timestamp 1
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_677
timestamp 1
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_678
timestamp 1
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_679
timestamp 1
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_680
timestamp 1
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_681
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_682
timestamp 1
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_683
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_684
timestamp 1
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_685
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_686
timestamp 1
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_687
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_688
timestamp 1
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_689
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_690
timestamp 1
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_691
timestamp 1
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_692
timestamp 1
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_693
timestamp 1
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_694
timestamp 1
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_695
timestamp 1
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_696
timestamp 1
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_697
timestamp 1
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_698
timestamp 1
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_699
timestamp 1
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_700
timestamp 1
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_701
timestamp 1
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_702
timestamp 1
transform 1 0 60352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_703
timestamp 1
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_704
timestamp 1
transform 1 0 65504 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_705
timestamp 1
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_706
timestamp 1
transform 1 0 70656 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_707
timestamp 1
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_708
timestamp 1
transform 1 0 75808 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_709
timestamp 1
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_710
timestamp 1
transform 1 0 80960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_711
timestamp 1
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_712
timestamp 1
transform 1 0 86112 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_713
timestamp 1
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_714
timestamp 1
transform 1 0 91264 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_715
timestamp 1
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_716
timestamp 1
transform 1 0 96416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_717
timestamp 1
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_718
timestamp 1
transform 1 0 101568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_719
timestamp 1
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_720
timestamp 1
transform 1 0 106720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_721
timestamp 1
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_1101
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_1102
timestamp 1
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_1_722
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_1103
timestamp 1
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_723
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_1104
timestamp 1
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_1_724
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_1105
timestamp 1
transform 1 0 109204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_725
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_1106
timestamp 1
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_1_726
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_2_1107
timestamp 1
transform 1 0 109204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_727
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_1108
timestamp 1
transform 1 0 106628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_1_728
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_2_1109
timestamp 1
transform 1 0 109204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_729
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_1110
timestamp 1
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_1_730
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_2_1111
timestamp 1
transform 1 0 109204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_731
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_1112
timestamp 1
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_1_732
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_2_1113
timestamp 1
transform 1 0 109204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_733
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_1114
timestamp 1
transform 1 0 106628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_1_734
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_2_1115
timestamp 1
transform 1 0 109204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_735
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_1116
timestamp 1
transform 1 0 106628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_1_736
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_2_1117
timestamp 1
transform 1 0 109204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_737
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_1118
timestamp 1
transform 1 0 106628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_1_738
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_2_1119
timestamp 1
transform 1 0 109204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_739
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_1120
timestamp 1
transform 1 0 106628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_1_740
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_2_1121
timestamp 1
transform 1 0 109204 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_741
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_1122
timestamp 1
transform 1 0 106628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_1_742
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_2_1123
timestamp 1
transform 1 0 109204 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_743
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_1124
timestamp 1
transform 1 0 106628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_1_744
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_2_1125
timestamp 1
transform 1 0 109204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_745
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_1126
timestamp 1
transform 1 0 106628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_1_746
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_2_1127
timestamp 1
transform 1 0 109204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_747
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_1128
timestamp 1
transform 1 0 106628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_1_748
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_2_1129
timestamp 1
transform 1 0 109204 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_749
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_1130
timestamp 1
transform 1 0 106628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_1_750
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_2_1131
timestamp 1
transform 1 0 109204 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_751
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_1132
timestamp 1
transform 1 0 106628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_1_752
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_2_1133
timestamp 1
transform 1 0 109204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_753
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_1134
timestamp 1
transform 1 0 106628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_1_754
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_2_1135
timestamp 1
transform 1 0 109204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_755
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_1136
timestamp 1
transform 1 0 106628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_1_756
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_2_1137
timestamp 1
transform 1 0 109204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_757
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_1138
timestamp 1
transform 1 0 106628 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_1_758
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_2_1139
timestamp 1
transform 1 0 109204 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_759
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_1140
timestamp 1
transform 1 0 106628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1_760
timestamp 1
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_2_1141
timestamp 1
transform 1 0 109204 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_761
timestamp 1
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_1142
timestamp 1
transform 1 0 106628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1_762
timestamp 1
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_2_1143
timestamp 1
transform 1 0 109204 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_763
timestamp 1
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_1144
timestamp 1
transform 1 0 106628 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1_764
timestamp 1
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_2_1145
timestamp 1
transform 1 0 109204 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_765
timestamp 1
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_1146
timestamp 1
transform 1 0 106628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1_766
timestamp 1
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_2_1147
timestamp 1
transform 1 0 109204 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_767
timestamp 1
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_1148
timestamp 1
transform 1 0 106628 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1_768
timestamp 1
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_2_1149
timestamp 1
transform 1 0 109204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_769
timestamp 1
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_1150
timestamp 1
transform 1 0 106628 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1_770
timestamp 1
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_2_1151
timestamp 1
transform 1 0 109204 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_771
timestamp 1
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_1152
timestamp 1
transform 1 0 106628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1_772
timestamp 1
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_2_1153
timestamp 1
transform 1 0 109204 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_773
timestamp 1
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_1154
timestamp 1
transform 1 0 106628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1_774
timestamp 1
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_2_1155
timestamp 1
transform 1 0 109204 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_775
timestamp 1
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_1156
timestamp 1
transform 1 0 106628 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1_776
timestamp 1
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_2_1157
timestamp 1
transform 1 0 109204 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_777
timestamp 1
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_1158
timestamp 1
transform 1 0 106628 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1_778
timestamp 1
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_2_1159
timestamp 1
transform 1 0 109204 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_779
timestamp 1
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_1160
timestamp 1
transform 1 0 106628 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1_780
timestamp 1
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_2_1161
timestamp 1
transform 1 0 109204 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_781
timestamp 1
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_1162
timestamp 1
transform 1 0 106628 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1_782
timestamp 1
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_2_1163
timestamp 1
transform 1 0 109204 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_783
timestamp 1
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_1164
timestamp 1
transform 1 0 106628 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1_784
timestamp 1
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_2_1165
timestamp 1
transform 1 0 109204 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_785
timestamp 1
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_1166
timestamp 1
transform 1 0 106628 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1_786
timestamp 1
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_2_1167
timestamp 1
transform 1 0 109204 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_787
timestamp 1
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_1168
timestamp 1
transform 1 0 106628 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1_788
timestamp 1
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_2_1169
timestamp 1
transform 1 0 109204 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_789
timestamp 1
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_1170
timestamp 1
transform 1 0 106628 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1_790
timestamp 1
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_2_1171
timestamp 1
transform 1 0 109204 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_791
timestamp 1
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_1172
timestamp 1
transform 1 0 106628 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1_792
timestamp 1
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_2_1173
timestamp 1
transform 1 0 109204 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_793
timestamp 1
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_1174
timestamp 1
transform 1 0 106628 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1_794
timestamp 1
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_2_1175
timestamp 1
transform 1 0 109204 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_795
timestamp 1
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_1176
timestamp 1
transform 1 0 106628 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1_796
timestamp 1
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_2_1177
timestamp 1
transform 1 0 109204 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_797
timestamp 1
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_1178
timestamp 1
transform 1 0 106628 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1_798
timestamp 1
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_2_1179
timestamp 1
transform 1 0 109204 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_799
timestamp 1
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_1180
timestamp 1
transform 1 0 106628 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1_800
timestamp 1
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_2_1181
timestamp 1
transform 1 0 109204 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_801
timestamp 1
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_1182
timestamp 1
transform 1 0 106628 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1_802
timestamp 1
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_2_1183
timestamp 1
transform 1 0 109204 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_803
timestamp 1
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_1184
timestamp 1
transform 1 0 106628 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1_804
timestamp 1
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_2_1185
timestamp 1
transform 1 0 109204 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_805
timestamp 1
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_1186
timestamp 1
transform 1 0 106628 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1_806
timestamp 1
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_2_1187
timestamp 1
transform 1 0 109204 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_807
timestamp 1
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_1188
timestamp 1
transform 1 0 106628 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1_808
timestamp 1
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_2_1189
timestamp 1
transform 1 0 109204 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_809
timestamp 1
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_1190
timestamp 1
transform 1 0 106628 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1_810
timestamp 1
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_2_1191
timestamp 1
transform 1 0 109204 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_811
timestamp 1
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_1192
timestamp 1
transform 1 0 106628 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1_812
timestamp 1
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_2_1193
timestamp 1
transform 1 0 109204 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_813
timestamp 1
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_1194
timestamp 1
transform 1 0 106628 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1_814
timestamp 1
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_2_1195
timestamp 1
transform 1 0 109204 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_815
timestamp 1
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_1196
timestamp 1
transform 1 0 106628 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1_816
timestamp 1
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_2_1197
timestamp 1
transform 1 0 109204 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_817
timestamp 1
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_1198
timestamp 1
transform 1 0 106628 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1_818
timestamp 1
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_2_1199
timestamp 1
transform 1 0 109204 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_819
timestamp 1
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_1200
timestamp 1
transform 1 0 106628 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1_820
timestamp 1
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_2_1201
timestamp 1
transform 1 0 109204 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_821
timestamp 1
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_1202
timestamp 1
transform 1 0 106628 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1_822
timestamp 1
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_2_1203
timestamp 1
transform 1 0 109204 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_823
timestamp 1
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_1204
timestamp 1
transform 1 0 106628 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1_824
timestamp 1
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_2_1205
timestamp 1
transform 1 0 109204 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_825
timestamp 1
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_1206
timestamp 1
transform 1 0 106628 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1_826
timestamp 1
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_2_1207
timestamp 1
transform 1 0 109204 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_827
timestamp 1
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_1208
timestamp 1
transform 1 0 106628 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_828
timestamp 1
transform 1 0 3680 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_829
timestamp 1
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_830
timestamp 1
transform 1 0 8832 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_831
timestamp 1
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_832
timestamp 1
transform 1 0 13984 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_833
timestamp 1
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_834
timestamp 1
transform 1 0 19136 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_835
timestamp 1
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_836
timestamp 1
transform 1 0 24288 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_837
timestamp 1
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_838
timestamp 1
transform 1 0 29440 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_839
timestamp 1
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_840
timestamp 1
transform 1 0 34592 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_841
timestamp 1
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_842
timestamp 1
transform 1 0 39744 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_843
timestamp 1
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_844
timestamp 1
transform 1 0 44896 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_845
timestamp 1
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_846
timestamp 1
transform 1 0 50048 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_847
timestamp 1
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_848
timestamp 1
transform 1 0 55200 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_849
timestamp 1
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_850
timestamp 1
transform 1 0 60352 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_851
timestamp 1
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_852
timestamp 1
transform 1 0 65504 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_853
timestamp 1
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_854
timestamp 1
transform 1 0 70656 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_855
timestamp 1
transform 1 0 73232 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_856
timestamp 1
transform 1 0 75808 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_857
timestamp 1
transform 1 0 78384 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_858
timestamp 1
transform 1 0 80960 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_859
timestamp 1
transform 1 0 83536 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_860
timestamp 1
transform 1 0 86112 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_861
timestamp 1
transform 1 0 88688 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_862
timestamp 1
transform 1 0 91264 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_863
timestamp 1
transform 1 0 93840 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_864
timestamp 1
transform 1 0 96416 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_865
timestamp 1
transform 1 0 98992 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_866
timestamp 1
transform 1 0 101568 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_867
timestamp 1
transform 1 0 104144 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_868
timestamp 1
transform 1 0 106720 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_869
timestamp 1
transform 1 0 109296 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_870
timestamp 1
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_871
timestamp 1
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_872
timestamp 1
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_873
timestamp 1
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_874
timestamp 1
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_875
timestamp 1
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_876
timestamp 1
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_877
timestamp 1
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_878
timestamp 1
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_879
timestamp 1
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_880
timestamp 1
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_881
timestamp 1
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_882
timestamp 1
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_883
timestamp 1
transform 1 0 70656 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_884
timestamp 1
transform 1 0 75808 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_885
timestamp 1
transform 1 0 80960 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_886
timestamp 1
transform 1 0 86112 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_887
timestamp 1
transform 1 0 91264 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_888
timestamp 1
transform 1 0 96416 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_889
timestamp 1
transform 1 0 101568 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_890
timestamp 1
transform 1 0 106720 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_891
timestamp 1
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_892
timestamp 1
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_893
timestamp 1
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_894
timestamp 1
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_895
timestamp 1
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_896
timestamp 1
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_897
timestamp 1
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_898
timestamp 1
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_899
timestamp 1
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_900
timestamp 1
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_901
timestamp 1
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_902
timestamp 1
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_903
timestamp 1
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_904
timestamp 1
transform 1 0 73232 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_905
timestamp 1
transform 1 0 78384 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_906
timestamp 1
transform 1 0 83536 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_907
timestamp 1
transform 1 0 88688 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_908
timestamp 1
transform 1 0 93840 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_909
timestamp 1
transform 1 0 98992 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_910
timestamp 1
transform 1 0 104144 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_911
timestamp 1
transform 1 0 109296 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_912
timestamp 1
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_913
timestamp 1
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_914
timestamp 1
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_915
timestamp 1
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_916
timestamp 1
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_917
timestamp 1
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_918
timestamp 1
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_919
timestamp 1
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_920
timestamp 1
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_921
timestamp 1
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_922
timestamp 1
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_923
timestamp 1
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_924
timestamp 1
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_925
timestamp 1
transform 1 0 70656 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_926
timestamp 1
transform 1 0 75808 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_927
timestamp 1
transform 1 0 80960 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_928
timestamp 1
transform 1 0 86112 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_929
timestamp 1
transform 1 0 91264 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_930
timestamp 1
transform 1 0 96416 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_931
timestamp 1
transform 1 0 101568 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_932
timestamp 1
transform 1 0 106720 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_933
timestamp 1
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_934
timestamp 1
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_935
timestamp 1
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_936
timestamp 1
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_937
timestamp 1
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_938
timestamp 1
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_939
timestamp 1
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_940
timestamp 1
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_941
timestamp 1
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_942
timestamp 1
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_943
timestamp 1
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_944
timestamp 1
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_945
timestamp 1
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_946
timestamp 1
transform 1 0 73232 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_947
timestamp 1
transform 1 0 78384 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_948
timestamp 1
transform 1 0 83536 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_949
timestamp 1
transform 1 0 88688 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_950
timestamp 1
transform 1 0 93840 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_951
timestamp 1
transform 1 0 98992 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_952
timestamp 1
transform 1 0 104144 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_953
timestamp 1
transform 1 0 109296 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_954
timestamp 1
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_955
timestamp 1
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_956
timestamp 1
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_957
timestamp 1
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_958
timestamp 1
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_959
timestamp 1
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_960
timestamp 1
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_961
timestamp 1
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_962
timestamp 1
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_963
timestamp 1
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_964
timestamp 1
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_965
timestamp 1
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_966
timestamp 1
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_967
timestamp 1
transform 1 0 70656 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_968
timestamp 1
transform 1 0 75808 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_969
timestamp 1
transform 1 0 80960 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_970
timestamp 1
transform 1 0 86112 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_971
timestamp 1
transform 1 0 91264 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_972
timestamp 1
transform 1 0 96416 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_973
timestamp 1
transform 1 0 101568 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_974
timestamp 1
transform 1 0 106720 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_975
timestamp 1
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_976
timestamp 1
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_977
timestamp 1
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_978
timestamp 1
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_979
timestamp 1
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_980
timestamp 1
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_981
timestamp 1
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_982
timestamp 1
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_983
timestamp 1
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_984
timestamp 1
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_985
timestamp 1
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_986
timestamp 1
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_987
timestamp 1
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_988
timestamp 1
transform 1 0 73232 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_989
timestamp 1
transform 1 0 78384 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_990
timestamp 1
transform 1 0 83536 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_991
timestamp 1
transform 1 0 88688 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_992
timestamp 1
transform 1 0 93840 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_993
timestamp 1
transform 1 0 98992 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_994
timestamp 1
transform 1 0 104144 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_995
timestamp 1
transform 1 0 109296 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_996
timestamp 1
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_997
timestamp 1
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_998
timestamp 1
transform 1 0 13984 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_999
timestamp 1
transform 1 0 19136 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1000
timestamp 1
transform 1 0 24288 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1001
timestamp 1
transform 1 0 29440 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1002
timestamp 1
transform 1 0 34592 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1003
timestamp 1
transform 1 0 39744 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1004
timestamp 1
transform 1 0 44896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1005
timestamp 1
transform 1 0 50048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1006
timestamp 1
transform 1 0 55200 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1007
timestamp 1
transform 1 0 60352 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1008
timestamp 1
transform 1 0 65504 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1009
timestamp 1
transform 1 0 70656 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1010
timestamp 1
transform 1 0 75808 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1011
timestamp 1
transform 1 0 80960 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1012
timestamp 1
transform 1 0 86112 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1013
timestamp 1
transform 1 0 91264 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1014
timestamp 1
transform 1 0 96416 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1015
timestamp 1
transform 1 0 101568 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1016
timestamp 1
transform 1 0 106720 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1017
timestamp 1
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1018
timestamp 1
transform 1 0 11408 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1019
timestamp 1
transform 1 0 16560 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1020
timestamp 1
transform 1 0 21712 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1021
timestamp 1
transform 1 0 26864 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1022
timestamp 1
transform 1 0 32016 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1023
timestamp 1
transform 1 0 37168 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1024
timestamp 1
transform 1 0 42320 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1025
timestamp 1
transform 1 0 47472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1026
timestamp 1
transform 1 0 52624 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1027
timestamp 1
transform 1 0 57776 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1028
timestamp 1
transform 1 0 62928 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1029
timestamp 1
transform 1 0 68080 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1030
timestamp 1
transform 1 0 73232 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1031
timestamp 1
transform 1 0 78384 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1032
timestamp 1
transform 1 0 83536 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1033
timestamp 1
transform 1 0 88688 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1034
timestamp 1
transform 1 0 93840 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1035
timestamp 1
transform 1 0 98992 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1036
timestamp 1
transform 1 0 104144 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_1037
timestamp 1
transform 1 0 109296 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1038
timestamp 1
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1039
timestamp 1
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1040
timestamp 1
transform 1 0 13984 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1041
timestamp 1
transform 1 0 19136 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1042
timestamp 1
transform 1 0 24288 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1043
timestamp 1
transform 1 0 29440 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1044
timestamp 1
transform 1 0 34592 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1045
timestamp 1
transform 1 0 39744 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1046
timestamp 1
transform 1 0 44896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1047
timestamp 1
transform 1 0 50048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1048
timestamp 1
transform 1 0 55200 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1049
timestamp 1
transform 1 0 60352 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1050
timestamp 1
transform 1 0 65504 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1051
timestamp 1
transform 1 0 70656 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1052
timestamp 1
transform 1 0 75808 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1053
timestamp 1
transform 1 0 80960 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1054
timestamp 1
transform 1 0 86112 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1055
timestamp 1
transform 1 0 91264 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1056
timestamp 1
transform 1 0 96416 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1057
timestamp 1
transform 1 0 101568 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1058
timestamp 1
transform 1 0 106720 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1059
timestamp 1
transform 1 0 3680 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1060
timestamp 1
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1061
timestamp 1
transform 1 0 8832 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1062
timestamp 1
transform 1 0 11408 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1063
timestamp 1
transform 1 0 13984 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1064
timestamp 1
transform 1 0 16560 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1065
timestamp 1
transform 1 0 19136 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1066
timestamp 1
transform 1 0 21712 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1067
timestamp 1
transform 1 0 24288 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1068
timestamp 1
transform 1 0 26864 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1069
timestamp 1
transform 1 0 29440 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1070
timestamp 1
transform 1 0 32016 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1071
timestamp 1
transform 1 0 34592 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1072
timestamp 1
transform 1 0 37168 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1073
timestamp 1
transform 1 0 39744 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1074
timestamp 1
transform 1 0 42320 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1075
timestamp 1
transform 1 0 44896 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1076
timestamp 1
transform 1 0 47472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1077
timestamp 1
transform 1 0 50048 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1078
timestamp 1
transform 1 0 52624 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1079
timestamp 1
transform 1 0 55200 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1080
timestamp 1
transform 1 0 57776 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1081
timestamp 1
transform 1 0 60352 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1082
timestamp 1
transform 1 0 62928 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1083
timestamp 1
transform 1 0 65504 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1084
timestamp 1
transform 1 0 68080 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1085
timestamp 1
transform 1 0 70656 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1086
timestamp 1
transform 1 0 73232 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1087
timestamp 1
transform 1 0 75808 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1088
timestamp 1
transform 1 0 78384 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1089
timestamp 1
transform 1 0 80960 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1090
timestamp 1
transform 1 0 83536 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1091
timestamp 1
transform 1 0 86112 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1092
timestamp 1
transform 1 0 88688 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1093
timestamp 1
transform 1 0 91264 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1094
timestamp 1
transform 1 0 93840 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1095
timestamp 1
transform 1 0 96416 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1096
timestamp 1
transform 1 0 98992 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1097
timestamp 1
transform 1 0 101568 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1098
timestamp 1
transform 1 0 104144 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1099
timestamp 1
transform 1 0 106720 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1100
timestamp 1
transform 1 0 109296 0 -1 71808
box -38 -48 130 592
<< labels >>
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 addr0[0]
port 0 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 addr0[1]
port 1 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 addr0[2]
port 2 nsew signal input
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 addr0[3]
port 3 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 addr0[4]
port 4 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 addr0[5]
port 5 nsew signal input
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 addr0[6]
port 6 nsew signal input
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 addr0[7]
port 7 nsew signal input
flabel metal3 s 111200 10208 112000 10328 0 FreeSans 480 0 0 0 clk
port 8 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 csb0
port 9 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 din0[0]
port 10 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 din0[10]
port 11 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 din0[11]
port 12 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 din0[12]
port 13 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 din0[13]
port 14 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 din0[14]
port 15 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 din0[15]
port 16 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 din0[1]
port 17 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 din0[2]
port 18 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 din0[3]
port 19 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 din0[4]
port 20 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 din0[5]
port 21 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 din0[6]
port 22 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 din0[7]
port 23 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 din0[8]
port 24 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 din0[9]
port 25 nsew signal input
flabel metal3 s 111200 31288 112000 31408 0 FreeSans 480 0 0 0 rst
port 26 nsew signal input
flabel metal2 s 44454 73200 44510 74000 0 FreeSans 224 90 0 0 sine_out[0]
port 27 nsew signal output
flabel metal2 s 65706 73200 65762 74000 0 FreeSans 224 90 0 0 sine_out[10]
port 28 nsew signal output
flabel metal2 s 67638 73200 67694 74000 0 FreeSans 224 90 0 0 sine_out[11]
port 29 nsew signal output
flabel metal2 s 69570 73200 69626 74000 0 FreeSans 224 90 0 0 sine_out[12]
port 30 nsew signal output
flabel metal2 s 71502 73200 71558 74000 0 FreeSans 224 90 0 0 sine_out[13]
port 31 nsew signal output
flabel metal2 s 74078 73200 74134 74000 0 FreeSans 224 90 0 0 sine_out[14]
port 32 nsew signal output
flabel metal2 s 77298 73200 77354 74000 0 FreeSans 224 90 0 0 sine_out[15]
port 33 nsew signal output
flabel metal2 s 47030 73200 47086 74000 0 FreeSans 224 90 0 0 sine_out[1]
port 34 nsew signal output
flabel metal2 s 49606 73200 49662 74000 0 FreeSans 224 90 0 0 sine_out[2]
port 35 nsew signal output
flabel metal2 s 51538 73200 51594 74000 0 FreeSans 224 90 0 0 sine_out[3]
port 36 nsew signal output
flabel metal2 s 53470 73200 53526 74000 0 FreeSans 224 90 0 0 sine_out[4]
port 37 nsew signal output
flabel metal2 s 55402 73200 55458 74000 0 FreeSans 224 90 0 0 sine_out[5]
port 38 nsew signal output
flabel metal2 s 57334 73200 57390 74000 0 FreeSans 224 90 0 0 sine_out[6]
port 39 nsew signal output
flabel metal2 s 59266 73200 59322 74000 0 FreeSans 224 90 0 0 sine_out[7]
port 40 nsew signal output
flabel metal2 s 61198 73200 61254 74000 0 FreeSans 224 90 0 0 sine_out[8]
port 41 nsew signal output
flabel metal2 s 63130 73200 63186 74000 0 FreeSans 224 90 0 0 sine_out[9]
port 42 nsew signal output
flabel metal4 s 4208 2128 4528 71856 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 34928 2128 35248 7880 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 34928 65650 35248 71856 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 65648 2128 65968 8064 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 65648 65776 65968 71856 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 96368 2128 96688 8064 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 96368 65650 96688 71856 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 1056 5346 110908 5666 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 1056 35982 110908 36302 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 1056 66618 110908 66938 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 107020 7024 107340 66416 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 4868 2128 5188 71856 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 8064 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 35588 65650 35908 71856 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 66308 2128 66628 8064 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 66308 65650 66628 71856 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 97028 2128 97348 8064 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 97028 65650 97348 71856 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal5 s 1056 6006 110908 6326 0 FreeSans 2560 0 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal5 s 1056 36642 110908 36962 0 FreeSans 2560 0 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal5 s 1056 67278 110908 67598 0 FreeSans 2560 0 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 107756 7024 108076 66416 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
rlabel via4 101806 36142 101806 36142 0 vccd1
rlabel via4 101110 36802 101110 36802 0 vssd1
rlabel metal1 104558 55930 104558 55930 0 _000_
rlabel metal1 104512 53754 104512 53754 0 _001_
rlabel metal1 104558 41242 104558 41242 0 _002_
rlabel metal1 105938 31994 105938 31994 0 _003_
rlabel metal1 105432 30090 105432 30090 0 _004_
rlabel metal1 104512 27098 104512 27098 0 _005_
rlabel metal1 104742 23562 104742 23562 0 _006_
rlabel metal2 104374 20060 104374 20060 0 _007_
rlabel metal1 58420 65926 58420 65926 0 _008_
rlabel metal1 60398 67320 60398 67320 0 _009_
rlabel metal1 62606 65926 62606 65926 0 _010_
rlabel metal2 64906 66368 64906 66368 0 _011_
rlabel metal1 66240 66198 66240 66198 0 _012_
rlabel metal1 67758 66198 67758 66198 0 _013_
rlabel metal2 69598 66708 69598 66708 0 _014_
rlabel metal2 71438 66708 71438 66708 0 _015_
rlabel metal2 73462 66368 73462 66368 0 _016_
rlabel metal1 75900 66198 75900 66198 0 _017_
rlabel metal2 102994 61778 102994 61778 0 _018_
rlabel metal1 104788 54298 104788 54298 0 _019_
rlabel metal1 104788 43690 104788 43690 0 _020_
rlabel metal1 104512 36550 104512 36550 0 _021_
rlabel metal2 104466 34136 104466 34136 0 _022_
rlabel metal1 104604 31926 104604 31926 0 _023_
rlabel metal1 104689 25942 104689 25942 0 _024_
rlabel metal2 104926 22984 104926 22984 0 _025_
rlabel metal2 44758 66980 44758 66980 0 _026_
rlabel metal2 50554 66436 50554 66436 0 _027_
rlabel metal1 52486 66232 52486 66232 0 _028_
rlabel metal1 54004 66198 54004 66198 0 _029_
rlabel metal1 55522 66198 55522 66198 0 _030_
rlabel metal2 58006 66470 58006 66470 0 _031_
rlabel metal1 104926 24378 104926 24378 0 _032_
rlabel metal1 104328 41106 104328 41106 0 _033_
rlabel metal1 105340 30158 105340 30158 0 _034_
rlabel metal1 105156 26962 105156 26962 0 _035_
rlabel metal1 104696 24174 104696 24174 0 _036_
rlabel metal2 104742 22797 104742 22797 0 _037_
rlabel metal1 104650 23698 104650 23698 0 _038_
rlabel metal2 23506 8551 23506 8551 0 addr0[0]
rlabel metal2 24518 3831 24518 3831 0 addr0[1]
rlabel metal3 9476 34000 9476 34000 0 addr0[2]
rlabel metal3 2039 35428 2039 35428 0 addr0[3]
rlabel metal3 9476 36742 9476 36742 0 addr0[4]
rlabel metal3 1855 38148 1855 38148 0 addr0[5]
rlabel metal3 9476 39516 9476 39516 0 addr0[6]
rlabel metal3 3787 41548 3787 41548 0 addr0[7]
rlabel metal1 82110 65960 82110 65960 0 clk
rlabel metal1 57730 66096 57730 66096 0 clknet_0_clk
rlabel metal1 44298 67354 44298 67354 0 clknet_1_0__leaf_clk
rlabel metal4 95890 63779 95890 63779 0 clknet_1_1__leaf_clk
rlabel metal3 2039 15708 2039 15708 0 csb0
rlabel via3 25829 8092 25829 8092 0 din0[0]
rlabel metal2 37398 3831 37398 3831 0 din0[10]
rlabel via3 38709 8092 38709 8092 0 din0[11]
rlabel metal2 39974 3831 39974 3831 0 din0[12]
rlabel metal2 41262 3831 41262 3831 0 din0[13]
rlabel via2 42182 7531 42182 7531 0 din0[14]
rlabel metal2 43194 3831 43194 3831 0 din0[15]
rlabel metal2 27094 3831 27094 3831 0 din0[1]
rlabel metal2 28382 3831 28382 3831 0 din0[2]
rlabel metal3 29187 8092 29187 8092 0 din0[3]
rlabel metal2 30314 3831 30314 3831 0 din0[4]
rlabel via3 31624 9724 31624 9724 0 din0[5]
rlabel via3 32867 8092 32867 8092 0 din0[6]
rlabel metal2 34178 3831 34178 3831 0 din0[7]
rlabel metal2 35282 7803 35282 7803 0 din0[8]
rlabel via2 36386 7531 36386 7531 0 din0[9]
rlabel metal2 110354 32198 110354 32198 0 net1
rlabel metal2 49542 69462 49542 69462 0 net10
rlabel metal1 51566 67354 51566 67354 0 net11
rlabel metal1 53498 66810 53498 66810 0 net12
rlabel metal1 55430 67354 55430 67354 0 net13
rlabel metal1 57316 67354 57316 67354 0 net14
rlabel metal2 59662 69462 59662 69462 0 net15
rlabel metal1 61548 67354 61548 67354 0 net16
rlabel metal1 63204 71570 63204 71570 0 net17
rlabel metal1 58098 66164 58098 66164 0 net18
rlabel metal1 72542 66130 72542 66130 0 net19
rlabel metal2 45126 69360 45126 69360 0 net2
rlabel metal2 102902 59534 102902 59534 0 net20
rlabel metal3 102279 59738 102279 59738 0 net21
rlabel metal2 104558 56202 104558 56202 0 net22
rlabel metal1 105202 30226 105202 30226 0 net23
rlabel metal2 104742 19788 104742 19788 0 net24
rlabel metal2 105662 32538 105662 32538 0 net25
rlabel metal1 65642 71570 65642 71570 0 net3
rlabel metal1 67574 71570 67574 71570 0 net4
rlabel metal2 69966 69462 69966 69462 0 net5
rlabel metal1 71852 67354 71852 67354 0 net6
rlabel metal1 73876 66470 73876 66470 0 net7
rlabel metal1 76774 71570 76774 71570 0 net8
rlabel metal2 47334 69360 47334 69360 0 net9
rlabel metal2 110538 31569 110538 31569 0 rst
rlabel metal1 44574 71706 44574 71706 0 sine_out[0]
rlabel metal1 65872 71706 65872 71706 0 sine_out[10]
rlabel metal1 67804 71706 67804 71706 0 sine_out[11]
rlabel metal1 69690 71706 69690 71706 0 sine_out[12]
rlabel metal1 71622 71706 71622 71706 0 sine_out[13]
rlabel metal1 74244 71706 74244 71706 0 sine_out[14]
rlabel metal1 77464 71706 77464 71706 0 sine_out[15]
rlabel metal1 47150 71706 47150 71706 0 sine_out[1]
rlabel metal1 49772 71706 49772 71706 0 sine_out[2]
rlabel metal1 51704 71706 51704 71706 0 sine_out[3]
rlabel metal1 53636 71706 53636 71706 0 sine_out[4]
rlabel metal1 55568 71706 55568 71706 0 sine_out[5]
rlabel metal1 57500 71706 57500 71706 0 sine_out[6]
rlabel metal1 59386 71706 59386 71706 0 sine_out[7]
rlabel metal1 61318 71706 61318 71706 0 sine_out[8]
rlabel metal1 63296 71706 63296 71706 0 sine_out[9]
rlabel metal4 36107 63915 36107 63915 0 sine_out_temp\[0\]
rlabel metal4 61088 63983 61088 63983 0 sine_out_temp\[10\]
rlabel metal4 63572 64595 63572 64595 0 sine_out_temp\[11\]
rlabel metal4 66059 63983 66059 63983 0 sine_out_temp\[12\]
rlabel metal4 68540 64527 68540 64527 0 sine_out_temp\[13\]
rlabel metal4 71051 63983 71051 63983 0 sine_out_temp\[14\]
rlabel metal4 73547 63983 73547 63983 0 sine_out_temp\[15\]
rlabel metal4 38603 63779 38603 63779 0 sine_out_temp\[1\]
rlabel metal4 41099 63847 41099 63847 0 sine_out_temp\[2\]
rlabel metal4 43608 63915 43608 63915 0 sine_out_temp\[3\]
rlabel metal3 47909 66300 47909 66300 0 sine_out_temp\[4\]
rlabel metal4 48587 63983 48587 63983 0 sine_out_temp\[5\]
rlabel metal2 55706 66929 55706 66929 0 sine_out_temp\[6\]
rlabel metal2 58190 65501 58190 65501 0 sine_out_temp\[7\]
rlabel metal4 56051 64260 56051 64260 0 sine_out_temp\[8\]
rlabel metal4 58571 63983 58571 63983 0 sine_out_temp\[9\]
rlabel metal4 87342 63915 87342 63915 0 tcout\[0\]
rlabel metal4 86174 63847 86174 63847 0 tcout\[1\]
rlabel metal3 102279 25060 102279 25060 0 tcout\[2\]
rlabel metal3 102279 23360 102279 23360 0 tcout\[3\]
rlabel metal3 102279 22232 102279 22232 0 tcout\[4\]
rlabel metal1 104428 25126 104428 25126 0 tcout\[5\]
rlabel metal1 104282 23766 104282 23766 0 tcout\[6\]
rlabel metal1 104328 19686 104328 19686 0 tcout\[7\]
<< properties >>
string FIXED_BBOX 0 0 112000 74000
<< end >>
