sine_table[1] = {
16'h9127,
16'h901f,
16'h8f1e,
16'h8e25,
16'h8d34,
16'h8c4b,
16'h8b6a,
16'h8a90,
16'h89bf,
16'h88f6,
16'h8835,
16'h877c,
16'h86cc,
16'h8624,
16'h8584,
16'h84ed,
16'h845e,
16'h83d7,
16'h8359,
16'h82e4,
16'h8277,
16'h8212,
16'h81b7,
16'h8164,
16'h8119,
16'h80d8,
16'h809f,
16'h806f,
16'h8047,
16'h8028,
16'h8013,
16'h8005,
16'h8001,
16'h8005,
16'h8013,
16'h8028,
16'h8047,
16'h806f,
16'h809f,
16'h80d8,
16'h8119,
16'h8164,
16'h81b7,
16'h8212,
16'h8277,
16'h82e4,
16'h8359,
16'h83d7,
16'h845e,
16'h84ed,
16'h8584,
16'h8624,
16'h86cc,
16'h877c,
16'h8835,
16'h88f6,
16'h89bf,
16'h8a90,
16'h8b6a,
16'h8c4b,
16'h8d34,
16'h8e25,
16'h8f1e,
16'h901f,
16'h9127,
16'h9237,
16'h934e,
16'h946d,
16'h9593,
16'h96c1,
16'h97f5,
16'h9931,
16'h9a74,
16'h9bbe,
16'h9d0f,
16'h9e66,
16'h9fc4,
16'ha129,
16'ha295,
16'ha406,
16'ha57e,
16'ha6fc,
16'ha881,
16'haa0b,
16'hab9b,
16'had31,
16'haecd,
16'hb06e,
16'hb215,
16'hb3c1,
16'hb572,
16'hb728,
16'hb8e4,
16'hbaa4,
16'hbc69,
16'hbe32,
16'hc000,
16'hc1d3,
16'hc3aa,
16'hc585,
16'hc764,
16'hc946,
16'hcb2d,
16'hcd17,
16'hcf05,
16'hd0f6,
16'hd2ea,
16'hd4e1,
16'hd6db,
16'hd8d8,
16'hdad8,
16'hdcdb,
16'hdedf,
16'he0e6,
16'he2ef,
16'he4fb,
16'he707,
16'he916,
16'heb26,
16'hed38,
16'hef4b,
16'hf15f,
16'hf374,
16'hf58a,
16'hf7a1,
16'hf9b8,
16'hfbd0,
16'hfde8,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000,
16'h0000
};