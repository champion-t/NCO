VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 98.060 BY 108.780 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 95.440 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 95.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 94.060 68.040 98.060 68.640 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 94.060 71.440 98.060 72.040 ;
    END
  END rst
  PIN sine_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 94.060 61.240 98.060 61.840 ;
    END
  END sine_out[0]
  PIN sine_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END sine_out[10]
  PIN sine_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END sine_out[11]
  PIN sine_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END sine_out[12]
  PIN sine_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END sine_out[13]
  PIN sine_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END sine_out[14]
  PIN sine_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END sine_out[15]
  PIN sine_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END sine_out[1]
  PIN sine_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 94.060 37.440 98.060 38.040 ;
    END
  END sine_out[2]
  PIN sine_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 104.780 58.330 108.780 ;
    END
  END sine_out[3]
  PIN sine_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END sine_out[4]
  PIN sine_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 104.780 39.010 108.780 ;
    END
  END sine_out[5]
  PIN sine_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END sine_out[6]
  PIN sine_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END sine_out[7]
  PIN sine_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 104.780 48.670 108.780 ;
    END
  END sine_out[8]
  PIN sine_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END sine_out[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 92.650 95.390 ;
      LAYER li1 ;
        RECT 5.520 10.795 92.460 95.285 ;
      LAYER met1 ;
        RECT 4.210 10.640 92.460 95.440 ;
      LAYER met2 ;
        RECT 4.230 104.500 38.450 104.780 ;
        RECT 39.290 104.500 48.110 104.780 ;
        RECT 48.950 104.500 57.770 104.780 ;
        RECT 58.610 104.500 90.980 104.780 ;
        RECT 4.230 4.280 90.980 104.500 ;
        RECT 4.230 4.000 44.890 4.280 ;
        RECT 45.730 4.000 57.770 4.280 ;
        RECT 58.610 4.000 90.980 4.280 ;
      LAYER met3 ;
        RECT 3.990 82.640 94.060 95.365 ;
        RECT 4.400 81.240 94.060 82.640 ;
        RECT 3.990 79.240 94.060 81.240 ;
        RECT 4.400 77.840 94.060 79.240 ;
        RECT 3.990 72.440 94.060 77.840 ;
        RECT 4.400 71.040 93.660 72.440 ;
        RECT 3.990 69.040 94.060 71.040 ;
        RECT 4.400 67.640 93.660 69.040 ;
        RECT 3.990 62.240 94.060 67.640 ;
        RECT 3.990 60.840 93.660 62.240 ;
        RECT 3.990 58.840 94.060 60.840 ;
        RECT 4.400 57.440 94.060 58.840 ;
        RECT 3.990 48.640 94.060 57.440 ;
        RECT 4.400 47.240 94.060 48.640 ;
        RECT 3.990 41.840 94.060 47.240 ;
        RECT 4.400 40.440 94.060 41.840 ;
        RECT 3.990 38.440 94.060 40.440 ;
        RECT 4.400 37.040 93.660 38.440 ;
        RECT 3.990 35.040 94.060 37.040 ;
        RECT 4.400 33.640 94.060 35.040 ;
        RECT 3.990 10.715 94.060 33.640 ;
      LAYER met4 ;
        RECT 14.095 19.215 20.640 91.625 ;
        RECT 23.040 19.215 23.940 91.625 ;
        RECT 26.340 19.215 88.025 91.625 ;
  END
END counter
END LIBRARY

