* NGSPICE file created from counter.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

.subckt counter VGND VPWR clk rst sine_out[0] sine_out[10] sine_out[11] sine_out[12]
+ sine_out[13] sine_out[14] sine_out[15] sine_out[1] sine_out[2] sine_out[3] sine_out[4]
+ sine_out[5] sine_out[6] sine_out[7] sine_out[8] sine_out[9]
XTAP_TAPCELL_ROW_24_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_501_ _338_ net23 _350_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__a21bo_1
X_432_ net75 net70 VGND VGND VPWR VPWR _375_ sky130_fd_sc_hd__xnor2_4
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_415_ net74 _347_ net58 VGND VGND VPWR VPWR _358_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_680_ net52 net24 _380_ VGND VGND VPWR VPWR _244_ sky130_fd_sc_hd__or3_1
XFILLER_29_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_594_ _159_ _161_ net39 VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__a21o_1
X_663_ _226_ _227_ net39 VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__a21oi_1
X_732_ net36 _286_ VGND VGND VPWR VPWR _292_ sky130_fd_sc_hd__nand2_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput7 net7 VGND VGND VPWR VPWR sine_out[14] sky130_fd_sc_hd__buf_2
X_646_ _046_ _086_ _166_ net46 VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__a31o_1
X_577_ _061_ _144_ net21 VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__a21oi_1
X_715_ _268_ _271_ _273_ _276_ VGND VGND VPWR VPWR _277_ sky130_fd_sc_hd__a22o_1
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_431_ net77 net74 VGND VGND VPWR VPWR _374_ sky130_fd_sc_hd__or2_2
XFILLER_13_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_500_ net26 _345_ _382_ _356_ _350_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__o32a_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire19 _137_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
X_629_ _076_ _184_ VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__nand2_1
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_414_ net27 net67 VGND VGND VPWR VPWR _357_ sky130_fd_sc_hd__nand2_1
XFILLER_5_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_662_ _383_ _044_ _358_ _377_ VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__a211o_1
X_731_ _288_ _290_ net20 VGND VGND VPWR VPWR _291_ sky130_fd_sc_hd__a21oi_1
X_593_ _134_ _160_ VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_645_ net38 _205_ _209_ _196_ _201_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__a311o_1
Xoutput8 net8 VGND VGND VPWR VPWR sine_out[15] sky130_fd_sc_hd__buf_2
X_576_ _383_ _120_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__nand2_1
X_714_ net22 _055_ _222_ _274_ _275_ VGND VGND VPWR VPWR _276_ sky130_fd_sc_hd__o32a_1
Xoutput10 net10 VGND VGND VPWR VPWR sine_out[2] sky130_fd_sc_hd__buf_2
X_430_ net45 net41 VGND VGND VPWR VPWR _373_ sky130_fd_sc_hd__nand2b_1
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_628_ _021_ _032_ _134_ net46 VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__o211ai_1
X_559_ _349_ net23 VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ net51 net70 VGND VGND VPWR VPWR _356_ sky130_fd_sc_hd__or2_2
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_592_ net46 net71 _348_ _045_ net42 VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__o311a_1
X_661_ net22 _225_ _369_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__or3b_1
X_730_ net31 _289_ VGND VGND VPWR VPWR _290_ sky130_fd_sc_hd__nand2_1
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput11 net11 VGND VGND VPWR VPWR sine_out[3] sky130_fd_sc_hd__buf_2
X_644_ net38 _205_ _209_ _201_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__a31o_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_575_ _139_ _142_ net33 VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__o21a_1
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput9 net9 VGND VGND VPWR VPWR sine_out[1] sky130_fd_sc_hd__buf_2
X_713_ net29 _023_ _063_ net41 VGND VGND VPWR VPWR _275_ sky130_fd_sc_hd__a31o_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_489_ _372_ _053_ _058_ _376_ net37 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__a221o_1
X_558_ _349_ _381_ _036_ net57 VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__a31o_1
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_627_ net25 _190_ _193_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__a21oi_1
XFILLER_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_412_ net59 _350_ _342_ net48 VGND VGND VPWR VPWR _355_ sky130_fd_sc_hd__a211o_1
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_591_ net46 _151_ _158_ _026_ net42 VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__a221o_1
X_660_ net67 _383_ _359_ net59 VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__o211a_1
X_789_ net1 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__inv_2
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_712_ _041_ _088_ _099_ _217_ net44 VGND VGND VPWR VPWR _274_ sky130_fd_sc_hd__o311a_1
Xoutput12 net12 VGND VGND VPWR VPWR sine_out[4] sky130_fd_sc_hd__buf_2
X_643_ net46 _158_ _206_ _208_ net32 VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__a311o_1
X_574_ _035_ _141_ _140_ net49 VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__o211a_1
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_488_ net75 net26 _018_ _054_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__a31o_1
X_557_ _336_ _375_ _051_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__a21o_1
X_626_ _181_ _186_ _192_ net35 VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__o211a_1
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_411_ net65 net74 net78 VGND VGND VPWR VPWR _354_ sky130_fd_sc_hd__and3b_2
X_609_ _380_ _032_ VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__nor2_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_590_ _089_ _157_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__nand2_1
X_788_ net1 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__inv_2
Xoutput13 net13 VGND VGND VPWR VPWR sine_out[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_573_ _380_ _052_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_642_ _339_ _379_ _207_ _357_ net29 VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__o2111a_1
X_711_ net37 _272_ VGND VGND VPWR VPWR _273_ sky130_fd_sc_hd__nor2_1
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_625_ _187_ _191_ net20 VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__a21o_1
X_556_ net34 _118_ _124_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__or3_1
X_487_ net78 net74 net66 VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_20_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ net75 net70 VGND VGND VPWR VPWR _353_ sky130_fd_sc_hd__nand2_2
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_608_ _148_ _172_ _173_ _174_ VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__a22oi_1
X_539_ _106_ _107_ _372_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__o21a_1
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout70 net72 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_787_ net1 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_572_ net67 _001_ net58 VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__a21o_1
Xoutput14 net14 VGND VGND VPWR VPWR sine_out[6] sky130_fd_sc_hd__buf_2
X_641_ net77 _342_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__nand2_1
X_710_ _356_ _179_ net21 VGND VGND VPWR VPWR _272_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_555_ _357_ _376_ _123_ _121_ _372_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__a32o_1
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_486_ net66 _353_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__nand2_1
X_624_ _346_ _361_ net23 net44 VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_20_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_607_ _383_ _044_ net29 VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_538_ _065_ _089_ net27 VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_469_ _020_ _027_ _028_ _029_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__a32o_1
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_4
Xfanout60 tcout\[3\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_786_ net1 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_571_ _119_ _138_ net31 VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__o21a_1
X_640_ _343_ _370_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__and2_1
XFILLER_16_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR sine_out[7] sky130_fd_sc_hd__buf_2
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_769_ net35 _325_ _324_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__mux2_1
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_554_ net23 _122_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__nand2_1
X_485_ net51 net75 VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__and2b_2
X_623_ _186_ _189_ _181_ VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_606_ net63 _383_ _368_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__a21o_1
X_468_ net31 _034_ _037_ _033_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__a31o_1
X_537_ _378_ _022_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__nor2_1
X_399_ net65 net73 net56 VGND VGND VPWR VPWR _342_ sky130_fd_sc_hd__nor3b_2
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout50 tcout\[4\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout72 tcout\[1\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xfanout61 net62 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_8
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_785_ net1 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput16 net16 VGND VGND VPWR VPWR sine_out[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_570_ net58 _345_ net19 VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__nor3_1
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_699_ _260_ _261_ _029_ VGND VGND VPWR VPWR _262_ sky130_fd_sc_hd__o21a_1
X_768_ net20 _248_ net25 VGND VGND VPWR VPWR _325_ sky130_fd_sc_hd__o21a_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_484_ _383_ _045_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__nor2_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_622_ _187_ _188_ net41 VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__a21o_1
X_553_ net62 _375_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__nand2_4
X_605_ net29 _078_ _116_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__and3_1
X_398_ net65 net73 VGND VGND VPWR VPWR _341_ sky130_fd_sc_hd__or2_2
X_467_ net50 net57 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nor2_1
X_536_ net34 _097_ _103_ _104_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__or4_1
Xfanout40 tcout\[6\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout73 net74 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xfanout62 net69 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xfanout51 net55 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_519_ _336_ _001_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__nand2_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_784_ net1 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput17 net17 VGND VGND VPWR VPWR sine_out[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_767_ net38 _373_ _078_ _321_ _323_ VGND VGND VPWR VPWR _324_ sky130_fd_sc_hd__o311a_1
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_698_ _086_ _206_ net46 VGND VGND VPWR VPWR _261_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_552_ _374_ _120_ _119_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__a21o_1
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_483_ _051_ _052_ net26 _361_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a2bb2o_1
X_621_ net51 _346_ _361_ net44 VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_3_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_604_ net45 _115_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__nor2_1
X_397_ net64 net71 VGND VGND VPWR VPWR _340_ sky130_fd_sc_hd__nor2_2
X_466_ net28 _036_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__nand2_1
X_535_ _018_ _022_ _024_ _376_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__o211a_1
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout30 net31 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout74 tcout\[1\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
Xfanout41 net43 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xfanout63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xfanout52 net54 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_449_ net58 _019_ _017_ net49 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__o211ai_1
X_518_ net61 _375_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_783_ net1 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_766_ _319_ _322_ _030_ VGND VGND VPWR VPWR _323_ sky130_fd_sc_hd__a21o_1
X_697_ _346_ net23 _259_ net24 net49 VGND VGND VPWR VPWR _260_ sky130_fd_sc_hd__o221a_1
X_551_ net58 _345_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_620_ _338_ _032_ _066_ _078_ VGND VGND VPWR VPWR _187_ sky130_fd_sc_hd__nand4_1
X_482_ net76 net63 net53 VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__o21ai_2
X_749_ _029_ _307_ _305_ _302_ VGND VGND VPWR VPWR _308_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_3_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_603_ net36 _162_ _170_ _150_ _156_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__a32o_1
X_396_ net63 net53 VGND VGND VPWR VPWR _339_ sky130_fd_sc_hd__and2b_2
X_465_ net73 net66 net78 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand3b_1
X_534_ _038_ _056_ _100_ _102_ tcout\[5\] VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__a221oi_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
Xfanout31 _334_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
Xfanout20 _030_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xfanout53 net54 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
Xfanout64 net69 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
Xfanout75 net76 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_8
X_517_ net49 _359_ _086_ net43 VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__a31oi_1
X_448_ _345_ _018_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_782_ net25 _331_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_765_ _165_ _220_ net30 VGND VGND VPWR VPWR _322_ sky130_fd_sc_hd__o21ai_1
X_696_ net58 _374_ _381_ VGND VGND VPWR VPWR _259_ sky130_fd_sc_hd__o21ai_1
X_550_ net77 _359_ _383_ net67 net58 VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_481_ net75 net70 net61 VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_748_ _148_ _172_ _306_ net46 VGND VGND VPWR VPWR _307_ sky130_fd_sc_hd__a22o_1
X_679_ net32 _242_ VGND VGND VPWR VPWR _243_ sky130_fd_sc_hd__and2_1
X_464_ net74 net67 net77 VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__and3b_1
X_602_ net33 _027_ _163_ _169_ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__a31o_1
X_533_ _379_ _044_ net31 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__a21oi_2
X_395_ net73 net56 VGND VGND VPWR VPWR _338_ sky130_fd_sc_hd__nand2b_4
Xfanout43 tcout\[5\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xfanout21 _377_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
Xfanout32 _333_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
Xfanout76 net79 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_4
Xfanout54 net55 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout65 net68 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
X_516_ net77 _368_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__or2_1
X_447_ net61 net70 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_0_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_781_ _331_ _332_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_7_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_695_ _251_ _257_ VGND VGND VPWR VPWR _258_ sky130_fd_sc_hd__nand2_1
X_764_ net33 _046_ _319_ _320_ net34 VGND VGND VPWR VPWR _321_ sky130_fd_sc_hd__a221o_1
XFILLER_7_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_480_ net75 net70 net61 VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_747_ _341_ _349_ _157_ _283_ VGND VGND VPWR VPWR _306_ sky130_fd_sc_hd__a31o_1
X_678_ net29 _042_ _179_ _241_ _066_ VGND VGND VPWR VPWR _242_ sky130_fd_sc_hd__a32o_1
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_601_ net34 _164_ _168_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__or3b_1
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_394_ net1 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
X_463_ net58 _019_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nand2_1
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_532_ _379_ _044_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__nand2_1
Xfanout33 _333_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xfanout22 _373_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
Xfanout55 net60 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout44 net47 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xfanout77 net79 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
X_446_ _341_ _001_ net27 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a21o_1
XFILLER_13_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout66 net68 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_515_ net56 _353_ _351_ net31 VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__o211ai_1
X_429_ net32 net49 VGND VGND VPWR VPWR _372_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_23_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_780_ net43 _329_ net40 VGND VGND VPWR VPWR _332_ sky130_fd_sc_hd__a21oi_1
Xinput1 rst VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_763_ net45 _147_ VGND VGND VPWR VPWR _320_ sky130_fd_sc_hd__or2_1
X_694_ net33 _252_ _254_ _256_ VGND VGND VPWR VPWR _257_ sky130_fd_sc_hd__a211o_1
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_746_ net48 _303_ _304_ _028_ VGND VGND VPWR VPWR _305_ sky130_fd_sc_hd__o211a_1
X_677_ net72 _344_ _345_ _382_ net26 VGND VGND VPWR VPWR _241_ sky130_fd_sc_hd__a2111o_1
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_393_ net35 VGND VGND VPWR VPWR _337_ sky130_fd_sc_hd__inv_2
XFILLER_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_600_ _046_ _166_ _167_ net21 VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__a31o_1
X_462_ _340_ _382_ _031_ _343_ net47 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__o311a_1
X_531_ net57 _035_ _098_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__or3_1
X_729_ net57 _089_ _122_ _081_ VGND VGND VPWR VPWR _289_ sky130_fd_sc_hd__a31o_1
Xfanout45 net47 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xfanout34 _328_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xfanout67 net68 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
Xfanout78 net79 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_514_ net41 _077_ _083_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__o21ai_1
Xfanout23 _367_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
Xfanout56 net57 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
X_445_ _364_ _386_ net43 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__mux2_1
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_428_ net58 net24 VGND VGND VPWR VPWR _371_ sky130_fd_sc_hd__nand2_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_762_ net30 _157_ VGND VGND VPWR VPWR _319_ sky130_fd_sc_hd__or2_1
X_693_ net19 _244_ _255_ _372_ VGND VGND VPWR VPWR _256_ sky130_fd_sc_hd__o211a_1
XFILLER_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_745_ _334_ net59 net68 net74 VGND VGND VPWR VPWR _304_ sky130_fd_sc_hd__or4_1
XFILLER_7_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_676_ net43 _236_ _238_ _239_ VGND VGND VPWR VPWR _240_ sky130_fd_sc_hd__o22ai_1
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_461_ net77 net67 net59 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__a21bo_2
X_392_ net62 VGND VGND VPWR VPWR _336_ sky130_fd_sc_hd__inv_2
X_530_ _336_ _382_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__nor2_1
X_659_ _216_ _218_ _221_ _223_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__o211ai_1
X_728_ _101_ _287_ net31 _098_ VGND VGND VPWR VPWR _288_ sky130_fd_sc_hd__a211o_1
Xfanout35 tcout\[7\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xfanout24 _352_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
Xfanout46 net47 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xfanout79 tcout\[0\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
Xfanout68 net69 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_1
Xfanout57 net60 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_2
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_444_ net31 _369_ _371_ _385_ VGND VGND VPWR VPWR _386_ sky130_fd_sc_hd__a31o_1
X_513_ net21 _082_ _080_ net39 VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__o211a_1
XFILLER_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_427_ net76 net54 VGND VGND VPWR VPWR _370_ sky130_fd_sc_hd__nand2_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_761_ net25 _318_ _317_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_692_ net26 _350_ net24 VGND VGND VPWR VPWR _255_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_17_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_744_ net28 _002_ _044_ VGND VGND VPWR VPWR _303_ sky130_fd_sc_hd__a21oi_1
X_675_ _379_ _031_ net22 VGND VGND VPWR VPWR _239_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_460_ net76 net69 net55 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a21boi_2
X_391_ net56 VGND VGND VPWR VPWR _335_ sky130_fd_sc_hd__inv_2
X_589_ net63 net72 net53 VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__a21oi_2
X_658_ net28 _122_ _089_ _372_ VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__o211ai_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_727_ net65 _379_ _383_ net56 VGND VGND VPWR VPWR _287_ sky130_fd_sc_hd__a22o_1
Xfanout47 tcout\[4\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
Xfanout36 tcout\[7\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xfanout25 _337_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
Xfanout58 net60 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xfanout69 tcout\[2\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_512_ _338_ _344_ _081_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__o21ba_1
X_443_ net55 _344_ _354_ _384_ net48 VGND VGND VPWR VPWR _385_ sky130_fd_sc_hd__o311a_1
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_426_ net67 net24 _368_ VGND VGND VPWR VPWR _369_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_409_ net77 net74 VGND VGND VPWR VPWR _352_ sky130_fd_sc_hd__and2_1
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_691_ net21 _253_ net38 VGND VGND VPWR VPWR _254_ sky130_fd_sc_hd__o21ai_1
X_760_ net28 _021_ net25 VGND VGND VPWR VPWR _318_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_743_ _296_ _298_ _301_ _328_ VGND VGND VPWR VPWR _302_ sky130_fd_sc_hd__a31oi_1
X_674_ _336_ _383_ _022_ VGND VGND VPWR VPWR _238_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_390_ net45 VGND VGND VPWR VPWR _334_ sky130_fd_sc_hd__inv_2
X_588_ _153_ _155_ net36 VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__a21oi_1
X_726_ _280_ _281_ _282_ _285_ VGND VGND VPWR VPWR _286_ sky130_fd_sc_hd__a31o_1
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_657_ _089_ _122_ net27 VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__a21oi_1
Xfanout37 net40 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
Xfanout59 net60 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
Xfanout48 net50 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
Xfanout26 net28 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_511_ net23 _042_ _350_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_442_ _339_ _375_ VGND VGND VPWR VPWR _384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_709_ net22 _054_ _270_ _269_ net37 VGND VGND VPWR VPWR _271_ sky130_fd_sc_hd__o311a_1
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_425_ net64 net71 net53 VGND VGND VPWR VPWR _368_ sky130_fd_sc_hd__o21bai_2
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_408_ net56 _350_ VGND VGND VPWR VPWR _351_ sky130_fd_sc_hd__nand2_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_690_ net76 _368_ _370_ VGND VGND VPWR VPWR _253_ sky130_fd_sc_hd__o21a_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_673_ net21 _051_ _220_ net37 VGND VGND VPWR VPWR _237_ sky130_fd_sc_hd__o31ai_1
X_742_ net29 _299_ _300_ VGND VGND VPWR VPWR _301_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_587_ net20 _154_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__nand2_1
X_656_ _219_ _220_ _376_ VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__o21ai_1
X_725_ net22 _062_ _283_ _284_ net34 VGND VGND VPWR VPWR _285_ sky130_fd_sc_hd__o311a_1
Xfanout38 net40 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
Xfanout49 net50 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
Xfanout27 net28 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
X_441_ net74 net77 VGND VGND VPWR VPWR _383_ sky130_fd_sc_hd__nand2b_4
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_510_ _078_ _079_ net22 VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__a21o_1
X_639_ net30 _202_ _204_ VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__a21o_1
X_708_ net26 _050_ _088_ _099_ VGND VGND VPWR VPWR _270_ sky130_fd_sc_hd__o22a_1
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_424_ net56 net73 VGND VGND VPWR VPWR _367_ sky130_fd_sc_hd__nand2b_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ net75 net61 VGND VGND VPWR VPWR _350_ sky130_fd_sc_hd__xnor2_4
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_741_ net48 _347_ _023_ net32 VGND VGND VPWR VPWR _300_ sky130_fd_sc_hd__o31a_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_672_ _334_ _021_ _055_ _096_ _235_ VGND VGND VPWR VPWR _236_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_724_ net60 _377_ _018_ VGND VGND VPWR VPWR _284_ sky130_fd_sc_hd__or3_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_586_ _102_ _134_ _141_ _146_ net39 VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__a221o_1
X_655_ net52 _021_ VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__nor2_1
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout39 net40 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_440_ net72 net75 VGND VGND VPWR VPWR _382_ sky130_fd_sc_hd__and2b_1
Xfanout28 _335_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
X_569_ net77 tcout\[1\] net67 VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__nor3b_1
X_638_ _370_ _122_ _203_ net41 VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__a31o_1
X_707_ _023_ _063_ net21 VGND VGND VPWR VPWR _269_ sky130_fd_sc_hd__a21o_1
X_423_ net52 net71 VGND VGND VPWR VPWR _366_ sky130_fd_sc_hd__and2b_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_406_ net79 net68 VGND VGND VPWR VPWR _349_ sky130_fd_sc_hd__or2_2
XFILLER_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_740_ _018_ _055_ _042_ VGND VGND VPWR VPWR _299_ sky130_fd_sc_hd__o21a_1
X_671_ net27 net65 _379_ net50 VGND VGND VPWR VPWR _235_ sky130_fd_sc_hd__a31o_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_585_ net49 _151_ _152_ net43 VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__a211o_1
X_654_ _340_ net18 VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_18_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_723_ _057_ _179_ VGND VGND VPWR VPWR _283_ sky130_fd_sc_hd__nor2_1
Xfanout29 net31 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
Xfanout18 _001_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
X_637_ _349_ net23 net46 _338_ VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__o211a_1
X_706_ net44 _266_ _267_ net41 VGND VGND VPWR VPWR _268_ sky130_fd_sc_hd__a211o_1
X_499_ net32 _064_ _068_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__and3_1
X_568_ _337_ _125_ _136_ _113_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__a31o_1
X_422_ net64 net24 VGND VGND VPWR VPWR _365_ sky130_fd_sc_hd__nand2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_405_ net76 net63 VGND VGND VPWR VPWR _348_ sky130_fd_sc_hd__nor2_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_670_ _232_ _234_ net35 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_584_ _352_ _032_ _369_ net31 VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__o211a_1
XFILLER_17_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_653_ net44 _365_ _207_ _217_ net41 VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__a41o_1
X_722_ _038_ _278_ _279_ net39 VGND VGND VPWR VPWR _282_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_9_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_636_ net54 _089_ _122_ _120_ _374_ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__a32o_1
X_705_ _340_ net18 net29 net52 VGND VGND VPWR VPWR _267_ sky130_fd_sc_hd__o211a_1
X_498_ _354_ _067_ _066_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__o21ai_1
X_567_ _372_ _129_ _131_ _135_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__a22o_1
X_421_ _355_ _358_ _363_ net49 VGND VGND VPWR VPWR _364_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_619_ net34 _183_ _185_ VGND VGND VPWR VPWR _186_ sky130_fd_sc_hd__and3_1
XFILLER_25_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_404_ net78 net66 VGND VGND VPWR VPWR _347_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_22_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_583_ _035_ _141_ _362_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_721_ _341_ _001_ _049_ _239_ VGND VGND VPWR VPWR _281_ sky130_fd_sc_hd__a31o_1
X_652_ net18 _041_ VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_635_ _197_ _198_ _200_ VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__o21ai_1
X_704_ net79 net52 _197_ VGND VGND VPWR VPWR _266_ sky130_fd_sc_hd__a21o_1
X_566_ _102_ _134_ _133_ net20 VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_497_ net55 _374_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nand2_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_420_ _346_ _362_ VGND VGND VPWR VPWR _363_ sky130_fd_sc_hd__nand2_1
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_549_ _114_ _117_ net32 VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__o21a_1
X_618_ net23 _042_ _184_ net21 VGND VGND VPWR VPWR _185_ sky130_fd_sc_hd__a31o_1
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_403_ net61 net75 VGND VGND VPWR VPWR _346_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_19_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_797_ clknet_1_1__leaf_clk _007_ _015_ VGND VGND VPWR VPWR tcout\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_582_ net34 _143_ _145_ _149_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__or4_1
X_651_ net52 _346_ _122_ _215_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__a31oi_1
X_720_ _351_ _127_ _377_ VGND VGND VPWR VPWR _280_ sky130_fd_sc_hd__a21o_1
X_703_ net25 _258_ _262_ _265_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__o31a_1
XFILLER_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_634_ _055_ net19 _176_ _199_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__or4b_1
X_565_ _366_ _041_ _350_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_496_ net57 _336_ _378_ net48 VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__o31a_1
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_548_ _366_ _025_ _055_ _116_ net46 VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__o311a_1
X_617_ net61 _375_ _359_ net51 VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__o211ai_2
X_479_ net51 _359_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nand2_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_402_ net65 net78 VGND VGND VPWR VPWR _345_ sky130_fd_sc_hd__and2b_2
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_796_ clknet_1_1__leaf_clk _006_ _014_ VGND VGND VPWR VPWR tcout\[6\] sky130_fd_sc_hd__dfrtp_1
X_650_ net24 _041_ _051_ net26 net45 VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__a221o_1
X_779_ net40 net43 _329_ VGND VGND VPWR VPWR _331_ sky130_fd_sc_hd__and3_1
X_581_ _372_ _146_ _148_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__and3_1
XFILLER_3_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_702_ _251_ _257_ _264_ net36 VGND VGND VPWR VPWR _265_ sky130_fd_sc_hd__a31o_1
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_633_ net37 _373_ VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__nor2_1
X_564_ net47 _132_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_495_ net65 _379_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nand2_1
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_547_ net52 net64 net71 VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__nand3b_1
X_478_ net47 _047_ _043_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__o21ai_1
X_616_ _122_ _147_ _182_ net22 VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__a211o_1
X_401_ net76 net62 VGND VGND VPWR VPWR _344_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_19_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_795_ clknet_1_1__leaf_clk _005_ _013_ VGND VGND VPWR VPWR tcout\[5\] sky130_fd_sc_hd__dfrtp_1
X_580_ _340_ _051_ _052_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_4_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_778_ net33 _329_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_29_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_701_ _260_ _263_ _029_ VGND VGND VPWR VPWR _264_ sky130_fd_sc_hd__o21ai_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_632_ _028_ _102_ VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_563_ _350_ _356_ _375_ _045_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__o22a_1
X_494_ _357_ _061_ _063_ net48 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__a31o_1
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_546_ net53 net63 net72 VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__and3b_1
X_477_ net76 _341_ _046_ _031_ net18 VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__a32oi_1
XTAP_TAPCELL_ROW_1_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ net62 net18 _050_ net26 VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__o211a_1
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_400_ net54 _340_ VGND VGND VPWR VPWR _343_ sky130_fd_sc_hd__nand2_1
X_529_ net78 net66 net73 VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__nor3b_1
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_794_ clknet_1_0__leaf_clk _004_ _012_ VGND VGND VPWR VPWR tcout\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_777_ _329_ _330_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__and2b_1
X_700_ net78 _095_ _076_ VGND VGND VPWR VPWR _263_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_631_ net28 _349_ _381_ _036_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__and4_1
X_493_ net26 net18 VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__nand2_1
X_562_ net39 net32 _130_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__or3_1
XFILLER_29_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_476_ net71 _044_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__nand2_1
X_545_ net27 _019_ _355_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_614_ net41 _175_ _180_ net37 VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_459_ net37 net42 VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__or2_1
X_528_ _341_ _062_ _096_ net22 VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__a211oi_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_793_ clknet_1_0__leaf_clk _003_ _011_ VGND VGND VPWR VPWR tcout\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_776_ net24 _044_ net49 VGND VGND VPWR VPWR _330_ sky130_fd_sc_hd__a21o_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_630_ _194_ _195_ net20 VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_492_ net55 _375_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_561_ net57 _019_ _032_ _088_ net48 VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__o221a_1
X_759_ _045_ _078_ _199_ _314_ _316_ VGND VGND VPWR VPWR _317_ sky130_fd_sc_hd__a311o_1
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_613_ _376_ _177_ _178_ _179_ VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__a2bb2o_1
X_475_ net52 net63 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__nand2_2
X_544_ net39 _108_ _112_ net35 _105_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_28_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_389_ net43 VGND VGND VPWR VPWR _333_ sky130_fd_sc_hd__inv_2
X_458_ net37 net41 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__nor2_2
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_527_ net65 net18 _095_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_792_ clknet_1_0__leaf_clk _002_ _010_ VGND VGND VPWR VPWR tcout\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_775_ net50 net24 _044_ VGND VGND VPWR VPWR _329_ sky130_fd_sc_hd__and3_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_491_ net77 _018_ net27 VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__a21o_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_560_ _126_ _127_ _128_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_758_ net30 _339_ _115_ _315_ _029_ VGND VGND VPWR VPWR _316_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_17_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_689_ net44 _062_ _079_ _171_ VGND VGND VPWR VPWR _252_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_474_ net59 net67 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__and2_2
X_612_ net75 net61 net70 net51 VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__o31ai_4
X_543_ net43 _109_ _110_ _111_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__o31ai_1
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_526_ net65 net73 net57 VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_388_ net39 VGND VGND VPWR VPWR _328_ sky130_fd_sc_hd__inv_2
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_457_ net39 net33 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__nor2_1
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_509_ _336_ _375_ _032_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_5_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_791_ clknet_1_1__leaf_clk net18 _009_ VGND VGND VPWR VPWR tcout\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_774_ _347_ _367_ _032_ _338_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__o211ai_1
XFILLER_28_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_490_ net32 _048_ _059_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__a21o_1
X_688_ net49 _144_ _166_ _250_ VGND VGND VPWR VPWR _251_ sky130_fd_sc_hd__a31o_1
X_757_ _115_ _165_ net29 VGND VGND VPWR VPWR _315_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_5_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_473_ _018_ _031_ _041_ net24 net30 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a221o_1
X_611_ net44 _353_ _361_ VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__and3_1
X_542_ net57 _374_ _381_ net21 VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__a31o_1
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_387_ net79 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_456_ _021_ _022_ _026_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_525_ net35 _084_ _094_ _060_ _073_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__a32o_1
X_508_ net76 net71 net63 net52 VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_15_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ net67 net74 VGND VGND VPWR VPWR _381_ sky130_fd_sc_hd__nand2b_1
XFILLER_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_790_ clknet_1_0__leaf_clk _000_ _008_ VGND VGND VPWR VPWR tcout\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_773_ net20 _248_ net35 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__o21a_1
XFILLER_28_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_687_ net49 _023_ _028_ VGND VGND VPWR VPWR _250_ sky130_fd_sc_hd__o21ai_1
X_756_ _310_ _311_ _313_ VGND VGND VPWR VPWR _314_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_5_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_610_ _380_ _032_ net42 _353_ _368_ VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__o2111a_1
X_472_ net51 net61 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__or2_1
X_541_ _339_ _344_ _382_ _338_ net44 VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__o311a_1
X_739_ _342_ net22 _297_ VGND VGND VPWR VPWR _298_ sky130_fd_sc_hd__or3b_1
XFILLER_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_455_ net46 _025_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nor2_1
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_524_ _376_ _024_ _090_ _093_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_30_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_438_ net63 net71 VGND VGND VPWR VPWR _380_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_15_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ _362_ _075_ _076_ _074_ net44 VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__a32o_1
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_772_ _325_ net35 _327_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_755_ _376_ _312_ net34 VGND VGND VPWR VPWR _313_ sky130_fd_sc_hd__a21oi_1
X_686_ _249_ net25 _247_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__mux2_1
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_471_ net51 net62 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nor2_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_540_ net27 _057_ _076_ _362_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__o211a_1
X_669_ net37 _224_ _233_ _029_ _228_ VGND VGND VPWR VPWR _234_ sky130_fd_sc_hd__a221o_1
X_738_ net27 _345_ _360_ _018_ _022_ VGND VGND VPWR VPWR _297_ sky130_fd_sc_hd__o32a_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_454_ net52 _353_ _361_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_523_ _085_ _087_ _092_ _372_ net39 VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_18_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_506_ net48 _055_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__nor2_1
X_437_ net78 net73 VGND VGND VPWR VPWR _379_ sky130_fd_sc_hd__nand2b_2
XFILLER_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_771_ _029_ _248_ _319_ _326_ VGND VGND VPWR VPWR _327_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_754_ net26 _346_ _018_ _353_ _339_ VGND VGND VPWR VPWR _312_ sky130_fd_sc_hd__a32o_1
X_685_ net35 _248_ VGND VGND VPWR VPWR _249_ sky130_fd_sc_hd__and2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_599_ _349_ _157_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__nand2_1
X_470_ net34 _016_ _040_ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__o21bai_1
X_668_ net45 _366_ _021_ _229_ VGND VGND VPWR VPWR _233_ sky130_fd_sc_hd__o31ai_1
X_737_ _184_ _295_ net21 VGND VGND VPWR VPWR _296_ sky130_fd_sc_hd__a21o_1
XFILLER_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_453_ net56 _378_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__nand2_1
X_522_ _347_ net23 _383_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__a31o_1
Xoutput2 net2 VGND VGND VPWR VPWR sine_out[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_505_ _347_ _349_ _049_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__a21o_1
X_436_ net78 net73 VGND VGND VPWR VPWR _378_ sky130_fd_sc_hd__and2b_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_419_ net27 _360_ VGND VGND VPWR VPWR _362_ sky130_fd_sc_hd__nand2_1
X_770_ net45 _147_ net38 net42 VGND VGND VPWR VPWR _326_ sky130_fd_sc_hd__o211a_1
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_753_ net28 _051_ _165_ net45 VGND VGND VPWR VPWR _311_ sky130_fd_sc_hd__a211o_1
X_684_ _021_ _038_ VGND VGND VPWR VPWR _248_ sky130_fd_sc_hd__nand2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_736_ net57 _360_ _021_ VGND VGND VPWR VPWR _295_ sky130_fd_sc_hd__or3_1
X_598_ _339_ net18 VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__nand2_1
X_667_ net37 _224_ _228_ _231_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__a211oi_1
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_452_ net51 net70 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__nand2_2
X_521_ _347_ net23 VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__nor2_1
XFILLER_16_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_719_ net48 _354_ _057_ net32 VGND VGND VPWR VPWR _279_ sky130_fd_sc_hd__o31ai_1
Xoutput3 net3 VGND VGND VPWR VPWR sine_out[10] sky130_fd_sc_hd__buf_2
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_435_ net41 net45 VGND VGND VPWR VPWR _377_ sky130_fd_sc_hd__nand2_2
XFILLER_9_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_504_ net51 net70 _361_ _055_ _054_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_418_ net70 net61 VGND VGND VPWR VPWR _361_ sky130_fd_sc_hd__nand2b_2
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_752_ net45 _309_ net42 VGND VGND VPWR VPWR _310_ sky130_fd_sc_hd__a21o_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_683_ _237_ _240_ _243_ _246_ VGND VGND VPWR VPWR _247_ sky130_fd_sc_hd__o22a_1
XFILLER_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_597_ _339_ _353_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__and2_1
X_666_ _229_ _230_ net20 VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_735_ _291_ _292_ _294_ net36 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__o22a_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_520_ _065_ _089_ net56 VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__a21o_1
X_649_ net25 _211_ _214_ _210_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__o2bb2a_1
Xoutput4 net4 VGND VGND VPWR VPWR sine_out[11] sky130_fd_sc_hd__buf_2
X_718_ _018_ _022_ net48 _338_ VGND VGND VPWR VPWR _278_ sky130_fd_sc_hd__o211a_1
X_451_ net78 net66 net56 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_24_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_434_ net32 net29 VGND VGND VPWR VPWR _376_ sky130_fd_sc_hd__nor2_4
X_503_ _069_ _072_ _337_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__o21a_1
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_417_ net73 net65 VGND VGND VPWR VPWR _360_ sky130_fd_sc_hd__and2b_1
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_682_ _372_ _206_ _244_ _245_ net38 VGND VGND VPWR VPWR _246_ sky130_fd_sc_hd__a221o_1
X_751_ _359_ _051_ net28 VGND VGND VPWR VPWR _309_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_596_ _146_ _148_ net22 VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_665_ _356_ _179_ net44 VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__a21o_1
XFILLER_6_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_734_ net20 _293_ _286_ VGND VGND VPWR VPWR _294_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_27_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ net76 net64 net71 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__nor3_4
Xoutput5 net5 VGND VGND VPWR VPWR sine_out[12] sky130_fd_sc_hd__buf_2
XFILLER_15_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_648_ net35 _213_ VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__nand2_1
X_579_ _340_ _052_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__nor2_1
X_717_ _354_ _057_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _375_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
X_502_ _376_ _070_ _071_ _372_ net34 VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__a221o_1
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_416_ net63 net71 VGND VGND VPWR VPWR _359_ sky130_fd_sc_hd__nand2_2
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_681_ _051_ _052_ _376_ VGND VGND VPWR VPWR _245_ sky130_fd_sc_hd__o21a_1
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_750_ _249_ net25 _308_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__mux2_1
X_595_ _035_ _052_ _140_ VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_664_ _049_ _173_ net29 VGND VGND VPWR VPWR _229_ sky130_fd_sc_hd__a21o_1
X_733_ _128_ _222_ _235_ _288_ VGND VGND VPWR VPWR _293_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_16_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput6 net6 VGND VGND VPWR VPWR sine_out[13] sky130_fd_sc_hd__buf_2
XFILLER_15_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_647_ _194_ _212_ net20 VGND VGND VPWR VPWR _213_ sky130_fd_sc_hd__a21o_1
X_578_ net69 net18 _354_ net58 VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__a211o_1
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_716_ net25 _249_ _277_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__mux2_1
.ends

