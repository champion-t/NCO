VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 509.810 BY 520.530 ;
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END addr0[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 505.810 20.440 509.810 21.040 ;
    END
  END clk
  PIN csb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END csb0
  PIN din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END din0[15]
  PIN din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END din0[1]
  PIN din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END din0[2]
  PIN din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END din0[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 505.810 129.240 509.810 129.840 ;
    END
  END rst
  PIN sine_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END sine_out[0]
  PIN sine_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 293.110 516.530 293.390 520.530 ;
    END
  END sine_out[10]
  PIN sine_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 505.810 312.840 509.810 313.440 ;
    END
  END sine_out[11]
  PIN sine_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 505.810 309.440 509.810 310.040 ;
    END
  END sine_out[12]
  PIN sine_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 505.810 299.240 509.810 299.840 ;
    END
  END sine_out[13]
  PIN sine_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 505.810 306.040 509.810 306.640 ;
    END
  END sine_out[14]
  PIN sine_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 505.810 302.640 509.810 303.240 ;
    END
  END sine_out[15]
  PIN sine_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END sine_out[1]
  PIN sine_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 516.530 216.110 520.530 ;
    END
  END sine_out[2]
  PIN sine_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 516.530 225.770 520.530 ;
    END
  END sine_out[3]
  PIN sine_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 516.530 238.650 520.530 ;
    END
  END sine_out[4]
  PIN sine_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 516.530 248.310 520.530 ;
    END
  END sine_out[5]
  PIN sine_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 516.530 254.750 520.530 ;
    END
  END sine_out[6]
  PIN sine_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 516.530 264.410 520.530 ;
    END
  END sine_out[7]
  PIN sine_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 516.530 277.290 520.530 ;
    END
  END sine_out[8]
  PIN sine_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 516.530 286.950 520.530 ;
    END
  END sine_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 299.170 22.640 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 299.170 176.240 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 298.250 329.840 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 298.250 483.440 508.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 504.400 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 504.400 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 504.400 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 504.400 487.870 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.500 10.640 7.300 302.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 494.620 10.640 496.220 302.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 298.250 25.940 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 298.250 179.540 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 298.250 333.140 508.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 298.250 486.740 508.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 504.400 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 504.400 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 504.400 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 504.400 491.170 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.340 10.640 9.140 302.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 498.300 10.640 499.900 302.160 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 504.350 508.830 ;
      LAYER li1 ;
        RECT 5.520 10.795 504.160 508.725 ;
      LAYER met1 ;
        RECT 4.210 10.640 504.160 508.880 ;
      LAYER met2 ;
        RECT 4.230 516.250 215.550 517.210 ;
        RECT 216.390 516.250 225.210 517.210 ;
        RECT 226.050 516.250 238.090 517.210 ;
        RECT 238.930 516.250 247.750 517.210 ;
        RECT 248.590 516.250 254.190 517.210 ;
        RECT 255.030 516.250 263.850 517.210 ;
        RECT 264.690 516.250 276.730 517.210 ;
        RECT 277.570 516.250 286.390 517.210 ;
        RECT 287.230 516.250 292.830 517.210 ;
        RECT 293.670 516.250 502.690 517.210 ;
        RECT 4.230 4.280 502.690 516.250 ;
        RECT 4.230 4.000 86.750 4.280 ;
        RECT 87.590 4.000 93.190 4.280 ;
        RECT 94.030 4.000 99.630 4.280 ;
        RECT 100.470 4.000 102.850 4.280 ;
        RECT 103.690 4.000 109.290 4.280 ;
        RECT 110.130 4.000 115.730 4.280 ;
        RECT 116.570 4.000 122.170 4.280 ;
        RECT 123.010 4.000 128.610 4.280 ;
        RECT 129.450 4.000 135.050 4.280 ;
        RECT 135.890 4.000 138.270 4.280 ;
        RECT 139.110 4.000 144.710 4.280 ;
        RECT 145.550 4.000 151.150 4.280 ;
        RECT 151.990 4.000 157.590 4.280 ;
        RECT 158.430 4.000 164.030 4.280 ;
        RECT 164.870 4.000 167.250 4.280 ;
        RECT 168.090 4.000 173.690 4.280 ;
        RECT 174.530 4.000 180.130 4.280 ;
        RECT 180.970 4.000 186.570 4.280 ;
        RECT 187.410 4.000 502.690 4.280 ;
      LAYER met3 ;
        RECT 3.990 313.840 505.810 508.805 ;
        RECT 3.990 312.440 505.410 313.840 ;
        RECT 3.990 310.440 505.810 312.440 ;
        RECT 4.400 309.040 505.410 310.440 ;
        RECT 3.990 307.040 505.810 309.040 ;
        RECT 4.400 305.640 505.410 307.040 ;
        RECT 3.990 303.640 505.810 305.640 ;
        RECT 3.990 302.240 505.410 303.640 ;
        RECT 3.990 300.240 505.810 302.240 ;
        RECT 3.990 298.840 505.410 300.240 ;
        RECT 3.990 177.840 505.810 298.840 ;
        RECT 4.400 176.440 505.810 177.840 ;
        RECT 3.990 167.640 505.810 176.440 ;
        RECT 4.400 166.240 505.810 167.640 ;
        RECT 3.990 164.240 505.810 166.240 ;
        RECT 4.400 162.840 505.810 164.240 ;
        RECT 3.990 154.040 505.810 162.840 ;
        RECT 4.400 152.640 505.810 154.040 ;
        RECT 3.990 147.240 505.810 152.640 ;
        RECT 4.400 145.840 505.810 147.240 ;
        RECT 3.990 140.440 505.810 145.840 ;
        RECT 4.400 139.040 505.810 140.440 ;
        RECT 3.990 130.240 505.810 139.040 ;
        RECT 3.990 128.840 505.410 130.240 ;
        RECT 3.990 48.640 505.810 128.840 ;
        RECT 4.400 47.240 505.810 48.640 ;
        RECT 3.990 21.440 505.810 47.240 ;
        RECT 3.990 20.040 505.410 21.440 ;
        RECT 3.990 10.715 505.810 20.040 ;
      LAYER met4 ;
        RECT 20.000 298.770 20.640 385.385 ;
        RECT 23.040 298.770 23.940 385.385 ;
        RECT 20.000 297.850 23.940 298.770 ;
        RECT 26.340 298.770 174.240 385.385 ;
        RECT 176.640 298.770 177.540 385.385 ;
        RECT 26.340 297.850 177.540 298.770 ;
        RECT 179.940 297.850 327.840 385.385 ;
        RECT 330.240 297.850 331.140 385.385 ;
        RECT 333.540 297.850 479.900 385.385 ;
        RECT 20.000 13.775 479.900 297.850 ;
  END
END counter
END LIBRARY

